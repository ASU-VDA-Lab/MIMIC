module fake_netlist_5_1742_n_1743 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1743);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1743;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_2),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_29),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_21),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_47),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_54),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_56),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_33),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_36),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_50),
.Y(n_167)
);

BUFx8_ASAP7_75t_SL g168 ( 
.A(n_95),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_72),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_29),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_30),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_38),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_53),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_126),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_49),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_57),
.Y(n_187)
);

BUFx8_ASAP7_75t_SL g188 ( 
.A(n_42),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_92),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_45),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_58),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_73),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_14),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_137),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_9),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_27),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_68),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_55),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_23),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_45),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_35),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_20),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_34),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_122),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_74),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_143),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_80),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_18),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_37),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_148),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_81),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_39),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_113),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_129),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_112),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_66),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_25),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_21),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_20),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_128),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_13),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_18),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_89),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_59),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_97),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_114),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_61),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_12),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_30),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_15),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_5),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_109),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_6),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_138),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_149),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_96),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_82),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_26),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_142),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_64),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_32),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_36),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_1),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_7),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_93),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_14),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_15),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_67),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_117),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_139),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_86),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_98),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_120),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_85),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_51),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_17),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_76),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_28),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_40),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_102),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_121),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_104),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_13),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_1),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_151),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_40),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_100),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_33),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_44),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_83),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_25),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_28),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_46),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_123),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_35),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_41),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_222),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_182),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_188),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_172),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_198),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_154),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_222),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_164),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_222),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_156),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_156),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_175),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_215),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_175),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_238),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_177),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_169),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_238),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_235),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_169),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_235),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_247),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_178),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_272),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_177),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_191),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_182),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_155),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_215),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_162),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_211),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_165),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_199),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_213),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_221),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_169),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_190),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_237),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_240),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_166),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_224),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_248),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_212),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_160),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_270),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_232),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_177),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_286),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_233),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_234),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_167),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_190),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_173),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_174),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_245),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_249),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_161),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_161),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_205),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_229),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_229),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_179),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_320),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_309),
.B(n_214),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_317),
.B(n_194),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_319),
.B(n_205),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_335),
.B(n_159),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_307),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_310),
.B(n_169),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_194),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_319),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_321),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_321),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_312),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_L g418 ( 
.A(n_342),
.B(n_166),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_380),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_369),
.B(n_243),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_380),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_347),
.B(n_159),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_347),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_352),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_359),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_243),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_356),
.B(n_214),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_316),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_313),
.A2(n_226),
.B1(n_289),
.B2(n_281),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_329),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_184),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_329),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_332),
.B(n_159),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_365),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_391),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_357),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_445),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_445),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_332),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_383),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_408),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_386),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_409),
.A2(n_226),
.B1(n_314),
.B2(n_377),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_404),
.B(n_338),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_389),
.B(n_365),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_393),
.B(n_343),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_418),
.A2(n_367),
.B1(n_374),
.B2(n_373),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_404),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_444),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_395),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

CKINVDCx6p67_ASAP7_75t_R g476 ( 
.A(n_385),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

NOR2x1p5_ASAP7_75t_L g480 ( 
.A(n_400),
.B(n_367),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_398),
.A2(n_356),
.B1(n_344),
.B2(n_346),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_373),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_398),
.B(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_169),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_399),
.B(n_393),
.C(n_435),
.Y(n_490)
);

BUFx8_ASAP7_75t_SL g491 ( 
.A(n_408),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_398),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_411),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_399),
.A2(n_355),
.B1(n_368),
.B2(n_366),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_401),
.B(n_353),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_403),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_339),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_407),
.B(n_197),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_407),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_411),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_326),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_388),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_444),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_192),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_388),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_427),
.B(n_370),
.Y(n_519)
);

OA22x2_ASAP7_75t_L g520 ( 
.A1(n_446),
.A2(n_340),
.B1(n_334),
.B2(n_379),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_394),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

NOR2x1p5_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_176),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_446),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_443),
.A2(n_364),
.B1(n_348),
.B2(n_361),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_396),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_394),
.B(n_220),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_345),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_394),
.B(n_254),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_421),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_409),
.B(n_315),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_441),
.B(n_209),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_410),
.B(n_334),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_435),
.B(n_350),
.C(n_349),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_394),
.B(n_157),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_410),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

BUFx8_ASAP7_75t_SL g545 ( 
.A(n_441),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_402),
.B(n_158),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_429),
.B(n_447),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_447),
.B(n_429),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_443),
.B(n_170),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_384),
.A2(n_264),
.B1(n_195),
.B2(n_256),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_412),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_402),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_423),
.Y(n_555)
);

AND2x2_ASAP7_75t_SL g556 ( 
.A(n_384),
.B(n_192),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_412),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_413),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_413),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_414),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_385),
.A2(n_281),
.B1(n_227),
.B2(n_209),
.Y(n_563)
);

NOR2x1p5_ASAP7_75t_L g564 ( 
.A(n_422),
.B(n_176),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_414),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_415),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_422),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_417),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_415),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_434),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_406),
.B(n_227),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_406),
.B(n_279),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_406),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_402),
.B(n_163),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_417),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_416),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_406),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_434),
.B(n_265),
.Y(n_579)
);

INVxp33_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_420),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_420),
.A2(n_261),
.B1(n_266),
.B2(n_267),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_424),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_417),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_430),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_430),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_424),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_402),
.B(n_180),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_442),
.B(n_279),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_440),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_431),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_387),
.B(n_170),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_437),
.Y(n_596)
);

AO21x2_ASAP7_75t_L g597 ( 
.A1(n_437),
.A2(n_216),
.B(n_285),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_437),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_387),
.B(n_171),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_487),
.A2(n_289),
.B1(n_299),
.B2(n_260),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_492),
.A2(n_299),
.B1(n_244),
.B2(n_241),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_505),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_492),
.B(n_341),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_525),
.B(n_171),
.Y(n_604)
);

NAND2x1_ASAP7_75t_L g605 ( 
.A(n_503),
.B(n_387),
.Y(n_605)
);

INVxp33_ASAP7_75t_SL g606 ( 
.A(n_451),
.Y(n_606)
);

INVx8_ASAP7_75t_L g607 ( 
.A(n_500),
.Y(n_607)
);

AND2x6_ASAP7_75t_SL g608 ( 
.A(n_536),
.B(n_354),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_486),
.B(n_230),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_567),
.B(n_341),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_489),
.B(n_177),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_567),
.A2(n_210),
.B1(n_242),
.B2(n_236),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_520),
.A2(n_207),
.B1(n_231),
.B2(n_218),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_472),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_520),
.A2(n_196),
.B1(n_201),
.B2(n_185),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_525),
.B(n_556),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_489),
.B(n_177),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_556),
.B(n_230),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_490),
.A2(n_570),
.B1(n_504),
.B2(n_483),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_470),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_532),
.A2(n_208),
.B1(n_228),
.B2(n_225),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_454),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_548),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_453),
.B(n_363),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_458),
.A2(n_204),
.B1(n_246),
.B2(n_223),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_587),
.B(n_202),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_454),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_583),
.B(n_302),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_583),
.B(n_302),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_583),
.B(n_303),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_455),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_505),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_587),
.B(n_253),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_453),
.B(n_257),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_459),
.B(n_363),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_452),
.B(n_303),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_517),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_459),
.B(n_464),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_455),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_464),
.B(n_468),
.Y(n_640)
);

BUFx5_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_457),
.B(n_177),
.Y(n_642)
);

AND2x6_ASAP7_75t_SL g643 ( 
.A(n_500),
.B(n_358),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_520),
.A2(n_277),
.B1(n_274),
.B2(n_271),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_470),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_461),
.A2(n_259),
.B1(n_177),
.B2(n_192),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_451),
.B(n_168),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_458),
.A2(n_467),
.B1(n_564),
.B2(n_550),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_489),
.B(n_181),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_456),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_474),
.B(n_417),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_472),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_514),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_580),
.B(n_239),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_456),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_461),
.B(n_438),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_537),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_471),
.B(n_306),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_477),
.B(n_324),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_509),
.B(n_306),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_538),
.B(n_276),
.C(n_250),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_509),
.B(n_183),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_537),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_462),
.B(n_438),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_501),
.B(n_186),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_462),
.B(n_426),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_463),
.B(n_426),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_463),
.B(n_426),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_539),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_531),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_589),
.B(n_187),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_543),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_474),
.B(n_438),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_531),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_482),
.B(n_438),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_543),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_589),
.B(n_251),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_482),
.B(n_426),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_460),
.B(n_239),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_477),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_466),
.B(n_324),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_500),
.Y(n_685)
);

NAND2x1_ASAP7_75t_L g686 ( 
.A(n_503),
.B(n_426),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_551),
.B(n_189),
.Y(n_687)
);

OAI221xp5_ASAP7_75t_L g688 ( 
.A1(n_496),
.A2(n_287),
.B1(n_252),
.B2(n_255),
.C(n_292),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_498),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_573),
.B(n_325),
.Y(n_690)
);

AOI21x1_ASAP7_75t_L g691 ( 
.A1(n_542),
.A2(n_331),
.B(n_328),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_500),
.B(n_239),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_579),
.A2(n_304),
.B1(n_305),
.B2(n_275),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_488),
.B(n_426),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_552),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_466),
.B(n_325),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_488),
.B(n_493),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_498),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_499),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_552),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_540),
.B(n_193),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_493),
.A2(n_283),
.B1(n_200),
.B2(n_203),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_499),
.B(n_438),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_502),
.A2(n_192),
.B1(n_304),
.B2(n_305),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_557),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_549),
.B(n_298),
.C(n_297),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_563),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_582),
.B(n_206),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_502),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_476),
.Y(n_710)
);

BUFx12f_ASAP7_75t_SL g711 ( 
.A(n_579),
.Y(n_711)
);

AOI221xp5_ASAP7_75t_L g712 ( 
.A1(n_473),
.A2(n_291),
.B1(n_268),
.B2(n_327),
.C(n_331),
.Y(n_712)
);

AO221x1_ASAP7_75t_L g713 ( 
.A1(n_573),
.A2(n_192),
.B1(n_557),
.B2(n_576),
.C(n_560),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_590),
.B(n_282),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_560),
.B(n_438),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_561),
.B(n_280),
.Y(n_717)
);

INVx8_ASAP7_75t_L g718 ( 
.A(n_466),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_554),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_562),
.B(n_428),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_564),
.A2(n_278),
.B1(n_219),
.B2(n_258),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_579),
.B(n_328),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_579),
.B(n_327),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_508),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_565),
.A2(n_288),
.B1(n_262),
.B2(n_296),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_508),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_466),
.B(n_217),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_SL g728 ( 
.A1(n_473),
.A2(n_263),
.B1(n_269),
.B2(n_273),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_R g729 ( 
.A(n_577),
.B(n_514),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_566),
.B(n_294),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_524),
.Y(n_731)
);

BUFx5_ASAP7_75t_L g732 ( 
.A(n_596),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_SL g733 ( 
.A(n_514),
.B(n_290),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_523),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_566),
.B(n_428),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_569),
.B(n_428),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_569),
.A2(n_428),
.B1(n_426),
.B2(n_4),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_489),
.B(n_428),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_428),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_576),
.B(n_144),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_578),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_578),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_581),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_591),
.B(n_141),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_591),
.B(n_134),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_526),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_469),
.B(n_130),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_523),
.B(n_3),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_515),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_469),
.B(n_127),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_494),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_478),
.B(n_116),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_595),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_494),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_497),
.B(n_10),
.C(n_11),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_480),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_515),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_516),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_516),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_518),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_523),
.B(n_10),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_530),
.B(n_11),
.Y(n_762)
);

NOR2x1p5_ASAP7_75t_L g763 ( 
.A(n_476),
.B(n_16),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_478),
.B(n_115),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_596),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_533),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_610),
.B(n_522),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_610),
.B(n_479),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_623),
.B(n_519),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_603),
.B(n_641),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_683),
.B(n_572),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_614),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_614),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_602),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_673),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_632),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_653),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_603),
.B(n_479),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_614),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_754),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_641),
.B(n_481),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_756),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_689),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_649),
.B(n_599),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_653),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_719),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_619),
.B(n_465),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_751),
.A2(n_640),
.B(n_638),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_641),
.B(n_638),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_606),
.Y(n_790)
);

BUFx4f_ASAP7_75t_L g791 ( 
.A(n_607),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_637),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_481),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_620),
.B(n_546),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_677),
.B(n_510),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_641),
.B(n_640),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_660),
.A2(n_489),
.B1(n_510),
.B2(n_597),
.Y(n_797)
);

INVx6_ASAP7_75t_L g798 ( 
.A(n_683),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_723),
.Y(n_799)
);

OR2x2_ASAP7_75t_SL g800 ( 
.A(n_669),
.B(n_491),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_645),
.Y(n_801)
);

BUFx12f_ASAP7_75t_L g802 ( 
.A(n_643),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_754),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_654),
.B(n_574),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_654),
.B(n_588),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_698),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_699),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_495),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_697),
.B(n_495),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_718),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_SL g812 ( 
.A(n_600),
.B(n_577),
.C(n_545),
.Y(n_812)
);

AND2x6_ASAP7_75t_L g813 ( 
.A(n_740),
.B(n_485),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_718),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_656),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_609),
.B(n_485),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_659),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_719),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_646),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_697),
.B(n_484),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_665),
.B(n_675),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_754),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_679),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_722),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_607),
.B(n_484),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_700),
.B(n_489),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_705),
.B(n_597),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_682),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_SL g830 ( 
.A(n_712),
.B(n_598),
.C(n_594),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_616),
.A2(n_511),
.B1(n_597),
.B2(n_598),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_746),
.A2(n_511),
.B(n_593),
.C(n_592),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_707),
.A2(n_544),
.B1(n_506),
.B2(n_512),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_680),
.B(n_594),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_716),
.B(n_544),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_624),
.A2(n_544),
.B(n_506),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_711),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_684),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_628),
.B(n_535),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_741),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_629),
.B(n_535),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_731),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_742),
.B(n_475),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_630),
.B(n_674),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_661),
.B(n_593),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_743),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_751),
.A2(n_584),
.B(n_575),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_765),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_672),
.A2(n_475),
.B1(n_506),
.B2(n_512),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_661),
.B(n_592),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_655),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_624),
.B(n_475),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_734),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_635),
.B(n_568),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_739),
.A2(n_586),
.B1(n_585),
.B2(n_529),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_635),
.B(n_568),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_718),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_733),
.B(n_512),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_728),
.B(n_503),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_684),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_696),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_696),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_763),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_676),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_607),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_612),
.B(n_494),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_745),
.B(n_568),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_724),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_745),
.B(n_744),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_685),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_730),
.B(n_721),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_729),
.Y(n_872)
);

AND2x6_ASAP7_75t_L g873 ( 
.A(n_748),
.B(n_586),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_676),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_739),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_732),
.B(n_585),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_732),
.B(n_518),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_692),
.B(n_761),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_732),
.B(n_613),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_726),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_732),
.B(n_521),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_618),
.A2(n_521),
.B1(n_528),
.B2(n_559),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_636),
.B(n_528),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_749),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_678),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_663),
.B(n_494),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_690),
.B(n_553),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_601),
.A2(n_547),
.B1(n_529),
.B2(n_559),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_732),
.B(n_541),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_687),
.A2(n_541),
.B1(n_534),
.B2(n_553),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_739),
.Y(n_891)
);

INVx8_ASAP7_75t_L g892 ( 
.A(n_690),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_615),
.B(n_534),
.Y(n_893)
);

AND2x6_ASAP7_75t_SL g894 ( 
.A(n_690),
.B(n_19),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_710),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_662),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_604),
.B(n_555),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_747),
.Y(n_898)
);

O2A1O1Ixp5_ASAP7_75t_L g899 ( 
.A1(n_717),
.A2(n_555),
.B(n_575),
.C(n_584),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_678),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_644),
.B(n_575),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_706),
.B(n_535),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_701),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_762),
.Y(n_904)
);

BUFx8_ASAP7_75t_SL g905 ( 
.A(n_648),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_681),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_634),
.B(n_558),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_SL g908 ( 
.A(n_693),
.B(n_22),
.C(n_23),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_625),
.B(n_558),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_727),
.B(n_558),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_681),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_715),
.B(n_558),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_621),
.B(n_558),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_714),
.B(n_24),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_747),
.B(n_513),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_667),
.B(n_513),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_608),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_626),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_633),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_664),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_715),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_757),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_720),
.B(n_513),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_755),
.B(n_79),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_758),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_688),
.B(n_26),
.C(n_31),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_759),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_702),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_622),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_760),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_708),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_720),
.B(n_513),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_735),
.B(n_513),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_627),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_753),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_642),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_631),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_735),
.B(n_507),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_639),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_736),
.B(n_507),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_L g941 ( 
.A(n_750),
.B(n_507),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_642),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_725),
.B(n_736),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_651),
.B(n_657),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_704),
.B(n_507),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_703),
.B(n_507),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_750),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_652),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_694),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_752),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_775),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_929),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_789),
.A2(n_737),
.B1(n_766),
.B2(n_647),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_777),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_824),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_SL g956 ( 
.A1(n_914),
.A2(n_764),
.B(n_752),
.C(n_650),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_819),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_838),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_796),
.A2(n_770),
.B(n_869),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_929),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_797),
.A2(n_703),
.B1(n_764),
.B2(n_670),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_810),
.B(n_686),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_770),
.A2(n_605),
.B(n_738),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_879),
.A2(n_668),
.B1(n_671),
.B2(n_670),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_864),
.B(n_666),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_878),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_918),
.B(n_666),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_774),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_776),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_788),
.A2(n_671),
.B(n_668),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_821),
.B(n_658),
.Y(n_971)
);

CKINVDCx10_ASAP7_75t_R g972 ( 
.A(n_800),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_SL g973 ( 
.A1(n_769),
.A2(n_713),
.B1(n_617),
.B2(n_611),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_829),
.Y(n_974)
);

OAI22x1_ASAP7_75t_L g975 ( 
.A1(n_787),
.A2(n_691),
.B1(n_658),
.B2(n_39),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_815),
.B(n_32),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_917),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_792),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_879),
.A2(n_43),
.B1(n_48),
.B2(n_75),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_795),
.B(n_43),
.Y(n_980)
);

BUFx2_ASAP7_75t_SL g981 ( 
.A(n_895),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_939),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_939),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_868),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_874),
.B(n_84),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_SL g986 ( 
.A1(n_871),
.A2(n_87),
.B(n_90),
.C(n_94),
.Y(n_986)
);

NOR2x1_ASAP7_75t_L g987 ( 
.A(n_853),
.B(n_99),
.Y(n_987)
);

CKINVDCx8_ASAP7_75t_R g988 ( 
.A(n_851),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_810),
.B(n_105),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_SL g990 ( 
.A(n_928),
.B(n_108),
.C(n_812),
.Y(n_990)
);

INVx6_ASAP7_75t_L g991 ( 
.A(n_865),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_931),
.B(n_799),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_935),
.A2(n_821),
.B1(n_875),
.B2(n_891),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_777),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_771),
.B(n_844),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_861),
.B(n_771),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_943),
.A2(n_784),
.B(n_904),
.C(n_924),
.Y(n_997)
);

INVx3_ASAP7_75t_SL g998 ( 
.A(n_872),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_875),
.A2(n_891),
.B1(n_820),
.B2(n_809),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_857),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_794),
.B(n_919),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_860),
.B(n_862),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_926),
.A2(n_908),
.B(n_924),
.C(n_834),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_858),
.B(n_859),
.C(n_841),
.Y(n_1004)
);

O2A1O1Ixp5_ASAP7_75t_L g1005 ( 
.A1(n_886),
.A2(n_866),
.B(n_913),
.C(n_910),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_801),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_903),
.A2(n_942),
.B(n_896),
.C(n_839),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_773),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_885),
.B(n_900),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_809),
.A2(n_767),
.B(n_803),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_880),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_817),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_906),
.B(n_911),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_823),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_920),
.B(n_826),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_767),
.A2(n_803),
.B(n_780),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_780),
.A2(n_803),
.B(n_808),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_813),
.A2(n_902),
.B1(n_845),
.B2(n_850),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_936),
.A2(n_845),
.B1(n_850),
.B2(n_830),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_773),
.B(n_779),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_875),
.A2(n_891),
.B1(n_846),
.B2(n_840),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_773),
.B(n_779),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_828),
.A2(n_816),
.B(n_867),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_836),
.A2(n_778),
.B(n_768),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_780),
.A2(n_803),
.B(n_781),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_785),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_848),
.A2(n_897),
.B(n_883),
.C(n_909),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_875),
.A2(n_891),
.B1(n_921),
.B2(n_901),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_944),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_SL g1030 ( 
.A(n_780),
.B(n_825),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_813),
.B(n_948),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_884),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_793),
.A2(n_867),
.B(n_907),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_870),
.B(n_782),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_907),
.A2(n_778),
.B(n_912),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_887),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_912),
.A2(n_876),
.B(n_877),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_950),
.A2(n_947),
.B(n_901),
.C(n_902),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_836),
.A2(n_768),
.B(n_856),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_857),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_813),
.B(n_949),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_893),
.A2(n_831),
.B(n_832),
.C(n_828),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_842),
.B(n_772),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_944),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_813),
.A2(n_887),
.B1(n_798),
.B2(n_805),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_837),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_922),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_785),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_852),
.A2(n_854),
.B(n_856),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_791),
.B(n_865),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_852),
.A2(n_854),
.B(n_893),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_786),
.B(n_818),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_798),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_791),
.A2(n_818),
.B1(n_786),
.B2(n_798),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_772),
.B(n_892),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_857),
.B(n_865),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_892),
.B(n_814),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_892),
.B(n_814),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_925),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_827),
.A2(n_783),
.B(n_811),
.C(n_806),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_927),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_898),
.B(n_807),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_804),
.A2(n_873),
.B1(n_916),
.B2(n_937),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_898),
.B(n_905),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_898),
.B(n_930),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_934),
.B(n_843),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_SL g1067 ( 
.A(n_833),
.B(n_827),
.C(n_882),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_899),
.A2(n_843),
.B(n_835),
.C(n_849),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_835),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_855),
.A2(n_915),
.B(n_941),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_881),
.A2(n_889),
.B(n_847),
.Y(n_1071)
);

CKINVDCx6p67_ASAP7_75t_R g1072 ( 
.A(n_802),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_822),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_822),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_945),
.B(n_923),
.Y(n_1075)
);

OAI22x1_ASAP7_75t_L g1076 ( 
.A1(n_894),
.A2(n_890),
.B1(n_863),
.B2(n_873),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_825),
.B(n_888),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_825),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_873),
.A2(n_923),
.B1(n_932),
.B2(n_933),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_873),
.A2(n_932),
.B1(n_933),
.B2(n_938),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_938),
.B(n_940),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_940),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_946),
.B(n_815),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_789),
.B(n_796),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_892),
.B(n_607),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_SL g1086 ( 
.A1(n_789),
.A2(n_796),
.B(n_492),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_775),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_857),
.Y(n_1088)
);

CKINVDCx16_ASAP7_75t_R g1089 ( 
.A(n_853),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_815),
.B(n_769),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1071),
.A2(n_970),
.B(n_1037),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_951),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_980),
.A2(n_966),
.B1(n_995),
.B2(n_1004),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_SL g1094 ( 
.A1(n_1003),
.A2(n_997),
.B1(n_979),
.B2(n_975),
.C(n_953),
.Y(n_1094)
);

AOI211x1_ASAP7_75t_L g1095 ( 
.A1(n_968),
.A2(n_1006),
.B(n_1012),
.C(n_978),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_SL g1096 ( 
.A1(n_966),
.A2(n_1001),
.B(n_979),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_969),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1050),
.B(n_996),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1090),
.B(n_957),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1029),
.B(n_1044),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1009),
.A2(n_1013),
.B1(n_971),
.B2(n_1019),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_SL g1102 ( 
.A1(n_1030),
.A2(n_985),
.B(n_1027),
.Y(n_1102)
);

NAND3x1_ASAP7_75t_L g1103 ( 
.A(n_1064),
.B(n_1057),
.C(n_1058),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_955),
.B(n_957),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1014),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1047),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1046),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1015),
.B(n_1036),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_SL g1109 ( 
.A(n_1054),
.B(n_993),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1061),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1086),
.A2(n_1042),
.B(n_1035),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_984),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1011),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_SL g1114 ( 
.A1(n_1038),
.A2(n_1053),
.B(n_961),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1033),
.A2(n_963),
.B(n_1023),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_988),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1053),
.A2(n_961),
.B(n_1054),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1049),
.A2(n_1051),
.B(n_964),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1036),
.B(n_958),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1000),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1032),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1059),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1077),
.A2(n_965),
.B1(n_1069),
.B2(n_953),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_967),
.B(n_1082),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_952),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1049),
.A2(n_1024),
.B(n_1010),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_960),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1024),
.A2(n_1039),
.B(n_956),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_982),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1066),
.B(n_965),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_983),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1039),
.A2(n_1051),
.B(n_1081),
.Y(n_1132)
);

OA21x2_ASAP7_75t_L g1133 ( 
.A1(n_1005),
.A2(n_1068),
.B(n_1080),
.Y(n_1133)
);

AND3x4_ASAP7_75t_L g1134 ( 
.A(n_990),
.B(n_987),
.C(n_972),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1075),
.A2(n_1079),
.B(n_964),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_999),
.A2(n_1016),
.B(n_1070),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1065),
.B(n_992),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_985),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1018),
.A2(n_993),
.B1(n_1007),
.B2(n_1045),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_1087),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_1089),
.B(n_981),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1073),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1002),
.B(n_1083),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1031),
.A2(n_1041),
.B(n_1063),
.Y(n_1144)
);

AO21x2_ASAP7_75t_L g1145 ( 
.A1(n_999),
.A2(n_1028),
.B(n_1067),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_998),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1034),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1060),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1028),
.A2(n_1021),
.B(n_986),
.C(n_976),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_973),
.A2(n_1021),
.B(n_1062),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_991),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_1070),
.A2(n_1052),
.B(n_1020),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_954),
.A2(n_1026),
.B(n_1048),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1022),
.A2(n_954),
.B(n_1048),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1074),
.A2(n_1078),
.B(n_1056),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1043),
.B(n_1026),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_994),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_994),
.B(n_974),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_962),
.A2(n_989),
.B(n_1055),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_962),
.A2(n_1085),
.B(n_989),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_977),
.B(n_1085),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_991),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1008),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_1000),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1076),
.A2(n_1008),
.A3(n_1085),
.B(n_1040),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1000),
.A2(n_1040),
.B(n_1088),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1040),
.B(n_1088),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1088),
.A2(n_796),
.B(n_789),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1072),
.A2(n_796),
.B(n_789),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_968),
.Y(n_1170)
);

NOR2x1_ASAP7_75t_SL g1171 ( 
.A(n_1054),
.B(n_1004),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_997),
.A2(n_1003),
.B(n_844),
.C(n_914),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_959),
.A2(n_796),
.B(n_789),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_SL g1174 ( 
.A(n_1054),
.B(n_1004),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_959),
.A2(n_796),
.B(n_789),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1084),
.A2(n_1009),
.B1(n_1013),
.B2(n_797),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_980),
.A2(n_787),
.B1(n_444),
.B2(n_995),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_959),
.A2(n_796),
.B(n_789),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1071),
.A2(n_970),
.B(n_1037),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_959),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_997),
.A2(n_1003),
.B(n_844),
.C(n_914),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_966),
.B(n_460),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_SL g1183 ( 
.A1(n_1030),
.A2(n_1003),
.B(n_1009),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_966),
.B(n_460),
.Y(n_1184)
);

NAND3x1_ASAP7_75t_L g1185 ( 
.A(n_980),
.B(n_444),
.C(n_563),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_968),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1084),
.B(n_1029),
.Y(n_1187)
);

AOI221x1_ASAP7_75t_L g1188 ( 
.A1(n_975),
.A2(n_993),
.B1(n_1028),
.B2(n_999),
.C(n_979),
.Y(n_1188)
);

NAND3x1_ASAP7_75t_L g1189 ( 
.A(n_980),
.B(n_444),
.C(n_563),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_980),
.A2(n_787),
.B(n_997),
.C(n_532),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_993),
.A2(n_784),
.B(n_871),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_959),
.A2(n_796),
.B(n_789),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1084),
.B(n_1029),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_966),
.B(n_824),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_968),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1084),
.B(n_1009),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_968),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_959),
.A2(n_796),
.B(n_789),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1084),
.A2(n_1009),
.B1(n_1013),
.B2(n_797),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_999),
.A2(n_1028),
.A3(n_1038),
.B(n_1042),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1053),
.B(n_810),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_997),
.A2(n_1042),
.B(n_1038),
.Y(n_1202)
);

NAND2x1_ASAP7_75t_L g1203 ( 
.A(n_1053),
.B(n_813),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_R g1204 ( 
.A(n_988),
.B(n_790),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1084),
.B(n_1029),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1084),
.B(n_1029),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1084),
.B(n_1009),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_968),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_997),
.A2(n_1003),
.B(n_844),
.C(n_914),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_1042),
.B(n_959),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_968),
.Y(n_1211)
);

CKINVDCx14_ASAP7_75t_R g1212 ( 
.A(n_1072),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_966),
.B(n_824),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1053),
.Y(n_1214)
);

NOR4xp25_ASAP7_75t_L g1215 ( 
.A(n_1003),
.B(n_787),
.C(n_997),
.D(n_753),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_959),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1071),
.A2(n_970),
.B(n_1037),
.Y(n_1217)
);

AOI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1003),
.A2(n_784),
.B(n_787),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1084),
.B(n_1029),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1086),
.A2(n_1042),
.B(n_959),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_968),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_999),
.A2(n_1028),
.A3(n_1038),
.B(n_1042),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1053),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1001),
.B(n_314),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_966),
.B(n_460),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1071),
.A2(n_970),
.B(n_1037),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1188),
.A2(n_1111),
.B(n_1210),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1190),
.A2(n_1181),
.B(n_1172),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1197),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1177),
.A2(n_1218),
.B1(n_1224),
.B2(n_1093),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1119),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1185),
.A2(n_1189),
.B1(n_1207),
.B2(n_1196),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1104),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1218),
.A2(n_1134),
.B1(n_1135),
.B2(n_1101),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1209),
.B(n_1094),
.C(n_1215),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1136),
.A2(n_1128),
.B(n_1111),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1215),
.A2(n_1094),
.B1(n_1135),
.B2(n_1202),
.C(n_1101),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_SL g1238 ( 
.A1(n_1171),
.A2(n_1174),
.B(n_1183),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1203),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1116),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1164),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1097),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1217),
.A2(n_1226),
.B(n_1180),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1147),
.B(n_1098),
.Y(n_1244)
);

CKINVDCx9p33_ASAP7_75t_R g1245 ( 
.A(n_1099),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1194),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1164),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1139),
.A2(n_1191),
.B1(n_1123),
.B2(n_1199),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1118),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1210),
.A2(n_1220),
.B(n_1126),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1216),
.A2(n_1138),
.B(n_1173),
.Y(n_1251)
);

AO21x2_ASAP7_75t_L g1252 ( 
.A1(n_1220),
.A2(n_1102),
.B(n_1132),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1187),
.B(n_1193),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1175),
.A2(n_1178),
.B(n_1192),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1098),
.B(n_1182),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1109),
.A2(n_1145),
.B(n_1150),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1198),
.A2(n_1144),
.B(n_1168),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1212),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1123),
.B(n_1176),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1160),
.A2(n_1159),
.B(n_1153),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1213),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1153),
.A2(n_1148),
.B(n_1139),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1152),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1176),
.A2(n_1199),
.B1(n_1161),
.B2(n_1169),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1155),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1164),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1105),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1145),
.A2(n_1150),
.B(n_1114),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1184),
.B(n_1225),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1170),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1152),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1149),
.A2(n_1117),
.B(n_1133),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1133),
.A2(n_1154),
.B(n_1155),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1130),
.A2(n_1219),
.B1(n_1096),
.B2(n_1108),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1100),
.A2(n_1124),
.B(n_1096),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1200),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1092),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1157),
.A2(n_1110),
.B(n_1106),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1107),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1161),
.A2(n_1141),
.B1(n_1156),
.B2(n_1143),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1186),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1201),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1200),
.B(n_1222),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1204),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1140),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1122),
.A2(n_1112),
.B1(n_1113),
.B2(n_1121),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1195),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1146),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1208),
.A2(n_1221),
.B(n_1211),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1120),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_SL g1292 ( 
.A(n_1120),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1142),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1095),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1129),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1200),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1131),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1222),
.A2(n_1158),
.B(n_1163),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1165),
.B(n_1214),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1151),
.A2(n_1162),
.B1(n_1167),
.B2(n_1214),
.Y(n_1300)
);

BUFx8_ASAP7_75t_L g1301 ( 
.A(n_1120),
.Y(n_1301)
);

OAI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1223),
.A2(n_532),
.B1(n_504),
.B2(n_1190),
.C(n_435),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1165),
.A2(n_1115),
.B(n_1091),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1223),
.A2(n_1190),
.B(n_1181),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1118),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1197),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1307)
);

OAI221xp5_ASAP7_75t_L g1308 ( 
.A1(n_1190),
.A2(n_532),
.B1(n_504),
.B2(n_435),
.C(n_1172),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1164),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_787),
.B1(n_980),
.B2(n_556),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1191),
.A2(n_1188),
.A3(n_1128),
.B(n_1136),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1196),
.B(n_1207),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1224),
.A2(n_1185),
.B1(n_1189),
.B2(n_1134),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1190),
.A2(n_1181),
.B(n_1172),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1197),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1137),
.B(n_1196),
.Y(n_1318)
);

AO21x1_ASAP7_75t_L g1319 ( 
.A1(n_1190),
.A2(n_1218),
.B(n_1135),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1164),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1177),
.A2(n_787),
.B1(n_980),
.B2(n_556),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1177),
.A2(n_787),
.B1(n_980),
.B2(n_556),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1197),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1188),
.A2(n_1111),
.B(n_1220),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1104),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1204),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1197),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_L g1328 ( 
.A(n_1182),
.B(n_790),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1136),
.A2(n_1128),
.B(n_1111),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1116),
.Y(n_1331)
);

CKINVDCx6p67_ASAP7_75t_R g1332 ( 
.A(n_1164),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1107),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1197),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1197),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1136),
.A2(n_1128),
.B(n_1111),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1137),
.B(n_1196),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1339)
);

BUFx10_ASAP7_75t_L g1340 ( 
.A(n_1116),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1098),
.B(n_1078),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1104),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1197),
.Y(n_1343)
);

INVx6_ASAP7_75t_L g1344 ( 
.A(n_1164),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1136),
.A2(n_1128),
.B(n_1111),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1159),
.B(n_1133),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1115),
.A2(n_1179),
.B(n_1091),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1136),
.A2(n_1128),
.B(n_1111),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1190),
.A2(n_1181),
.B(n_1172),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1196),
.B(n_1207),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1197),
.Y(n_1351)
);

AND2x2_ASAP7_75t_SL g1352 ( 
.A(n_1215),
.B(n_556),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1118),
.Y(n_1353)
);

BUFx8_ASAP7_75t_L g1354 ( 
.A(n_1147),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1164),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1231),
.B(n_1246),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1231),
.B(n_1299),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1234),
.A2(n_1310),
.B1(n_1322),
.B2(n_1321),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1273),
.A2(n_1316),
.B(n_1228),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1279),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1326),
.B(n_1286),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1280),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1314),
.B(n_1350),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1315),
.A2(n_1230),
.B1(n_1232),
.B2(n_1308),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1265),
.A2(n_1302),
.B1(n_1338),
.B2(n_1318),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1280),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1319),
.A2(n_1349),
.B(n_1304),
.C(n_1235),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_1326),
.B(n_1240),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1262),
.B(n_1253),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1250),
.A2(n_1254),
.B(n_1337),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1334),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1279),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1314),
.B(n_1350),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1334),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1253),
.B(n_1255),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1275),
.A2(n_1281),
.B(n_1256),
.C(n_1276),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1279),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1273),
.A2(n_1251),
.B(n_1254),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1354),
.Y(n_1379)
);

NOR2x1_ASAP7_75t_SL g1380 ( 
.A(n_1269),
.B(n_1252),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1244),
.B(n_1270),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1238),
.B(n_1263),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1241),
.A2(n_1267),
.B(n_1237),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1233),
.B(n_1325),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1341),
.B(n_1342),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1259),
.A2(n_1352),
.B1(n_1289),
.B2(n_1285),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1306),
.B(n_1317),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1241),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1341),
.B(n_1306),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1259),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1317),
.B(n_1323),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1241),
.A2(n_1267),
.B(n_1250),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1289),
.Y(n_1394)
);

AOI221x1_ASAP7_75t_SL g1395 ( 
.A1(n_1328),
.A2(n_1282),
.B1(n_1268),
.B2(n_1271),
.C(n_1288),
.Y(n_1395)
);

O2A1O1Ixp5_ASAP7_75t_L g1396 ( 
.A1(n_1260),
.A2(n_1249),
.B(n_1305),
.C(n_1353),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1323),
.B(n_1327),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1241),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1250),
.A2(n_1236),
.B(n_1329),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1248),
.A2(n_1260),
.B(n_1263),
.C(n_1293),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1238),
.A2(n_1227),
.B(n_1324),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1266),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1293),
.A2(n_1290),
.B(n_1300),
.C(n_1261),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1287),
.A2(n_1278),
.B1(n_1332),
.B2(n_1227),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1269),
.A2(n_1229),
.B(n_1336),
.C(n_1343),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_SL g1406 ( 
.A1(n_1227),
.A2(n_1324),
.B(n_1269),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1266),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1241),
.A2(n_1267),
.B(n_1324),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1327),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1267),
.A2(n_1355),
.B(n_1320),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1335),
.B(n_1351),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1335),
.A2(n_1351),
.B(n_1257),
.C(n_1296),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1298),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1297),
.B(n_1295),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1332),
.A2(n_1344),
.B1(n_1284),
.B2(n_1294),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1354),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1344),
.A2(n_1284),
.B1(n_1294),
.B2(n_1245),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1354),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1297),
.B(n_1295),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1340),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1277),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1277),
.B(n_1296),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_SL g1423 ( 
.A1(n_1311),
.A2(n_1257),
.B(n_1252),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1267),
.A2(n_1355),
.B(n_1320),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1344),
.A2(n_1247),
.B1(n_1309),
.B2(n_1283),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1247),
.A2(n_1309),
.B(n_1337),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1291),
.B(n_1340),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1345),
.A2(n_1348),
.B(n_1346),
.C(n_1272),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1344),
.B(n_1311),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1311),
.B(n_1348),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1292),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1258),
.A2(n_1274),
.B(n_1243),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1311),
.B(n_1301),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1346),
.A2(n_1239),
.B1(n_1240),
.B2(n_1331),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1346),
.A2(n_1239),
.B1(n_1331),
.B2(n_1264),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1301),
.B(n_1264),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1303),
.B(n_1264),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1292),
.A2(n_1301),
.B1(n_1307),
.B2(n_1312),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1307),
.Y(n_1439)
);

O2A1O1Ixp5_ASAP7_75t_L g1440 ( 
.A1(n_1312),
.A2(n_1347),
.B(n_1330),
.C(n_1333),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1313),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1313),
.B(n_1330),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1333),
.B(n_1339),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1339),
.B(n_1231),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1402),
.B(n_1407),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1444),
.B(n_1430),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1360),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1402),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1372),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1367),
.A2(n_1376),
.B(n_1364),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1357),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1376),
.A2(n_1400),
.B1(n_1367),
.B2(n_1384),
.C(n_1405),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1377),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1359),
.B(n_1429),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1358),
.A2(n_1365),
.B1(n_1387),
.B2(n_1357),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1421),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1363),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1373),
.B(n_1381),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1414),
.B(n_1419),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1437),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1383),
.B(n_1393),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1359),
.B(n_1380),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1437),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1383),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1413),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1442),
.Y(n_1466)
);

BUFx2_ASAP7_75t_SL g1467 ( 
.A(n_1361),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1404),
.A2(n_1403),
.B(n_1405),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_L g1469 ( 
.A(n_1426),
.B(n_1408),
.Y(n_1469)
);

OAI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1385),
.A2(n_1399),
.B(n_1382),
.C(n_1424),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1443),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1396),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1391),
.A2(n_1386),
.B1(n_1420),
.B2(n_1356),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1412),
.B(n_1370),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1413),
.B(n_1396),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1441),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1369),
.B(n_1375),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1409),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1435),
.B(n_1428),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1433),
.B(n_1409),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1417),
.B(n_1378),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1388),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1390),
.B(n_1392),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1411),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1389),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1439),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1432),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1432),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1449),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1465),
.B(n_1438),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1466),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1450),
.B(n_1434),
.C(n_1425),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1465),
.B(n_1415),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1448),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1450),
.A2(n_1418),
.B1(n_1379),
.B2(n_1416),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1454),
.B(n_1440),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1454),
.B(n_1459),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1476),
.B(n_1394),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1464),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1459),
.B(n_1440),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1459),
.B(n_1446),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1488),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1447),
.B(n_1453),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1446),
.B(n_1406),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1463),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1468),
.A2(n_1423),
.B(n_1401),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1486),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1448),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1509),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1493),
.A2(n_1476),
.B1(n_1468),
.B2(n_1455),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1505),
.B(n_1457),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1498),
.B(n_1471),
.Y(n_1514)
);

NAND2xp33_ASAP7_75t_R g1515 ( 
.A(n_1499),
.B(n_1484),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1493),
.A2(n_1452),
.B(n_1469),
.Y(n_1516)
);

OAI33xp33_ASAP7_75t_L g1517 ( 
.A1(n_1505),
.A2(n_1484),
.A3(n_1458),
.B1(n_1456),
.B2(n_1480),
.B3(n_1472),
.Y(n_1517)
);

AOI211xp5_ASAP7_75t_L g1518 ( 
.A1(n_1493),
.A2(n_1452),
.B(n_1470),
.C(n_1476),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1507),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1505),
.A2(n_1470),
.B1(n_1472),
.B2(n_1458),
.C(n_1477),
.Y(n_1520)
);

OAI211xp5_ASAP7_75t_L g1521 ( 
.A1(n_1496),
.A2(n_1469),
.B(n_1473),
.C(n_1480),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1491),
.B(n_1445),
.Y(n_1522)
);

OAI211xp5_ASAP7_75t_L g1523 ( 
.A1(n_1496),
.A2(n_1475),
.B(n_1481),
.C(n_1462),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1502),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1510),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1494),
.A2(n_1467),
.B1(n_1479),
.B2(n_1451),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1491),
.A2(n_1479),
.B(n_1410),
.Y(n_1527)
);

NAND2xp33_ASAP7_75t_R g1528 ( 
.A(n_1499),
.B(n_1427),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1509),
.B(n_1362),
.Y(n_1529)
);

NOR2x1_ASAP7_75t_SL g1530 ( 
.A(n_1508),
.B(n_1461),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1504),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1498),
.B(n_1460),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1500),
.B(n_1460),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_R g1534 ( 
.A(n_1500),
.B(n_1398),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1508),
.A2(n_1479),
.B(n_1474),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1504),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1498),
.B(n_1460),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1504),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1495),
.Y(n_1539)
);

NAND4xp25_ASAP7_75t_L g1540 ( 
.A(n_1491),
.B(n_1475),
.C(n_1478),
.D(n_1368),
.Y(n_1540)
);

NOR4xp25_ASAP7_75t_SL g1541 ( 
.A(n_1495),
.B(n_1451),
.C(n_1487),
.D(n_1467),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1494),
.A2(n_1477),
.B1(n_1475),
.B2(n_1482),
.C(n_1485),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1502),
.B(n_1483),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1510),
.B(n_1445),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1490),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1516),
.A2(n_1479),
.B(n_1474),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1514),
.B(n_1497),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1545),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1525),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1531),
.Y(n_1551)
);

NOR2xp67_ASAP7_75t_L g1552 ( 
.A(n_1535),
.B(n_1492),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_SL g1553 ( 
.A(n_1518),
.B(n_1512),
.C(n_1520),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1536),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1538),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1539),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1540),
.B(n_1371),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1522),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1534),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1521),
.A2(n_1479),
.B(n_1474),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1519),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1544),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1546),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1544),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1546),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1522),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1523),
.A2(n_1489),
.B(n_1503),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1530),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1532),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1534),
.Y(n_1571)
);

NOR2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1511),
.B(n_1500),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1572),
.B(n_1511),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1557),
.B(n_1542),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1550),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1557),
.B(n_1513),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1572),
.B(n_1559),
.Y(n_1577)
);

AND2x2_ASAP7_75t_SL g1578 ( 
.A(n_1568),
.B(n_1515),
.Y(n_1578)
);

AND2x2_ASAP7_75t_SL g1579 ( 
.A(n_1568),
.B(n_1529),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1549),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1572),
.B(n_1532),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1563),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1559),
.B(n_1537),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1549),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1562),
.B(n_1543),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1559),
.B(n_1537),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1524),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1562),
.B(n_1494),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1571),
.B(n_1502),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1549),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1533),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1527),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1550),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1556),
.Y(n_1596)
);

INVxp67_ASAP7_75t_SL g1597 ( 
.A(n_1558),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1533),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1553),
.A2(n_1479),
.B(n_1501),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1565),
.Y(n_1601)
);

CKINVDCx16_ASAP7_75t_R g1602 ( 
.A(n_1553),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1564),
.B(n_1533),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1556),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1563),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1551),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1560),
.A2(n_1517),
.B(n_1541),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1506),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1551),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1563),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1554),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1573),
.B(n_1563),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1573),
.B(n_1563),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1599),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1595),
.B(n_1554),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1573),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1597),
.B(n_1554),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1580),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1593),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1581),
.B(n_1566),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1578),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1577),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1577),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1578),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1574),
.B(n_1570),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1576),
.B(n_1570),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1575),
.B(n_1570),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1584),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1591),
.B(n_1566),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1600),
.A2(n_1560),
.B1(n_1547),
.B2(n_1528),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1589),
.B(n_1607),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1591),
.B(n_1566),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1583),
.B(n_1566),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1590),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1583),
.B(n_1586),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1586),
.Y(n_1644)
);

NOR2x2_ASAP7_75t_L g1645 ( 
.A(n_1582),
.B(n_1564),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1589),
.B(n_1566),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1621),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1618),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1594),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1618),
.Y(n_1650)
);

CKINVDCx16_ASAP7_75t_R g1651 ( 
.A(n_1617),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1612),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1625),
.B(n_1587),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1633),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1637),
.A2(n_1626),
.B1(n_1623),
.B2(n_1615),
.C(n_1627),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1645),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1612),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1620),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

AOI222xp33_ASAP7_75t_L g1660 ( 
.A1(n_1623),
.A2(n_1579),
.B1(n_1560),
.B2(n_1547),
.C1(n_1587),
.C2(n_1601),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1644),
.B(n_1628),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1614),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1615),
.B(n_1594),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1626),
.A2(n_1579),
.B1(n_1547),
.B2(n_1568),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1620),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1630),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1614),
.B(n_1582),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1633),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1630),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1631),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1671),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1651),
.A2(n_1634),
.B1(n_1568),
.B2(n_1643),
.Y(n_1673)
);

OR2x6_ASAP7_75t_L g1674 ( 
.A(n_1647),
.B(n_1639),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1659),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1655),
.A2(n_1634),
.B1(n_1624),
.B2(n_1643),
.C(n_1629),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1648),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1624),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1652),
.B(n_1640),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1658),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1659),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1659),
.Y(n_1683)
);

OAI32xp33_ASAP7_75t_L g1684 ( 
.A1(n_1664),
.A2(n_1656),
.A3(n_1663),
.B1(n_1662),
.B2(n_1657),
.Y(n_1684)
);

AOI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1660),
.A2(n_1616),
.B(n_1610),
.Y(n_1685)
);

AOI32xp33_ASAP7_75t_L g1686 ( 
.A1(n_1664),
.A2(n_1663),
.A3(n_1656),
.B1(n_1667),
.B2(n_1668),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1649),
.A2(n_1616),
.B(n_1619),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1654),
.A2(n_1552),
.B(n_1603),
.C(n_1640),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1654),
.Y(n_1689)
);

OAI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1653),
.A2(n_1636),
.B(n_1635),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1689),
.B(n_1668),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1674),
.B(n_1622),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1674),
.B(n_1680),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1674),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1661),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1682),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1686),
.A2(n_1646),
.B(n_1636),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1672),
.B(n_1635),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1682),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1675),
.B(n_1646),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1683),
.B(n_1687),
.Y(n_1701)
);

AOI211x1_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1684),
.B(n_1687),
.C(n_1673),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1697),
.A2(n_1673),
.B(n_1685),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1696),
.A2(n_1676),
.B1(n_1690),
.B2(n_1679),
.C(n_1681),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1694),
.A2(n_1677),
.B(n_1688),
.Y(n_1705)
);

AOI32xp33_ASAP7_75t_L g1706 ( 
.A1(n_1692),
.A2(n_1693),
.A3(n_1700),
.B1(n_1694),
.B2(n_1699),
.Y(n_1706)
);

NAND4xp25_ASAP7_75t_L g1707 ( 
.A(n_1691),
.B(n_1670),
.C(n_1665),
.D(n_1669),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1698),
.Y(n_1708)
);

NAND4xp25_ASAP7_75t_L g1709 ( 
.A(n_1693),
.B(n_1666),
.C(n_1622),
.D(n_1610),
.Y(n_1709)
);

OAI32xp33_ASAP7_75t_L g1710 ( 
.A1(n_1695),
.A2(n_1619),
.A3(n_1605),
.B1(n_1606),
.B2(n_1641),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1702),
.A2(n_1692),
.B1(n_1622),
.B2(n_1641),
.C(n_1632),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1708),
.B(n_1605),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1703),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1706),
.B(n_1609),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1704),
.A2(n_1631),
.B(n_1632),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1713),
.A2(n_1710),
.B(n_1709),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1712),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1714),
.B(n_1707),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1711),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1715),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1713),
.B(n_1705),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1606),
.B(n_1552),
.C(n_1642),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1717),
.B(n_1719),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1720),
.B(n_1638),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_R g1725 ( 
.A(n_1716),
.B(n_1638),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_L g1726 ( 
.A(n_1718),
.B(n_1642),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1723),
.B(n_1585),
.Y(n_1727)
);

NOR4xp75_ASAP7_75t_SL g1728 ( 
.A(n_1725),
.B(n_1608),
.C(n_1564),
.D(n_1569),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_L g1729 ( 
.A(n_1726),
.B(n_1374),
.C(n_1366),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1727),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1730),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1731),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1731),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_SL g1734 ( 
.A1(n_1733),
.A2(n_1730),
.B(n_1724),
.Y(n_1734)
);

XNOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1732),
.B(n_1729),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1734),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1735),
.A2(n_1722),
.B1(n_1728),
.B2(n_1569),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1736),
.A2(n_1564),
.B1(n_1569),
.B2(n_1596),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1737),
.B1(n_1569),
.B2(n_1564),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1592),
.B(n_1604),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1569),
.B1(n_1604),
.B2(n_1592),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1596),
.B1(n_1611),
.B2(n_1561),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1431),
.B(n_1552),
.C(n_1389),
.Y(n_1743)
);


endmodule