module fake_jpeg_20449_n_210 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_210);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_19),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_46),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_34),
.C(n_31),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_72),
.Y(n_74)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_51),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_30),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_24),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_21),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_44),
.B1(n_23),
.B2(n_16),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_94),
.B1(n_26),
.B2(n_25),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_44),
.B1(n_23),
.B2(n_20),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_69),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_97),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_30),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_31),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_104),
.B1(n_113),
.B2(n_93),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_50),
.B1(n_60),
.B2(n_68),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_114),
.B1(n_117),
.B2(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_87),
.B(n_21),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_60),
.B1(n_48),
.B2(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_118),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_119),
.B(n_97),
.Y(n_132)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_48),
.B1(n_72),
.B2(n_53),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_56),
.B1(n_53),
.B2(n_20),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_26),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_34),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_31),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_95),
.C(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_133),
.C(n_136),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_129),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_119),
.B1(n_107),
.B2(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_94),
.B1(n_79),
.B2(n_91),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_95),
.B1(n_90),
.B2(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_134),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_117),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_86),
.C(n_74),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_74),
.B1(n_92),
.B2(n_89),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_115),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_75),
.C(n_87),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_25),
.B(n_87),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_112),
.B(n_118),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_109),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_138),
.B1(n_129),
.B2(n_132),
.C(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_105),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_149),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_159),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_105),
.C(n_109),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_158),
.C(n_131),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_155),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_102),
.B(n_106),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_156),
.B(n_130),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_102),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_116),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_33),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_127),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_73),
.B(n_18),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_121),
.B1(n_134),
.B2(n_124),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_164),
.B1(n_73),
.B2(n_28),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_136),
.B1(n_127),
.B2(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_169),
.C(n_28),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_143),
.C(n_151),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_145),
.B1(n_128),
.B2(n_21),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_87),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_142),
.A3(n_153),
.B1(n_156),
.B2(n_158),
.C1(n_148),
.C2(n_144),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_177),
.B(n_178),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_161),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_180),
.B(n_168),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_152),
.A3(n_145),
.B1(n_147),
.B2(n_128),
.C1(n_77),
.C2(n_76),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_73),
.B(n_18),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_171),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_169),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_3),
.C(n_4),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_SL g187 ( 
.A(n_184),
.B(n_164),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_162),
.B(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_191),
.Y(n_196)
);

AOI31xp67_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_161),
.A3(n_162),
.B(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_7),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_197),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_176),
.B1(n_183),
.B2(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_176),
.B1(n_184),
.B2(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_189),
.B(n_197),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_204),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_7),
.C(n_8),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_10),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_195),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_203),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_207),
.B(n_11),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_201),
.C(n_202),
.Y(n_209)
);


endmodule