module real_jpeg_16640_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_0),
.Y(n_113)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_1),
.Y(n_309)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_2),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_3),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22x1_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_32),
.B1(n_95),
.B2(n_101),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_3),
.A2(n_32),
.B1(n_277),
.B2(n_281),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_3),
.A2(n_32),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_4),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_4),
.A2(n_119),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_4),
.A2(n_119),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_5),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_6),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_10),
.Y(n_48)
);

OAI22x1_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_48),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_10),
.A2(n_48),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_10),
.B(n_222),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g294 ( 
.A1(n_10),
.A2(n_295),
.A3(n_296),
.B1(n_299),
.B2(n_303),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_10),
.B(n_105),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_10),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_10),
.B(n_57),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_236),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_234),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_198),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_15),
.B(n_198),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_135),
.C(n_174),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_16),
.B(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_54),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_17),
.B(n_55),
.C(n_92),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_19),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_20),
.B(n_48),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_23),
.Y(n_133)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_28),
.B(n_38),
.Y(n_233)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_34),
.Y(n_232)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_47),
.Y(n_37)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_42),
.Y(n_144)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_48),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_48),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_48),
.B(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_51),
.A2(n_137),
.B1(n_141),
.B2(n_147),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_53),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_91),
.B1(n_92),
.B2(n_134),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_73),
.B(n_83),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_57),
.A2(n_73),
.B(n_83),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_57),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_57),
.B(n_276),
.Y(n_311)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_58),
.B(n_274),
.Y(n_273)
);

AOI22x1_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_68),
.Y(n_186)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_68),
.Y(n_298)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_68),
.Y(n_320)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_73),
.B(n_83),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_73),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_73),
.B(n_206),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_80),
.B2(n_82),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_83),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_90),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_114),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_93),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_94),
.B(n_124),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_100),
.Y(n_249)
);

BUFx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2x1p5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_105),
.B(n_115),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_105),
.B(n_220),
.Y(n_219)
);

AO22x2_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_119),
.B(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_124),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_135),
.A2(n_174),
.B1(n_175),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_135),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_148),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_136),
.B(n_148),
.Y(n_215)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_158),
.B(n_161),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_149),
.A2(n_163),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_153),
.Y(n_302)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_161),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_172),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_163),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_167),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_176),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_191),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_182),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_186),
.Y(n_323)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_191),
.B(n_316),
.Y(n_343)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_194),
.Y(n_315)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_214),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_213),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_204),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_205),
.B(n_275),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_226),
.B2(n_227),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_220),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_246),
.A3(n_250),
.B1(n_253),
.B2(n_259),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_289),
.B(n_375),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_286),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_240),
.B(n_286),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.C(n_270),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_241),
.B(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_244),
.A2(n_270),
.B1(n_271),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_244),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_263),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_245),
.B(n_263),
.Y(n_365)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_268),
.B(n_269),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_SL g341 ( 
.A(n_267),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_314),
.B(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_369),
.B(n_374),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_352),
.B(n_368),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_329),
.B(n_351),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_312),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_SL g351 ( 
.A(n_293),
.B(n_312),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_310),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_310),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_324),
.Y(n_312)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_327),
.C(n_367),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_346),
.B(n_350),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_342),
.B(n_345),
.Y(n_330)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_337),
.Y(n_331)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_344),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_349),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_366),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_366),
.Y(n_368)
);

XOR2x2_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_365),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_359),
.B2(n_360),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_360),
.C(n_365),
.Y(n_373)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_373),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_373),
.Y(n_374)
);


endmodule