module fake_jpeg_15088_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_38),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_52),
.B(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_18),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_24),
.B1(n_22),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_22),
.B1(n_24),
.B2(n_34),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_32),
.B(n_33),
.C(n_38),
.Y(n_59)
);

AO22x2_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_62),
.B1(n_57),
.B2(n_50),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_70),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_33),
.B1(n_45),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_34),
.B1(n_48),
.B2(n_54),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_52),
.B1(n_43),
.B2(n_19),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_77),
.Y(n_96)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_22),
.B1(n_24),
.B2(n_29),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_49),
.B1(n_28),
.B2(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_34),
.B1(n_24),
.B2(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_39),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_95),
.B1(n_103),
.B2(n_104),
.Y(n_125)
);

OAI22x1_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_107),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_27),
.B1(n_20),
.B2(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_102),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_49),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_83),
.B(n_25),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_60),
.B1(n_77),
.B2(n_21),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_57),
.C(n_38),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_39),
.B1(n_50),
.B2(n_32),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_35),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_35),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_65),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_121),
.B1(n_96),
.B2(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_127),
.Y(n_151)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_81),
.B1(n_59),
.B2(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_102),
.B1(n_105),
.B2(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_39),
.B1(n_110),
.B2(n_75),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_9),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_58),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_10),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_58),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_131),
.B(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_63),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_26),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_18),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_39),
.B(n_32),
.C(n_67),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_112),
.B(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_92),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_106),
.C(n_94),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_96),
.C(n_98),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_165),
.B1(n_168),
.B2(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_161),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_162),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_165),
.B1(n_168),
.B2(n_117),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_86),
.B1(n_109),
.B2(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_91),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_113),
.B1(n_32),
.B2(n_38),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_117),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_194),
.B1(n_195),
.B2(n_199),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_174),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

CKINVDCx12_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_177),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_128),
.C(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_178),
.Y(n_213)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_185),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_136),
.B(n_25),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_182),
.A2(n_145),
.B(n_152),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_140),
.B(n_169),
.C(n_167),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_188),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_196),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_136),
.B1(n_23),
.B2(n_16),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_23),
.B1(n_16),
.B2(n_120),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_141),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_116),
.B1(n_120),
.B2(n_87),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_141),
.B(n_26),
.Y(n_200)
);

XOR2x1_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_18),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_87),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_147),
.A2(n_38),
.B1(n_16),
.B2(n_35),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_148),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_221),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_144),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_222),
.B(n_228),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_146),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_209),
.C(n_229),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_158),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_224),
.B(n_196),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_170),
.B(n_139),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_140),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_193),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_190),
.B(n_166),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_164),
.B(n_155),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_152),
.C(n_35),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_199),
.B1(n_178),
.B2(n_188),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_223),
.B1(n_213),
.B2(n_204),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_236),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_225),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_181),
.B1(n_182),
.B2(n_180),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_249),
.B1(n_23),
.B2(n_10),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_183),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_241),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_176),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_242),
.B(n_210),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_212),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_247),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_203),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_238),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_189),
.C(n_192),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_23),
.C(n_16),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_228),
.A2(n_202),
.B(n_197),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_227),
.B(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_177),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_243),
.B(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_220),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_256),
.C(n_261),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_242),
.B1(n_256),
.B2(n_237),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_210),
.B1(n_214),
.B2(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_259),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_210),
.B(n_11),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_245),
.C(n_238),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_266),
.C(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_35),
.C(n_18),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_278),
.Y(n_291)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_1),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_282),
.B1(n_267),
.B2(n_11),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_241),
.C(n_232),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_275),
.C(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_234),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_0),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_6),
.C(n_14),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_281),
.B1(n_8),
.B2(n_13),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_254),
.B1(n_251),
.B2(n_266),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_6),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_8),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_252),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_292),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_11),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_35),
.C(n_3),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_5),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_273),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_5),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_283),
.CI(n_272),
.CON(n_298),
.SN(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.Y(n_311)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_5),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_280),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_286),
.C(n_277),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_291),
.B(n_304),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_272),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_312),
.Y(n_317)
);

NOR2x1_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_292),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_313),
.B1(n_305),
.B2(n_302),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_315),
.B(n_313),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_306),
.B(n_297),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_317),
.C(n_12),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_12),
.B(n_13),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_1),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_4),
.Y(n_324)
);


endmodule