module fake_ariane_1954_n_1846 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1846);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1846;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1806;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_114),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_76),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_71),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_65),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_31),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_44),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_97),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_59),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_23),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_60),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_44),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_90),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_78),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_95),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_36),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_63),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_59),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_20),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_63),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_133),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_40),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_22),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_110),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_144),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_61),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_45),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_23),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_31),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_2),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_55),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_154),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_127),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_121),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_149),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_51),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_106),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_52),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_15),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_40),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_108),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_19),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_139),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_79),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_171),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_51),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_142),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_85),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_146),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_93),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_124),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_94),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_120),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_14),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_42),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_27),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_33),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_41),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_17),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_104),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_166),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_168),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_52),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_174),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_164),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_64),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_46),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_74),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_81),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_145),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_118),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_62),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_21),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_16),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_101),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_60),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_62),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_96),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_39),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_107),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_159),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_56),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_119),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_170),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_98),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_34),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_37),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_162),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_1),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_132),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_115),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_65),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_10),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_143),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_123),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_113),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_167),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_12),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_155),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_24),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_102),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_75),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_100),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_131),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_57),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_26),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_129),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_57),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_15),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_158),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_99),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_22),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_10),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_134),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_32),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_58),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_176),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_122),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_126),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_136),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_83),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_173),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_77),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_12),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_156),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_55),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_53),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_73),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_43),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_140),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_6),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_47),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_9),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_24),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_26),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_56),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_49),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_3),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_157),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_50),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_47),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_35),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_181),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_207),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_223),
.B(n_1),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_207),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_182),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_207),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_186),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_179),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_205),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_207),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_208),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_257),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_211),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_219),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_216),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_179),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_220),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_286),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_200),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_253),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_219),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_219),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_219),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_229),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_300),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_253),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_286),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_293),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_232),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_233),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_185),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_222),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_293),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_244),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_198),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_222),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_259),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_259),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_254),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_260),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_256),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_260),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_330),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_193),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_330),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_200),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_258),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_203),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_209),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_340),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_217),
.B(n_3),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_340),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_217),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_269),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_270),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_187),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_189),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_280),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_212),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_276),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_213),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_218),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_231),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_238),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_279),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_200),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_255),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_282),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_291),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_264),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_275),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_292),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_183),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_187),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_277),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_283),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_287),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_267),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_200),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_294),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_297),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_201),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_295),
.Y(n_439)
);

BUFx2_ASAP7_75t_SL g440 ( 
.A(n_273),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_386),
.B(n_215),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_371),
.A2(n_206),
.B(n_202),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_354),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_386),
.B(n_329),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_356),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_371),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_356),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_387),
.B(n_372),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_386),
.B(n_221),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_357),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_L g455 ( 
.A(n_355),
.B(n_200),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_379),
.B(n_273),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_403),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_358),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_362),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_401),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_241),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_364),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_412),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_362),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_422),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_438),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_366),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_373),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_183),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_375),
.A2(n_245),
.B(n_242),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_378),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_409),
.B(n_273),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_385),
.B(n_404),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_385),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_355),
.B(n_215),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_393),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_399),
.A2(n_252),
.B(n_246),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_409),
.B(n_316),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_395),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_261),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_427),
.B(n_301),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_405),
.B(n_278),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_471),
.B(n_353),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_471),
.B(n_353),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_463),
.Y(n_520)
);

AND3x1_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_407),
.C(n_352),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_196),
.C(n_390),
.Y(n_522)
);

AND3x4_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_288),
.C(n_267),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_471),
.B(n_390),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_500),
.A2(n_364),
.B1(n_413),
.B2(n_334),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_455),
.B(n_183),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_477),
.Y(n_527)
);

AND3x2_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_414),
.C(n_439),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_493),
.B(n_183),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_514),
.B(n_439),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_504),
.A2(n_191),
.B1(n_192),
.B2(n_189),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_477),
.Y(n_533)
);

AND3x2_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_251),
.C(n_417),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_454),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_444),
.B(n_359),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_444),
.B(n_361),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_454),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_477),
.B(n_363),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_493),
.B(n_365),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_445),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_448),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_477),
.B(n_367),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_466),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_448),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_466),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_508),
.B(n_369),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_200),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_508),
.B(n_376),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_R g553 ( 
.A(n_458),
.B(n_383),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_508),
.B(n_188),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_450),
.Y(n_557)
);

AOI21x1_ASAP7_75t_L g558 ( 
.A1(n_463),
.A2(n_290),
.B(n_281),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_510),
.A2(n_321),
.B1(n_288),
.B2(n_333),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_514),
.B(n_418),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_468),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_468),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_450),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_468),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_458),
.B(n_384),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_458),
.B(n_389),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_450),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_513),
.B(n_418),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_462),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_462),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_500),
.A2(n_194),
.B1(n_345),
.B2(n_280),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_462),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_514),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_459),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_465),
.B(n_394),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_500),
.B(n_188),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_501),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_441),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_469),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_452),
.B(n_396),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_442),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_469),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_476),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_452),
.B(n_402),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_476),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_501),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_510),
.A2(n_321),
.B1(n_411),
.B2(n_410),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_500),
.A2(n_455),
.B1(n_442),
.B2(n_441),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_465),
.B(n_416),
.Y(n_597)
);

BUFx6f_ASAP7_75t_SL g598 ( 
.A(n_500),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_441),
.B(n_421),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_445),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_452),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_441),
.A2(n_437),
.B1(n_436),
.B2(n_424),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_476),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_479),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_479),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_479),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_481),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_442),
.A2(n_345),
.B1(n_280),
.B2(n_316),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_459),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_481),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_496),
.B(n_428),
.C(n_425),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_441),
.B(n_190),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_513),
.B(n_419),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_483),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_442),
.A2(n_345),
.B1(n_316),
.B2(n_432),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_445),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_445),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_483),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_496),
.B(n_419),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_483),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_483),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_517),
.B(n_190),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_480),
.B(n_200),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_516),
.Y(n_631)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_505),
.A2(n_311),
.B(n_308),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_442),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_483),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_501),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_443),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_480),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_501),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_501),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_445),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_516),
.B(n_420),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_480),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_517),
.B(n_420),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_517),
.A2(n_191),
.B1(n_192),
.B2(n_195),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_501),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_515),
.B(n_423),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_501),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_453),
.B(n_197),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_487),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_443),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_453),
.B(n_423),
.Y(n_651)
);

INVxp33_ASAP7_75t_L g652 ( 
.A(n_515),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_501),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_464),
.A2(n_195),
.B1(n_204),
.B2(n_343),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_464),
.B(n_197),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_502),
.B(n_426),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_446),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_480),
.B(n_250),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_487),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_498),
.B(n_426),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_506),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_502),
.B(n_431),
.Y(n_664)
);

BUFx4f_ASAP7_75t_L g665 ( 
.A(n_487),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_446),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_502),
.B(n_431),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_506),
.B(n_199),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_498),
.B(n_432),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_499),
.B(n_433),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_L g671 ( 
.A(n_536),
.B(n_499),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_636),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_579),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_536),
.B(n_509),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_538),
.B(n_503),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_646),
.B(n_503),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_646),
.B(n_503),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_591),
.A2(n_199),
.B1(n_265),
.B2(n_349),
.Y(n_678)
);

INVxp33_ASAP7_75t_L g679 ( 
.A(n_579),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_555),
.B(n_265),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_578),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_L g682 ( 
.A(n_550),
.B(n_509),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_636),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_512),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_626),
.B(n_512),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_537),
.B(n_480),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_520),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_578),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_526),
.A2(n_487),
.B1(n_507),
.B2(n_506),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_565),
.B(n_586),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_602),
.A2(n_349),
.B1(n_323),
.B2(n_312),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_520),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_627),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_555),
.B(n_506),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_602),
.B(n_507),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_518),
.B(n_506),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_650),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_620),
.B(n_507),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_555),
.B(n_506),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_526),
.A2(n_487),
.B1(n_507),
.B2(n_511),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_620),
.B(n_511),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_650),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_526),
.A2(n_487),
.B1(n_511),
.B2(n_505),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_552),
.B(n_343),
.C(n_204),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_620),
.B(n_511),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_631),
.B(n_511),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_597),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_560),
.B(n_511),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_519),
.B(n_511),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_556),
.Y(n_711)
);

BUFx8_ASAP7_75t_L g712 ( 
.A(n_577),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_596),
.A2(n_351),
.B1(n_350),
.B2(n_348),
.Y(n_713)
);

INVx8_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_560),
.B(n_511),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_560),
.B(n_505),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_651),
.B(n_447),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_524),
.B(n_307),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_561),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_658),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_523),
.A2(n_460),
.B1(n_495),
.B2(n_461),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_658),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_631),
.B(n_344),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_521),
.A2(n_335),
.B1(n_248),
.B2(n_214),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_631),
.B(n_344),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_561),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_662),
.A2(n_447),
.B(n_495),
.C(n_449),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_566),
.B(n_309),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_603),
.B(n_346),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_527),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_533),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_562),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_529),
.B(n_449),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_665),
.A2(n_460),
.B(n_451),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_597),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_523),
.A2(n_467),
.B1(n_451),
.B2(n_461),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_666),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_529),
.B(n_467),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_529),
.B(n_472),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_531),
.B(n_433),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_599),
.B(n_314),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_661),
.A2(n_577),
.B1(n_559),
.B2(n_544),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_533),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_562),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_541),
.B(n_315),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_SL g747 ( 
.A1(n_547),
.A2(n_388),
.B1(n_368),
.B2(n_408),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_531),
.B(n_360),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_583),
.B(n_346),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_529),
.B(n_472),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_583),
.B(n_347),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_529),
.B(n_474),
.Y(n_752)
);

OAI21xp33_ASAP7_75t_L g753 ( 
.A1(n_669),
.A2(n_348),
.B(n_347),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_539),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_540),
.B(n_317),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_529),
.B(n_474),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_666),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_545),
.B(n_318),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_564),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_529),
.B(n_475),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_564),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_598),
.A2(n_296),
.B1(n_338),
.B2(n_306),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_567),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_370),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_567),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_583),
.B(n_350),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_554),
.B(n_570),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_595),
.B(n_351),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_531),
.B(n_322),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_616),
.B(n_325),
.C(n_324),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_539),
.B(n_522),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_569),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_539),
.B(n_336),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_598),
.A2(n_230),
.B1(n_210),
.B2(n_184),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_530),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_530),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_531),
.B(n_381),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_661),
.A2(n_478),
.B1(n_475),
.B2(n_482),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_657),
.A2(n_398),
.B1(n_406),
.B2(n_400),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_532),
.B(n_478),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_657),
.A2(n_337),
.B1(n_341),
.B2(n_342),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_598),
.A2(n_225),
.B1(n_177),
.B2(n_178),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_648),
.B(n_482),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_654),
.B(n_180),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_535),
.Y(n_785)
);

INVx8_ASAP7_75t_L g786 ( 
.A(n_554),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_582),
.B(n_594),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_569),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_657),
.A2(n_382),
.B1(n_484),
.B2(n_490),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_657),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_554),
.B(n_484),
.Y(n_791)
);

INVx4_ASAP7_75t_SL g792 ( 
.A(n_581),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_571),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_525),
.B(n_570),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_571),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_572),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_656),
.B(n_488),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_573),
.B(n_224),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_535),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_572),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_549),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_618),
.B(n_488),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_641),
.B(n_226),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_629),
.B(n_490),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_627),
.B(n_4),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_543),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_554),
.B(n_491),
.Y(n_807)
);

AND2x6_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_188),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_582),
.B(n_480),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_544),
.B(n_4),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_544),
.B(n_5),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_534),
.Y(n_812)
);

BUFx6f_ASAP7_75t_SL g813 ( 
.A(n_554),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_543),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_670),
.B(n_227),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_643),
.B(n_228),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_664),
.B(n_235),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_554),
.B(n_491),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_588),
.B(n_5),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_588),
.A2(n_491),
.B1(n_480),
.B2(n_434),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_644),
.B(n_430),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_582),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_582),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_575),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_667),
.B(n_237),
.Y(n_825)
);

AND2x6_ASAP7_75t_SL g826 ( 
.A(n_547),
.B(n_575),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_588),
.B(n_6),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_665),
.A2(n_491),
.B(n_485),
.C(n_457),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_546),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_576),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_554),
.B(n_239),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_581),
.B(n_240),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_581),
.B(n_243),
.Y(n_833)
);

NOR2x1p5_ASAP7_75t_L g834 ( 
.A(n_553),
.B(n_247),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_581),
.A2(n_304),
.B1(n_249),
.B2(n_262),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_581),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_528),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_581),
.A2(n_305),
.B1(n_263),
.B2(n_266),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_581),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_668),
.B(n_580),
.C(n_576),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_546),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_741),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_690),
.B(n_633),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_768),
.A2(n_617),
.B(n_621),
.C(n_625),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_810),
.A2(n_665),
.B(n_580),
.C(n_587),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_790),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_790),
.B(n_633),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_682),
.B(n_611),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_675),
.B(n_622),
.Y(n_850)
);

BUFx4f_ASAP7_75t_L g851 ( 
.A(n_714),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_732),
.Y(n_853)
);

OAI21xp33_ASAP7_75t_L g854 ( 
.A1(n_678),
.A2(n_605),
.B(n_587),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_685),
.A2(n_600),
.B(n_542),
.Y(n_855)
);

AO21x1_ASAP7_75t_L g856 ( 
.A1(n_810),
.A2(n_633),
.B(n_558),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_SL g857 ( 
.A1(n_747),
.A2(n_319),
.B1(n_284),
.B2(n_289),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_673),
.B(n_548),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_716),
.A2(n_600),
.B(n_542),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_787),
.A2(n_600),
.B(n_542),
.Y(n_860)
);

O2A1O1Ixp5_ASAP7_75t_L g861 ( 
.A1(n_755),
.A2(n_609),
.B(n_617),
.C(n_621),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_755),
.B(n_605),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_607),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_801),
.Y(n_864)
);

AOI21x1_ASAP7_75t_L g865 ( 
.A1(n_707),
.A2(n_632),
.B(n_558),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_743),
.B(n_551),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_741),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_828),
.A2(n_624),
.B(n_640),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_676),
.A2(n_624),
.B(n_640),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_677),
.A2(n_717),
.B(n_710),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_758),
.B(n_607),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_758),
.B(n_608),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_735),
.A2(n_609),
.B(n_608),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_713),
.A2(n_625),
.B(n_628),
.C(n_548),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_732),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_696),
.A2(n_623),
.B(n_624),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_672),
.A2(n_623),
.B1(n_640),
.B2(n_628),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_690),
.B(n_557),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_696),
.A2(n_623),
.B(n_649),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_776),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_708),
.B(n_557),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_710),
.A2(n_614),
.B(n_563),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_701),
.A2(n_614),
.B(n_563),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_811),
.A2(n_632),
.B(n_660),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_736),
.B(n_568),
.Y(n_885)
);

CKINVDCx10_ASAP7_75t_R g886 ( 
.A(n_777),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_706),
.A2(n_699),
.B(n_694),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_687),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_679),
.B(n_568),
.Y(n_889)
);

AOI21xp33_ASAP7_75t_L g890 ( 
.A1(n_746),
.A2(n_649),
.B(n_574),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_698),
.A2(n_610),
.B(n_574),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_776),
.A2(n_615),
.B(n_584),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_681),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_822),
.B(n_594),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_683),
.A2(n_606),
.B1(n_584),
.B2(n_585),
.Y(n_895)
);

AOI21xp33_ASAP7_75t_L g896 ( 
.A1(n_746),
.A2(n_615),
.B(n_601),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_712),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_719),
.B(n_585),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_719),
.B(n_589),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_742),
.B(n_684),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_811),
.A2(n_589),
.B(n_590),
.C(n_592),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_742),
.B(n_590),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_807),
.A2(n_604),
.B(n_592),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_794),
.A2(n_606),
.B1(n_610),
.B2(n_593),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_697),
.B(n_702),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_785),
.A2(n_593),
.B(n_601),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_688),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_743),
.A2(n_551),
.B1(n_659),
.B2(n_630),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_785),
.A2(n_634),
.B(n_612),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_730),
.A2(n_634),
.B(n_612),
.C(n_604),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_792),
.B(n_642),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_721),
.B(n_635),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_704),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_692),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_711),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_704),
.Y(n_916)
);

AOI21xp33_ASAP7_75t_L g917 ( 
.A1(n_729),
.A2(n_663),
.B(n_660),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_799),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_723),
.B(n_635),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_738),
.A2(n_663),
.B1(n_655),
.B2(n_653),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_819),
.A2(n_827),
.B(n_757),
.C(n_725),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_818),
.A2(n_639),
.B(n_655),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_711),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_815),
.A2(n_653),
.B(n_647),
.C(n_645),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_819),
.B(n_594),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_769),
.B(n_638),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_799),
.A2(n_638),
.B(n_647),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_806),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_780),
.B(n_639),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_769),
.B(n_645),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_764),
.B(n_777),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_806),
.A2(n_594),
.B(n_630),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_724),
.B(n_594),
.Y(n_933)
);

NOR2x1_ASAP7_75t_L g934 ( 
.A(n_834),
.B(n_642),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_718),
.A2(n_642),
.B1(n_497),
.B2(n_492),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_814),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_814),
.A2(n_659),
.B(n_457),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_726),
.B(n_7),
.Y(n_938)
);

NOR2x1_ASAP7_75t_R g939 ( 
.A(n_748),
.B(n_268),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_827),
.B(n_619),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_712),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_829),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_820),
.A2(n_497),
.B1(n_492),
.B2(n_489),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_718),
.B(n_271),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_720),
.B(n_272),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_829),
.A2(n_457),
.B(n_485),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_720),
.B(n_727),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_841),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_714),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_822),
.B(n_619),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_841),
.A2(n_457),
.B(n_485),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_748),
.B(n_486),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_753),
.A2(n_485),
.B(n_8),
.C(n_9),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_671),
.A2(n_326),
.B1(n_285),
.B2(n_313),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_728),
.A2(n_637),
.B(n_619),
.Y(n_955)
);

AO21x1_ASAP7_75t_L g956 ( 
.A1(n_686),
.A2(n_250),
.B(n_274),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_727),
.B(n_298),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_733),
.B(n_299),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_733),
.A2(n_328),
.B(n_302),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_745),
.B(n_761),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_745),
.A2(n_331),
.B(n_303),
.Y(n_961)
);

AOI33xp33_ASAP7_75t_L g962 ( 
.A1(n_821),
.A2(n_7),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.B3(n_18),
.Y(n_962)
);

NOR2xp67_ASAP7_75t_L g963 ( 
.A(n_705),
.B(n_637),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_777),
.B(n_486),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_761),
.B(n_674),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_722),
.B(n_737),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_759),
.B(n_310),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_709),
.A2(n_327),
.B(n_332),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_695),
.B(n_11),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_715),
.A2(n_637),
.B(n_619),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_763),
.A2(n_637),
.B(n_619),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_765),
.A2(n_637),
.B(n_619),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_704),
.B(n_637),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_772),
.A2(n_456),
.B(n_470),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_778),
.B(n_13),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_788),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_793),
.A2(n_456),
.B(n_470),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_795),
.A2(n_456),
.B(n_470),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_778),
.B(n_18),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_796),
.A2(n_830),
.B(n_824),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_800),
.A2(n_456),
.B(n_470),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_786),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_802),
.B(n_21),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_729),
.B(n_25),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_704),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_789),
.A2(n_497),
.B1(n_492),
.B2(n_489),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_693),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_802),
.B(n_25),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_822),
.B(n_497),
.Y(n_989)
);

AO21x1_ASAP7_75t_L g990 ( 
.A1(n_805),
.A2(n_250),
.B(n_274),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_767),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_722),
.B(n_28),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_737),
.B(n_497),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_731),
.A2(n_456),
.B(n_470),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_771),
.B(n_28),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_689),
.A2(n_497),
.B1(n_492),
.B2(n_489),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_691),
.B(n_29),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_804),
.B(n_783),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_805),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_804),
.B(n_29),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_783),
.B(n_30),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_797),
.B(n_30),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_797),
.B(n_32),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_837),
.B(n_497),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_744),
.A2(n_816),
.B(n_817),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_820),
.B(n_33),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_825),
.A2(n_456),
.B(n_470),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_840),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_762),
.B(n_34),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_749),
.B(n_35),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_823),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_689),
.A2(n_497),
.B1(n_492),
.B2(n_489),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_751),
.B(n_36),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_766),
.B(n_38),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_784),
.A2(n_38),
.B(n_42),
.C(n_43),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_781),
.B(n_45),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_734),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_792),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_680),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_739),
.A2(n_470),
.B(n_456),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_803),
.B(n_48),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_812),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_822),
.A2(n_456),
.B(n_470),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_770),
.B(n_53),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_700),
.B(n_54),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_823),
.A2(n_473),
.B(n_234),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_700),
.A2(n_703),
.B(n_756),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_773),
.A2(n_54),
.B(n_58),
.C(n_61),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_774),
.B(n_492),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_740),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_703),
.B(n_492),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_750),
.A2(n_473),
.B(n_234),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_982),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_851),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_998),
.A2(n_782),
.B1(n_786),
.B2(n_813),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_897),
.Y(n_1036)
);

NAND2x2_ASAP7_75t_L g1037 ( 
.A(n_1024),
.B(n_826),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_851),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_843),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_976),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_984),
.A2(n_798),
.B(n_752),
.C(n_760),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_907),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_879),
.A2(n_809),
.B(n_791),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_852),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_SL g1045 ( 
.A1(n_925),
.A2(n_831),
.B(n_833),
.C(n_832),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_984),
.A2(n_779),
.B1(n_836),
.B2(n_838),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_842),
.B(n_792),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_900),
.A2(n_835),
.B(n_839),
.C(n_486),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_SL g1049 ( 
.A1(n_921),
.A2(n_813),
.B(n_808),
.C(n_274),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_900),
.B(n_492),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_966),
.B(n_808),
.Y(n_1051)
);

AND3x1_ASAP7_75t_SL g1052 ( 
.A(n_999),
.B(n_274),
.C(n_250),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_921),
.A2(n_489),
.B(n_486),
.C(n_188),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_888),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_893),
.A2(n_808),
.B1(n_489),
.B2(n_486),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_844),
.B(n_489),
.Y(n_1056)
);

AO21x1_ASAP7_75t_L g1057 ( 
.A1(n_925),
.A2(n_808),
.B(n_274),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_852),
.B(n_808),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_844),
.B(n_489),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1001),
.A2(n_1002),
.B1(n_1003),
.B2(n_1000),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_914),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_866),
.B(n_320),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_915),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_SL g1064 ( 
.A(n_949),
.B(n_486),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_842),
.B(n_486),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_897),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_867),
.B(n_486),
.Y(n_1067)
);

OAI22x1_ASAP7_75t_L g1068 ( 
.A1(n_992),
.A2(n_274),
.B1(n_250),
.B2(n_320),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_938),
.A2(n_320),
.B(n_236),
.C(n_234),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_880),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_898),
.A2(n_473),
.B(n_274),
.C(n_250),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_923),
.B(n_250),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_905),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_867),
.B(n_320),
.Y(n_1074)
);

OAI22x1_ASAP7_75t_L g1075 ( 
.A1(n_938),
.A2(n_236),
.B1(n_234),
.B2(n_72),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_941),
.B(n_67),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_907),
.B(n_236),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_983),
.A2(n_236),
.B1(n_473),
.B2(n_82),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_881),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_846),
.A2(n_473),
.B(n_80),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_846),
.A2(n_473),
.B(n_84),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_940),
.A2(n_473),
.B(n_87),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_878),
.B(n_473),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_931),
.B(n_163),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_864),
.B(n_68),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_949),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_952),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_898),
.A2(n_88),
.B(n_89),
.C(n_91),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_911),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_848),
.B(n_103),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_941),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_991),
.B(n_109),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_918),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_940),
.A2(n_111),
.B(n_117),
.Y(n_1094)
);

OAI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_988),
.A2(n_128),
.B(n_130),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1022),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_975),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_926),
.A2(n_160),
.B(n_1016),
.C(n_997),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_911),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_894),
.A2(n_876),
.B(n_871),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_947),
.B(n_960),
.Y(n_1101)
);

OAI22x1_ASAP7_75t_L g1102 ( 
.A1(n_995),
.A2(n_1009),
.B1(n_1006),
.B2(n_979),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_962),
.A2(n_995),
.B(n_872),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_858),
.B(n_889),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_894),
.A2(n_862),
.B(n_860),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_857),
.A2(n_866),
.B1(n_926),
.B2(n_889),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_885),
.B(n_965),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_982),
.Y(n_1108)
);

OAI21xp33_ASAP7_75t_SL g1109 ( 
.A1(n_908),
.A2(n_899),
.B(n_962),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_850),
.A2(n_1008),
.B(n_953),
.C(n_930),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_848),
.B(n_847),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_855),
.A2(n_859),
.B(n_902),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_918),
.B(n_928),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_886),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_933),
.A2(n_1015),
.B(n_1019),
.C(n_849),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_848),
.B(n_847),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_911),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_869),
.A2(n_868),
.B(n_901),
.Y(n_1118)
);

AO32x2_ASAP7_75t_L g1119 ( 
.A1(n_920),
.A2(n_1012),
.A3(n_996),
.B1(n_895),
.B2(n_877),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_964),
.B(n_863),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1010),
.A2(n_1014),
.B(n_1013),
.C(n_1021),
.Y(n_1121)
);

AOI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1005),
.A2(n_980),
.B1(n_887),
.B2(n_968),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_853),
.B(n_875),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_853),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_901),
.A2(n_882),
.B(n_891),
.Y(n_1125)
);

CKINVDCx8_ASAP7_75t_R g1126 ( 
.A(n_939),
.Y(n_1126)
);

AND3x1_ASAP7_75t_SL g1127 ( 
.A(n_987),
.B(n_1028),
.C(n_954),
.Y(n_1127)
);

OAI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_967),
.A2(n_969),
.B(n_854),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_875),
.B(n_913),
.Y(n_1129)
);

NAND2x1p5_ASAP7_75t_L g1130 ( 
.A(n_913),
.B(n_916),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_933),
.A2(n_1025),
.B(n_908),
.C(n_896),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_R g1132 ( 
.A(n_916),
.B(n_985),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1004),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_936),
.B(n_942),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_SL g1135 ( 
.A1(n_1031),
.A2(n_917),
.B(n_989),
.C(n_890),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_874),
.A2(n_861),
.B(n_845),
.C(n_910),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_929),
.A2(n_904),
.B(n_873),
.C(n_986),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_993),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_912),
.A2(n_919),
.B(n_1031),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_927),
.A2(n_909),
.B(n_989),
.Y(n_1140)
);

INVx5_ASAP7_75t_L g1141 ( 
.A(n_985),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1011),
.B(n_958),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_932),
.A2(n_1027),
.B(n_924),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_948),
.B(n_1017),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1011),
.A2(n_934),
.B1(n_944),
.B2(n_945),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_883),
.A2(n_994),
.B(n_856),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_SL g1147 ( 
.A1(n_892),
.A2(n_906),
.B(n_957),
.C(n_1029),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1018),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_948),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_935),
.A2(n_974),
.B(n_977),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_959),
.A2(n_961),
.B(n_943),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_950),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1030),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1030),
.B(n_1018),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_943),
.B(n_973),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_973),
.B(n_963),
.Y(n_1156)
);

INVx3_ASAP7_75t_SL g1157 ( 
.A(n_950),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_978),
.A2(n_981),
.B(n_884),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_990),
.B(n_946),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_955),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1007),
.A2(n_1023),
.B(n_971),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_865),
.A2(n_1020),
.B(n_922),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_903),
.Y(n_1163)
);

INVx3_ASAP7_75t_SL g1164 ( 
.A(n_956),
.Y(n_1164)
);

AOI22x1_ASAP7_75t_L g1165 ( 
.A1(n_1026),
.A2(n_1032),
.B1(n_951),
.B2(n_937),
.Y(n_1165)
);

CKINVDCx6p67_ASAP7_75t_R g1166 ( 
.A(n_972),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_970),
.A2(n_870),
.B(n_879),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_870),
.A2(n_879),
.B(n_998),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_966),
.B(n_866),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_870),
.A2(n_879),
.B(n_998),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_864),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_998),
.B(n_900),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_851),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_995),
.B(n_536),
.C(n_754),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_998),
.B(n_900),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_870),
.A2(n_879),
.B(n_998),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_842),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_900),
.B(n_998),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_852),
.B(n_949),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_870),
.A2(n_879),
.B(n_998),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_870),
.A2(n_879),
.B(n_998),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_984),
.A2(n_921),
.B(n_900),
.C(n_998),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_900),
.B(n_998),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1040),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1182),
.A2(n_1062),
.B(n_1175),
.C(n_1172),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1109),
.A2(n_1060),
.B(n_1080),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1034),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1105),
.A2(n_1100),
.B(n_1062),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1060),
.A2(n_1170),
.B(n_1168),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1054),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1106),
.A2(n_1103),
.B(n_1121),
.C(n_1098),
.Y(n_1194)
);

NAND4xp25_ASAP7_75t_SL g1195 ( 
.A(n_1046),
.B(n_1080),
.C(n_1081),
.D(n_1091),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1115),
.A2(n_1081),
.B(n_1128),
.C(n_1053),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1147),
.A2(n_1137),
.B(n_1131),
.Y(n_1197)
);

NAND3xp33_ASAP7_75t_L g1198 ( 
.A(n_1078),
.B(n_1169),
.C(n_1110),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1176),
.A2(n_1181),
.B(n_1180),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1078),
.B(n_1169),
.C(n_1041),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1163),
.A2(n_1068),
.A3(n_1146),
.B(n_1158),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1161),
.A2(n_1167),
.B(n_1112),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1140),
.A2(n_1125),
.B(n_1150),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1139),
.A2(n_1059),
.B(n_1056),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1102),
.A2(n_1048),
.A3(n_1057),
.B(n_1160),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1136),
.A2(n_1075),
.A3(n_1069),
.B(n_1142),
.Y(n_1206)
);

AOI31xp67_ASAP7_75t_L g1207 ( 
.A1(n_1050),
.A2(n_1145),
.A3(n_1083),
.B(n_1072),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1151),
.A2(n_1073),
.B(n_1095),
.C(n_1107),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1061),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1042),
.B(n_1177),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1104),
.B(n_1079),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1138),
.A2(n_1153),
.B1(n_1035),
.B2(n_1063),
.Y(n_1212)
);

AOI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1159),
.A2(n_1083),
.B(n_1043),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1174),
.A2(n_1101),
.B1(n_1155),
.B2(n_1087),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1171),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1064),
.A2(n_1101),
.B(n_1035),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1148),
.B(n_1034),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1092),
.A2(n_1072),
.A3(n_1113),
.B(n_1134),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1038),
.B(n_1096),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1038),
.B(n_1120),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_1154),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1036),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1070),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1085),
.B(n_1084),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1051),
.A2(n_1120),
.B(n_1090),
.C(n_1082),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1135),
.A2(n_1045),
.B(n_1094),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1122),
.A2(n_1165),
.B(n_1144),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1179),
.B(n_1047),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1049),
.A2(n_1097),
.B(n_1071),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1097),
.A2(n_1116),
.B(n_1111),
.C(n_1154),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1055),
.A2(n_1077),
.B(n_1127),
.Y(n_1231)
);

AOI221xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1123),
.A2(n_1133),
.B1(n_1067),
.B2(n_1074),
.C(n_1065),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1126),
.B(n_1157),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1093),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1156),
.A2(n_1129),
.B(n_1173),
.C(n_1033),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1124),
.B(n_1088),
.C(n_1141),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1164),
.A2(n_1152),
.B(n_1130),
.C(n_1033),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1066),
.B(n_1114),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1119),
.A2(n_1124),
.B(n_1130),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1149),
.A2(n_1124),
.B(n_1058),
.C(n_1141),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1044),
.B(n_1086),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1119),
.A2(n_1052),
.A3(n_1166),
.B(n_1108),
.Y(n_1242)
);

AO21x2_ASAP7_75t_L g1243 ( 
.A1(n_1132),
.A2(n_1119),
.B(n_1058),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1044),
.B(n_1086),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1076),
.B(n_1086),
.Y(n_1245)
);

OAI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1037),
.A2(n_1089),
.B1(n_1099),
.B2(n_1117),
.Y(n_1246)
);

NOR4xp25_ASAP7_75t_L g1247 ( 
.A(n_1089),
.B(n_1182),
.C(n_921),
.D(n_1103),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1040),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1182),
.A2(n_921),
.B(n_1109),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1042),
.B(n_673),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1060),
.A2(n_856),
.A3(n_1163),
.B(n_990),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1034),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1060),
.A2(n_856),
.A3(n_1163),
.B(n_990),
.Y(n_1255)
);

O2A1O1Ixp5_ASAP7_75t_L g1256 ( 
.A1(n_1060),
.A2(n_984),
.B(n_1081),
.C(n_1080),
.Y(n_1256)
);

AO21x1_ASAP7_75t_L g1257 ( 
.A1(n_1182),
.A2(n_1060),
.B(n_1062),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1062),
.A2(n_984),
.B1(n_1169),
.B2(n_966),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1062),
.A2(n_984),
.B1(n_1169),
.B2(n_966),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_SL g1260 ( 
.A1(n_1182),
.A2(n_1183),
.B(n_1178),
.C(n_1172),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1062),
.B(n_1169),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1262)
);

CKINVDCx6p67_ASAP7_75t_R g1263 ( 
.A(n_1036),
.Y(n_1263)
);

OAI22x1_ASAP7_75t_L g1264 ( 
.A1(n_1106),
.A2(n_523),
.B1(n_725),
.B2(n_966),
.Y(n_1264)
);

AND3x4_ASAP7_75t_L g1265 ( 
.A(n_1174),
.B(n_748),
.C(n_522),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1080),
.A2(n_1081),
.B(n_1146),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_1124),
.B(n_1141),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_SL g1273 ( 
.A1(n_1182),
.A2(n_1183),
.B(n_1178),
.C(n_1172),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1178),
.B(n_536),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1060),
.A2(n_856),
.A3(n_1163),
.B(n_990),
.Y(n_1276)
);

BUFx4f_ASAP7_75t_L g1277 ( 
.A(n_1034),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1040),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1091),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1178),
.B(n_536),
.Y(n_1282)
);

NOR2xp67_ASAP7_75t_SL g1283 ( 
.A(n_1036),
.B(n_536),
.Y(n_1283)
);

NOR4xp25_ASAP7_75t_L g1284 ( 
.A(n_1182),
.B(n_921),
.C(n_1103),
.D(n_962),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1042),
.B(n_673),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1040),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1042),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1182),
.A2(n_921),
.B(n_1109),
.Y(n_1289)
);

NAND3x1_ASAP7_75t_L g1290 ( 
.A(n_1178),
.B(n_984),
.C(n_962),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1039),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1080),
.A2(n_1081),
.B(n_1146),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1040),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1183),
.C(n_1178),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1089),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1042),
.Y(n_1302)
);

OAI22x1_ASAP7_75t_L g1303 ( 
.A1(n_1106),
.A2(n_523),
.B1(n_725),
.B2(n_966),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1034),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1062),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1183),
.C(n_1178),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1182),
.A2(n_984),
.B(n_1183),
.C(n_1178),
.Y(n_1307)
);

AOI211x1_ASAP7_75t_L g1308 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1183),
.C(n_1178),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1162),
.A2(n_1143),
.B(n_1118),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1062),
.A2(n_1178),
.B1(n_1183),
.B2(n_1106),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1040),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1042),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1042),
.B(n_673),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1040),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1042),
.B(n_549),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1040),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1040),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1040),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1182),
.A2(n_984),
.B(n_900),
.C(n_998),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1040),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1062),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1182),
.A2(n_1105),
.B(n_1172),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_SL g1327 ( 
.A1(n_1182),
.A2(n_1081),
.B(n_1080),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1264),
.A2(n_1303),
.B1(n_1195),
.B2(n_1259),
.Y(n_1328)
);

BUFx4f_ASAP7_75t_L g1329 ( 
.A(n_1263),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1258),
.A2(n_1259),
.B1(n_1261),
.B2(n_1224),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1261),
.A2(n_1188),
.B1(n_1327),
.B2(n_1198),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1274),
.A2(n_1282),
.B1(n_1258),
.B2(n_1312),
.Y(n_1332)
);

BUFx4_ASAP7_75t_R g1333 ( 
.A(n_1233),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1277),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1265),
.A2(n_1281),
.B1(n_1187),
.B2(n_1188),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1252),
.Y(n_1336)
);

BUFx12f_ASAP7_75t_L g1337 ( 
.A(n_1222),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1285),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1185),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1198),
.A2(n_1200),
.B1(n_1257),
.B2(n_1305),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1238),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1248),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1200),
.A2(n_1325),
.B1(n_1289),
.B2(n_1249),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1249),
.A2(n_1289),
.B1(n_1295),
.B2(n_1266),
.Y(n_1344)
);

BUFx8_ASAP7_75t_L g1345 ( 
.A(n_1245),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1266),
.A2(n_1295),
.B1(n_1287),
.B2(n_1278),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1184),
.A2(n_1301),
.B1(n_1291),
.B2(n_1250),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1311),
.B(n_1317),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1323),
.A2(n_1290),
.B1(n_1186),
.B2(n_1194),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1302),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1279),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1211),
.B(n_1297),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1286),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1288),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1306),
.A2(n_1307),
.B1(n_1308),
.B2(n_1314),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1315),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1190),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1319),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1296),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1277),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1210),
.B(n_1215),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1228),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1256),
.A2(n_1191),
.B(n_1192),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1223),
.A2(n_1234),
.B1(n_1243),
.B2(n_1294),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1231),
.A2(n_1233),
.B1(n_1214),
.B2(n_1324),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1190),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1221),
.A2(n_1214),
.B1(n_1313),
.B2(n_1318),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1251),
.A2(n_1326),
.B(n_1316),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1231),
.A2(n_1196),
.B(n_1197),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1244),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1254),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1283),
.A2(n_1246),
.B1(n_1232),
.B2(n_1284),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1320),
.A2(n_1322),
.B1(n_1321),
.B2(n_1193),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1219),
.Y(n_1374)
);

INVx6_ASAP7_75t_L g1375 ( 
.A(n_1254),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1212),
.A2(n_1197),
.B1(n_1284),
.B2(n_1209),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1230),
.A2(n_1208),
.B1(n_1309),
.B2(n_1300),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1217),
.Y(n_1378)
);

BUFx4f_ASAP7_75t_L g1379 ( 
.A(n_1298),
.Y(n_1379)
);

BUFx8_ASAP7_75t_L g1380 ( 
.A(n_1241),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1216),
.A2(n_1220),
.B1(n_1270),
.B2(n_1293),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1268),
.A2(n_1269),
.B1(n_1272),
.B2(n_1239),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1247),
.A2(n_1260),
.B(n_1273),
.Y(n_1383)
);

BUFx4f_ASAP7_75t_SL g1384 ( 
.A(n_1237),
.Y(n_1384)
);

BUFx8_ASAP7_75t_L g1385 ( 
.A(n_1247),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1232),
.A2(n_1267),
.B1(n_1235),
.B2(n_1225),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1226),
.A2(n_1229),
.B1(n_1236),
.B2(n_1267),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1236),
.A2(n_1229),
.B1(n_1240),
.B2(n_1204),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1226),
.A2(n_1206),
.B1(n_1199),
.B2(n_1203),
.Y(n_1389)
);

BUFx4_ASAP7_75t_R g1390 ( 
.A(n_1242),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1213),
.A2(n_1242),
.B1(n_1206),
.B2(n_1207),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1205),
.A2(n_1276),
.B1(n_1255),
.B2(n_1253),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1205),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1227),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1218),
.A2(n_1202),
.B1(n_1310),
.B2(n_1189),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1218),
.A2(n_1276),
.B1(n_1253),
.B2(n_1255),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1201),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1262),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1271),
.A2(n_1275),
.B1(n_1280),
.B2(n_1292),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1299),
.A2(n_1258),
.B1(n_1259),
.B2(n_1323),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1264),
.A2(n_966),
.B1(n_1303),
.B2(n_523),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1267),
.B(n_1304),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1195),
.A2(n_1274),
.B1(n_1282),
.B2(n_984),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1264),
.A2(n_966),
.B1(n_1303),
.B2(n_523),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1264),
.A2(n_966),
.B1(n_1303),
.B2(n_523),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1288),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1238),
.Y(n_1407)
);

BUFx4_ASAP7_75t_R g1408 ( 
.A(n_1233),
.Y(n_1408)
);

BUFx4_ASAP7_75t_SL g1409 ( 
.A(n_1281),
.Y(n_1409)
);

BUFx10_ASAP7_75t_L g1410 ( 
.A(n_1241),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1195),
.A2(n_966),
.B1(n_523),
.B2(n_1264),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1195),
.A2(n_966),
.B1(n_523),
.B2(n_1264),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1302),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1185),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1302),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1187),
.B(n_1184),
.Y(n_1416)
);

BUFx4_ASAP7_75t_SL g1417 ( 
.A(n_1281),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1187),
.B(n_1184),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1288),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1195),
.A2(n_966),
.B1(n_523),
.B2(n_1264),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1264),
.A2(n_966),
.B1(n_1303),
.B2(n_523),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1302),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1302),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1261),
.A2(n_1062),
.B1(n_1169),
.B2(n_966),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1281),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1261),
.A2(n_1062),
.B1(n_1169),
.B2(n_966),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1195),
.A2(n_966),
.B1(n_523),
.B2(n_1264),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1261),
.A2(n_1062),
.B1(n_1169),
.B2(n_966),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1195),
.A2(n_966),
.B1(n_523),
.B2(n_1264),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1277),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1261),
.A2(n_1062),
.B1(n_1169),
.B2(n_966),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1281),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1195),
.A2(n_966),
.B1(n_523),
.B2(n_1264),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1195),
.A2(n_1274),
.B1(n_1282),
.B2(n_984),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1222),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1258),
.A2(n_1259),
.B1(n_1323),
.B2(n_984),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1185),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1363),
.A2(n_1368),
.B(n_1391),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1384),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1397),
.Y(n_1440)
);

AOI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1368),
.A2(n_1363),
.B(n_1377),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1347),
.B(n_1352),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1344),
.B(n_1339),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1398),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1389),
.A2(n_1395),
.B(n_1346),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1384),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1344),
.B(n_1342),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1436),
.A2(n_1349),
.B(n_1403),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1425),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1394),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1437),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1351),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1353),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1359),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1389),
.A2(n_1395),
.B(n_1346),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1434),
.A2(n_1332),
.B1(n_1331),
.B2(n_1424),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1414),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1385),
.A2(n_1426),
.B1(n_1424),
.B2(n_1431),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1392),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1347),
.B(n_1376),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1396),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1406),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1422),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1382),
.A2(n_1381),
.B(n_1365),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1396),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1331),
.B(n_1376),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1400),
.A2(n_1388),
.B(n_1383),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1369),
.A2(n_1340),
.B(n_1387),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1343),
.B(n_1406),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1343),
.B(n_1419),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1432),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1385),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1419),
.B(n_1354),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1370),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1382),
.A2(n_1381),
.B(n_1365),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1373),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1390),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1393),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1330),
.B(n_1328),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1364),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1355),
.A2(n_1361),
.B(n_1418),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1386),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1367),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1367),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1372),
.A2(n_1348),
.B(n_1416),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1336),
.B(n_1338),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1387),
.A2(n_1328),
.B(n_1402),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1399),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1426),
.A2(n_1428),
.B(n_1431),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1413),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1415),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1409),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1428),
.B(n_1362),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1335),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1356),
.B(n_1423),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1420),
.B(n_1427),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1374),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1410),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1350),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1358),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1410),
.Y(n_1502)
);

AO21x1_ASAP7_75t_L g1503 ( 
.A1(n_1334),
.A2(n_1433),
.B(n_1429),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1401),
.B(n_1421),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1492),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1462),
.B(n_1378),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_SL g1507 ( 
.A1(n_1448),
.A2(n_1409),
.B(n_1417),
.C(n_1333),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1442),
.B(n_1357),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1449),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1442),
.B(n_1405),
.Y(n_1510)
);

NAND4xp25_ASAP7_75t_L g1511 ( 
.A(n_1448),
.B(n_1421),
.C(n_1404),
.D(n_1401),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1366),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1463),
.B(n_1341),
.Y(n_1513)
);

AOI211xp5_ASAP7_75t_L g1514 ( 
.A1(n_1456),
.A2(n_1360),
.B(n_1430),
.C(n_1408),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1494),
.A2(n_1379),
.B1(n_1329),
.B2(n_1430),
.C(n_1360),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1471),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1463),
.B(n_1329),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1473),
.B(n_1375),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1494),
.A2(n_1337),
.B1(n_1435),
.B2(n_1371),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1485),
.B(n_1380),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1452),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1380),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1499),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1443),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1462),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1438),
.A2(n_1345),
.B(n_1417),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1460),
.A2(n_1407),
.B(n_1466),
.C(n_1479),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1471),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1473),
.B(n_1407),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1495),
.B(n_1491),
.Y(n_1530)
);

BUFx8_ASAP7_75t_L g1531 ( 
.A(n_1471),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1474),
.B(n_1486),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1500),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_SL g1534 ( 
.A1(n_1468),
.A2(n_1503),
.B(n_1502),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1439),
.B(n_1446),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1438),
.A2(n_1467),
.B(n_1488),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1495),
.B(n_1491),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1440),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1466),
.A2(n_1479),
.B1(n_1503),
.B2(n_1468),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1485),
.B(n_1443),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1439),
.B(n_1446),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1467),
.A2(n_1468),
.B(n_1482),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1453),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1488),
.A2(n_1441),
.B(n_1450),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1490),
.B(n_1469),
.Y(n_1545)
);

CKINVDCx8_ASAP7_75t_R g1546 ( 
.A(n_1500),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1468),
.A2(n_1504),
.B1(n_1489),
.B2(n_1458),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1469),
.B(n_1470),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1470),
.B(n_1447),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1499),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1499),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1504),
.A2(n_1483),
.B1(n_1446),
.B2(n_1439),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1483),
.A2(n_1504),
.B(n_1487),
.C(n_1496),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1447),
.B(n_1498),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1498),
.B(n_1502),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1489),
.A2(n_1475),
.B1(n_1464),
.B2(n_1484),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1438),
.A2(n_1487),
.B(n_1441),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1497),
.A2(n_1475),
.B(n_1464),
.C(n_1496),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_L g1559 ( 
.A1(n_1497),
.A2(n_1484),
.B(n_1461),
.C(n_1465),
.Y(n_1559)
);

AND2x6_ASAP7_75t_L g1560 ( 
.A(n_1472),
.B(n_1477),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1489),
.A2(n_1475),
.B1(n_1464),
.B2(n_1493),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1536),
.B(n_1475),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1445),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1512),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1548),
.B(n_1445),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1549),
.B(n_1445),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1557),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1543),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1557),
.B(n_1445),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1545),
.B(n_1445),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1531),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1444),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1511),
.A2(n_1489),
.B1(n_1461),
.B2(n_1465),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1544),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1554),
.B(n_1455),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1561),
.B(n_1455),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1512),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1539),
.A2(n_1493),
.B1(n_1476),
.B2(n_1472),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1544),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1526),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1530),
.B(n_1455),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1538),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1525),
.B(n_1459),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1537),
.B(n_1455),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1538),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1547),
.A2(n_1476),
.B1(n_1493),
.B2(n_1480),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1542),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1455),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1524),
.B(n_1540),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1560),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1524),
.B(n_1459),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1592),
.B(n_1525),
.Y(n_1593)
);

AND2x2_ASAP7_75t_SL g1594 ( 
.A(n_1562),
.B(n_1540),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1564),
.Y(n_1596)
);

AOI33xp33_ASAP7_75t_L g1597 ( 
.A1(n_1574),
.A2(n_1556),
.A3(n_1558),
.B1(n_1555),
.B2(n_1454),
.B3(n_1457),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1572),
.B(n_1509),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_1570),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1572),
.Y(n_1600)
);

AOI211xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1565),
.A2(n_1507),
.B(n_1552),
.C(n_1541),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1586),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1574),
.A2(n_1510),
.B1(n_1553),
.B2(n_1559),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1569),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1592),
.B(n_1532),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1583),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1591),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1592),
.B(n_1558),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1586),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1582),
.B(n_1523),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1575),
.A2(n_1534),
.B(n_1520),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1586),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1582),
.B(n_1518),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1564),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1583),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1577),
.A2(n_1478),
.B1(n_1477),
.B2(n_1480),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1584),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.B(n_1552),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1451),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1451),
.Y(n_1621)
);

OAI31xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1577),
.A2(n_1508),
.A3(n_1522),
.B(n_1541),
.Y(n_1622)
);

AOI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1562),
.A2(n_1508),
.B(n_1527),
.C(n_1510),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1506),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1570),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1572),
.Y(n_1626)
);

NAND4xp25_ASAP7_75t_L g1627 ( 
.A(n_1562),
.B(n_1514),
.C(n_1522),
.D(n_1535),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_1551),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1570),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1628),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1599),
.B(n_1585),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_1588),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1593),
.B(n_1590),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1628),
.B(n_1611),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1585),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1602),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1595),
.B(n_1591),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1611),
.B(n_1585),
.Y(n_1640)
);

AND2x4_ASAP7_75t_SL g1641 ( 
.A(n_1600),
.B(n_1573),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1602),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1571),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1621),
.B(n_1571),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1593),
.B(n_1619),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1621),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1603),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1620),
.Y(n_1648)
);

BUFx4f_ASAP7_75t_L g1649 ( 
.A(n_1600),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1620),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1607),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1608),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1605),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1614),
.B(n_1571),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1625),
.B(n_1571),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1625),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1563),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1565),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1629),
.B(n_1576),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1595),
.B(n_1591),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1629),
.B(n_1576),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1619),
.B(n_1566),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1596),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1616),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1641),
.B(n_1624),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1664),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1656),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1657),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1658),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1664),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1645),
.B(n_1606),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1657),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1641),
.B(n_1643),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1656),
.Y(n_1674)
);

AND2x2_ASAP7_75t_SL g1675 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1656),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1641),
.B(n_1591),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1651),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1633),
.A2(n_1604),
.B1(n_1577),
.B2(n_1589),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1658),
.B(n_1600),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1651),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1645),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1633),
.B(n_1622),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1645),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1634),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1634),
.B(n_1603),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1648),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1638),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1648),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1656),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1634),
.B(n_1610),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1650),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1647),
.B(n_1613),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1647),
.B(n_1613),
.Y(n_1697)
);

NOR2xp67_ASAP7_75t_SL g1698 ( 
.A(n_1652),
.B(n_1572),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.B(n_1606),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1641),
.B(n_1601),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1656),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1635),
.B(n_1601),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1635),
.Y(n_1704)
);

NOR2x1_ASAP7_75t_SL g1705 ( 
.A(n_1662),
.B(n_1626),
.Y(n_1705)
);

NAND2x2_ASAP7_75t_L g1706 ( 
.A(n_1635),
.B(n_1505),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1632),
.B(n_1596),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1688),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1688),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1652),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1675),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_1699),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1703),
.A2(n_1652),
.B(n_1546),
.C(n_1623),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1702),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1671),
.B(n_1632),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1675),
.B(n_1643),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1682),
.B(n_1646),
.Y(n_1717)
);

NAND2x1_ASAP7_75t_L g1718 ( 
.A(n_1700),
.B(n_1639),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1679),
.B(n_1631),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1704),
.B(n_1631),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1705),
.B(n_1643),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1666),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1670),
.B(n_1631),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1669),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1705),
.B(n_1626),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1700),
.B(n_1673),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1677),
.B(n_1649),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1687),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1699),
.B(n_1644),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1673),
.B(n_1654),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_L g1733 ( 
.A(n_1686),
.B(n_1626),
.C(n_1519),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1678),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1698),
.B(n_1626),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1689),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1667),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1681),
.B(n_1672),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1668),
.B(n_1685),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1668),
.B(n_1644),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1667),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1694),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1711),
.A2(n_1516),
.B1(n_1528),
.B2(n_1598),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1725),
.B(n_1698),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1716),
.A2(n_1711),
.B(n_1720),
.Y(n_1747)
);

XNOR2x2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.B(n_1686),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1716),
.B(n_1677),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1680),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1727),
.B(n_1665),
.Y(n_1751)
);

AOI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1713),
.A2(n_1695),
.B(n_1707),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1712),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1712),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1665),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1708),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1733),
.A2(n_1597),
.B(n_1623),
.C(n_1604),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1726),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1718),
.A2(n_1693),
.B(n_1726),
.Y(n_1759)
);

OAI311xp33_ASAP7_75t_L g1760 ( 
.A1(n_1739),
.A2(n_1697),
.A3(n_1696),
.B1(n_1691),
.C1(n_1627),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1708),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1709),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1715),
.B(n_1707),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_SL g1764 ( 
.A(n_1718),
.B(n_1693),
.C(n_1578),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1726),
.B(n_1654),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1709),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1729),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1735),
.A2(n_1562),
.B(n_1578),
.C(n_1579),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1729),
.A2(n_1570),
.B1(n_1615),
.B2(n_1589),
.C(n_1663),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1734),
.B(n_1640),
.Y(n_1770)
);

NAND3xp33_ASAP7_75t_L g1771 ( 
.A(n_1757),
.B(n_1723),
.C(n_1739),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1748),
.A2(n_1589),
.B1(n_1732),
.B2(n_1714),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1751),
.B(n_1755),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1757),
.A2(n_1706),
.B1(n_1722),
.B2(n_1728),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1754),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1754),
.B(n_1723),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1753),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1748),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1746),
.Y(n_1779)
);

OAI32xp33_ASAP7_75t_L g1780 ( 
.A1(n_1747),
.A2(n_1738),
.A3(n_1715),
.B1(n_1736),
.B2(n_1744),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1751),
.B(n_1714),
.Y(n_1781)
);

OAI21xp33_ASAP7_75t_SL g1782 ( 
.A1(n_1759),
.A2(n_1722),
.B(n_1743),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1764),
.B(n_1736),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1755),
.B(n_1743),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1749),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1760),
.A2(n_1744),
.B1(n_1732),
.B2(n_1719),
.C(n_1717),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1756),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1750),
.B(n_1731),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1752),
.A2(n_1724),
.B(n_1738),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1778),
.Y(n_1791)
);

NOR2xp67_ASAP7_75t_L g1792 ( 
.A(n_1773),
.B(n_1763),
.Y(n_1792)
);

OAI322xp33_ASAP7_75t_L g1793 ( 
.A1(n_1771),
.A2(n_1763),
.A3(n_1758),
.B1(n_1767),
.B2(n_1766),
.C1(n_1761),
.C2(n_1762),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1772),
.A2(n_1768),
.B1(n_1769),
.B2(n_1745),
.C(n_1750),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1773),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1789),
.B(n_1765),
.Y(n_1796)
);

AOI211x1_ASAP7_75t_L g1797 ( 
.A1(n_1780),
.A2(n_1770),
.B(n_1765),
.C(n_1721),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1780),
.A2(n_1768),
.B(n_1742),
.C(n_1737),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1785),
.Y(n_1799)
);

OAI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1783),
.A2(n_1706),
.B1(n_1741),
.B2(n_1730),
.C(n_1740),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1789),
.B(n_1730),
.Y(n_1801)
);

AOI31xp33_ASAP7_75t_L g1802 ( 
.A1(n_1779),
.A2(n_1775),
.A3(n_1777),
.B(n_1774),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1792),
.B(n_1786),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1798),
.A2(n_1790),
.B(n_1787),
.Y(n_1804)
);

NAND4xp25_ASAP7_75t_L g1805 ( 
.A(n_1797),
.B(n_1786),
.C(n_1781),
.D(n_1785),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1799),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1795),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_L g1808 ( 
.A(n_1791),
.B(n_1776),
.C(n_1775),
.Y(n_1808)
);

NAND4xp25_ASAP7_75t_L g1809 ( 
.A(n_1800),
.B(n_1796),
.C(n_1801),
.D(n_1794),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1802),
.B(n_1784),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1793),
.B(n_1784),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1802),
.B(n_1788),
.Y(n_1812)
);

AOI211xp5_ASAP7_75t_L g1813 ( 
.A1(n_1804),
.A2(n_1782),
.B(n_1519),
.C(n_1737),
.Y(n_1813)
);

CKINVDCx16_ASAP7_75t_R g1814 ( 
.A(n_1810),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1811),
.A2(n_1812),
.B1(n_1806),
.B2(n_1803),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1807),
.Y(n_1816)
);

OAI321xp33_ASAP7_75t_L g1817 ( 
.A1(n_1809),
.A2(n_1742),
.A3(n_1627),
.B1(n_1741),
.B2(n_1740),
.C(n_1579),
.Y(n_1817)
);

AOI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1808),
.A2(n_1615),
.B1(n_1568),
.B2(n_1676),
.C(n_1674),
.Y(n_1818)
);

OAI211xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1805),
.A2(n_1701),
.B(n_1692),
.C(n_1676),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1816),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1815),
.A2(n_1649),
.B(n_1674),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1814),
.Y(n_1822)
);

OAI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1817),
.A2(n_1813),
.B1(n_1819),
.B2(n_1818),
.C1(n_1579),
.C2(n_1692),
.Y(n_1823)
);

AOI322xp5_ASAP7_75t_L g1824 ( 
.A1(n_1814),
.A2(n_1594),
.A3(n_1589),
.B1(n_1587),
.B2(n_1567),
.C1(n_1566),
.C2(n_1617),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1814),
.A2(n_1580),
.B1(n_1575),
.B2(n_1612),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1822),
.B(n_1701),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1820),
.A2(n_1649),
.B(n_1531),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1821),
.B(n_1630),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1823),
.B(n_1529),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1825),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1829),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1830),
.A2(n_1824),
.B1(n_1663),
.B2(n_1568),
.C(n_1649),
.Y(n_1832)
);

OR4x1_ASAP7_75t_L g1833 ( 
.A(n_1826),
.B(n_1550),
.C(n_1581),
.D(n_1653),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1831),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1834),
.Y(n_1835)
);

AND2x2_ASAP7_75t_SL g1836 ( 
.A(n_1835),
.B(n_1828),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1835),
.A2(n_1833),
.B1(n_1827),
.B2(n_1832),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1663),
.B1(n_1533),
.B2(n_1630),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1837),
.A2(n_1515),
.B1(n_1581),
.B2(n_1660),
.Y(n_1839)
);

OAI21x1_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1630),
.B(n_1636),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1839),
.Y(n_1841)
);

XNOR2xp5_ASAP7_75t_L g1842 ( 
.A(n_1841),
.B(n_1501),
.Y(n_1842)
);

OA21x2_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1840),
.B(n_1636),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1661),
.B1(n_1655),
.B2(n_1659),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1642),
.B1(n_1638),
.B2(n_1653),
.C(n_1639),
.Y(n_1845)
);

AOI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1515),
.B(n_1513),
.C(n_1517),
.Y(n_1846)
);


endmodule