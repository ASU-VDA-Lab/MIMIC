module real_jpeg_27846_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_0),
.A2(n_24),
.B1(n_52),
.B2(n_53),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_0),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_24),
.B1(n_58),
.B2(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_60),
.Y(n_95)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_47),
.B1(n_58),
.B2(n_60),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_47),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_4),
.A2(n_26),
.B1(n_30),
.B2(n_174),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_174),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_4),
.A2(n_58),
.B1(n_60),
.B2(n_174),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_6),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_25),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_30),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_6),
.A2(n_30),
.B(n_212),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_172),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_6),
.A2(n_11),
.B(n_58),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_78),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_6),
.A2(n_100),
.B1(n_118),
.B2(n_260),
.Y(n_262)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_26),
.B1(n_30),
.B2(n_45),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_45),
.B1(n_58),
.B2(n_60),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_114),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_114),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_9),
.A2(n_58),
.B1(n_60),
.B2(n_114),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_10),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_139),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_139),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_10),
.A2(n_58),
.B1(n_60),
.B2(n_139),
.Y(n_252)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_12),
.A2(n_36),
.B1(n_58),
.B2(n_60),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_122)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_85),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_83),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_20),
.A2(n_43),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_21),
.A2(n_32),
.B(n_82),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_25),
.B(n_28),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_28),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_22),
.B(n_172),
.CON(n_171),
.SN(n_171)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_25),
.A2(n_32),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_26),
.A2(n_30),
.B1(n_67),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_26),
.A2(n_33),
.B1(n_171),
.B2(n_185),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g210 ( 
.A1(n_26),
.A2(n_52),
.A3(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_28),
.B(n_30),
.Y(n_185)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_31),
.A2(n_44),
.B(n_48),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_32),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_48),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_75),
.C(n_80),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_39),
.A2(n_40),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.C(n_63),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_41),
.A2(n_42),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_43),
.A2(n_48),
.B1(n_113),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_43),
.A2(n_48),
.B1(n_138),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_49),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_49),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_49),
.A2(n_63),
.B1(n_309),
.B2(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_61),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_57),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_50),
.A2(n_106),
.B(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_50),
.A2(n_61),
.B(n_121),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_50),
.A2(n_57),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_50),
.A2(n_145),
.B(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_50),
.A2(n_57),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_50),
.A2(n_57),
.B1(n_219),
.B2(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_53),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_53),
.B(n_74),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_53),
.A2(n_56),
.B(n_172),
.C(n_239),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_105),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_57),
.B(n_172),
.Y(n_258)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_60),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_62),
.B(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_63),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_64),
.A2(n_77),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_65),
.A2(n_72),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_65),
.A2(n_72),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_65),
.A2(n_72),
.B1(n_168),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_65),
.A2(n_72),
.B1(n_197),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_78),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_79),
.B(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_77),
.A2(n_135),
.B(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_80),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_334),
.B(n_340),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_304),
.A3(n_326),
.B1(n_332),
.B2(n_333),
.C(n_342),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_157),
.B(n_303),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_140),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_89),
.B(n_140),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_115),
.C(n_125),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_90),
.A2(n_91),
.B1(n_115),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_107),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_109),
.C(n_111),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_93),
.B(n_104),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_94),
.A2(n_187),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_95),
.A2(n_103),
.B(n_130),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_95),
.A2(n_99),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_98),
.A2(n_118),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_101),
.Y(n_188)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_102),
.A2(n_118),
.B1(n_252),
.B2(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_102),
.B(n_172),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_115),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_124),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_117),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_120),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_117),
.A2(n_151),
.B(n_154),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_118),
.A2(n_128),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_125),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_134),
.C(n_136),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_126),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_131),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_134),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_155),
.B2(n_156),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_143),
.B(n_150),
.C(n_156),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B(n_149),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_149),
.B(n_306),
.C(n_316),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_149),
.A2(n_306),
.B1(n_307),
.B2(n_331),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_149),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_155),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_297),
.B(n_302),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_202),
.B(n_283),
.C(n_296),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_189),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_160),
.B(n_189),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_175),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_162),
.B(n_163),
.C(n_175),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_170),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_177),
.B(n_181),
.C(n_183),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_190),
.A2(n_191),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_282),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_275),
.B(n_281),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_230),
.B(n_274),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_221),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_206),
.B(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.C(n_217),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_207),
.A2(n_208),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_210),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_228),
.C(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_268),
.B(n_273),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_248),
.B(n_267),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_256),
.B(n_266),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_294),
.B2(n_295),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_318),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_318),
.Y(n_333)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_311),
.C(n_313),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_315),
.B1(n_320),
.B2(n_324),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_324),
.C(n_325),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_316),
.A2(n_317),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_337),
.Y(n_339)
);


endmodule