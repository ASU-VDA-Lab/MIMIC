module fake_jpeg_31460_n_369 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_369);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_369;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_54),
.A2(n_14),
.B(n_13),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_72),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_99),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_62),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_32),
.B1(n_34),
.B2(n_31),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_41),
.B1(n_25),
.B2(n_31),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_29),
.B1(n_28),
.B2(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_24),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_34),
.B1(n_26),
.B2(n_27),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_24),
.B1(n_19),
.B2(n_26),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_118),
.B1(n_47),
.B2(n_51),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_27),
.B(n_37),
.C(n_29),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_30),
.B(n_12),
.C(n_3),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_29),
.B1(n_28),
.B2(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_37),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_124),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_29),
.B1(n_28),
.B2(n_23),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_29),
.B1(n_28),
.B2(n_38),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_38),
.B1(n_17),
.B2(n_9),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_123),
.B1(n_0),
.B2(n_4),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_17),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_130),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_10),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_128),
.B(n_129),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_90),
.B(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_138),
.Y(n_186)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

NAND2x1p5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_62),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_9),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_80),
.A2(n_17),
.B1(n_47),
.B2(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_148),
.B1(n_152),
.B2(n_158),
.Y(n_168)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_159),
.B1(n_96),
.B2(n_105),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_17),
.B1(n_77),
.B2(n_30),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_151),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_98),
.A2(n_30),
.B1(n_12),
.B2(n_2),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_81),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_84),
.B(n_0),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_153),
.Y(n_198)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_30),
.B1(n_1),
.B2(n_3),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_157),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_98),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_162),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_7),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_4),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_119),
.C(n_91),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_166),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_82),
.A2(n_6),
.B(n_7),
.C(n_85),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_87),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_6),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_202),
.B(n_151),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_190),
.B1(n_191),
.B2(n_195),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_198),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_82),
.B(n_107),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_176),
.A2(n_135),
.B(n_131),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_134),
.A2(n_146),
.B1(n_100),
.B2(n_111),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_163),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_121),
.B1(n_117),
.B2(n_101),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_121),
.B1(n_117),
.B2(n_101),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_150),
.A2(n_119),
.B1(n_111),
.B2(n_109),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_95),
.B1(n_93),
.B2(n_109),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_196),
.A2(n_203),
.B1(n_158),
.B2(n_146),
.Y(n_222)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_134),
.B(n_105),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_142),
.A2(n_95),
.B1(n_105),
.B2(n_94),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_208),
.B(n_209),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_126),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_214),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_150),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_132),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_216),
.B(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_126),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_137),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_128),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_223),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_233),
.B1(n_238),
.B2(n_197),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_125),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_229),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_165),
.B(n_160),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_230),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_141),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_231),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_133),
.C(n_146),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_234),
.C(n_183),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_194),
.Y(n_229)
);

A2O1A1O1Ixp25_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_155),
.B(n_157),
.C(n_139),
.D(n_149),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_170),
.B(n_155),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_193),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_173),
.A2(n_155),
.B1(n_164),
.B2(n_161),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_202),
.C(n_195),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_201),
.B1(n_203),
.B2(n_196),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_186),
.B(n_157),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_174),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_244),
.B(n_252),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_171),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_177),
.C(n_201),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_234),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_232),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_263),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_201),
.A3(n_168),
.B1(n_157),
.B2(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_178),
.C(n_185),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_192),
.C(n_178),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_192),
.C(n_197),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_223),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_264),
.B(n_253),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_267),
.B1(n_229),
.B2(n_220),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_220),
.A2(n_136),
.B1(n_156),
.B2(n_182),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_206),
.A2(n_180),
.B1(n_169),
.B2(n_199),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_198),
.B1(n_180),
.B2(n_235),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_208),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_274),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_209),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_241),
.A2(n_239),
.B(n_228),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_282),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_273),
.B1(n_265),
.B2(n_259),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_233),
.B1(n_238),
.B2(n_222),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_216),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_286),
.B(n_287),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_291),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_225),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_217),
.C(n_226),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_260),
.C(n_266),
.Y(n_298)
);

BUFx12_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_236),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_296),
.A2(n_299),
.B1(n_313),
.B2(n_230),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_305),
.C(n_312),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_249),
.B1(n_252),
.B2(n_266),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_256),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_304),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_311),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_248),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_262),
.C(n_261),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_276),
.B(n_253),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_258),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_243),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_243),
.C(n_211),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_281),
.A2(n_282),
.B1(n_272),
.B2(n_275),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_274),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_318),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_317),
.B(n_320),
.Y(n_335)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_322),
.Y(n_341)
);

OAI322xp33_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_292),
.A3(n_295),
.B1(n_293),
.B2(n_246),
.C1(n_242),
.C2(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_297),
.B(n_247),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_302),
.C(n_305),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_313),
.B1(n_296),
.B2(n_299),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_289),
.C(n_280),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_288),
.C(n_285),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_283),
.C(n_294),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_174),
.C(n_189),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_332),
.B1(n_334),
.B2(n_337),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_301),
.B(n_294),
.C(n_308),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_87),
.B(n_145),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_301),
.B1(n_309),
.B2(n_314),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_270),
.B1(n_312),
.B2(n_254),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_294),
.B1(n_240),
.B2(n_237),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_237),
.B1(n_188),
.B2(n_169),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_338),
.B(n_145),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_321),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_189),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_340),
.B(n_329),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_326),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_348),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_315),
.B(n_328),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_347),
.B(n_331),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_345),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_335),
.A2(n_321),
.B(n_323),
.Y(n_346)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_346),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_336),
.B(n_154),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_334),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_332),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_354),
.B(n_355),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_337),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_356),
.B(n_358),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_347),
.A2(n_331),
.B(n_330),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_351),
.A2(n_344),
.B(n_340),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_361),
.A2(n_357),
.B(n_359),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_353),
.B(n_352),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_362),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_363),
.B(n_365),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_284),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_366),
.Y(n_367)
);

NAND2x1_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_364),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_365),
.Y(n_369)
);


endmodule