module fake_jpeg_8136_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_20;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_21),
.B1(n_30),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_54),
.B1(n_41),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_30),
.B2(n_39),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_24),
.B(n_30),
.C(n_21),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_35),
.B(n_34),
.C(n_19),
.Y(n_83)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_17),
.B1(n_38),
.B2(n_36),
.Y(n_81)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_89),
.B1(n_61),
.B2(n_37),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_38),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_77),
.B(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_34),
.CI(n_35),
.CON(n_76),
.SN(n_76)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_87),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_36),
.B(n_46),
.C(n_16),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_38),
.B1(n_29),
.B2(n_19),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_84),
.B(n_90),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_34),
.B(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp67_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_17),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_55),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_97),
.B(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_110),
.B1(n_112),
.B2(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_51),
.B1(n_37),
.B2(n_39),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_100),
.B1(n_108),
.B2(n_116),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_35),
.A3(n_42),
.B1(n_39),
.B2(n_37),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_106),
.Y(n_131)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_55),
.B1(n_35),
.B2(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_39),
.B1(n_37),
.B2(n_42),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_47),
.B1(n_59),
.B2(n_34),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_57),
.B1(n_48),
.B2(n_44),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_36),
.B1(n_65),
.B2(n_45),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_78),
.B1(n_33),
.B2(n_28),
.Y(n_145)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_46),
.B1(n_44),
.B2(n_31),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_74),
.B1(n_85),
.B2(n_100),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_91),
.B1(n_70),
.B2(n_71),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_136),
.B1(n_140),
.B2(n_114),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_76),
.B(n_27),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_136),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_88),
.C(n_91),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_99),
.C(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_13),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_128),
.Y(n_158)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_130),
.B1(n_103),
.B2(n_115),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_43),
.B(n_31),
.C(n_28),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_14),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_74),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_71),
.B1(n_70),
.B2(n_66),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_27),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_0),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_116),
.B(n_95),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_96),
.A2(n_66),
.B1(n_78),
.B2(n_49),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_144),
.B1(n_103),
.B2(n_98),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_93),
.A2(n_78),
.B1(n_43),
.B2(n_16),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_150),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_153),
.C(n_159),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_166),
.B1(n_168),
.B2(n_130),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_154),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_139),
.A2(n_111),
.B(n_117),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_155),
.B1(n_163),
.B2(n_15),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_102),
.C(n_98),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_171),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_27),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_28),
.B1(n_23),
.B2(n_20),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_141),
.C(n_121),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_122),
.C(n_142),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_23),
.B1(n_20),
.B2(n_27),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_134),
.B(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_0),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_184),
.B1(n_193),
.B2(n_155),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_125),
.B(n_130),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_185),
.B(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_119),
.B1(n_125),
.B2(n_126),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_188),
.C(n_197),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_124),
.C(n_129),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_171),
.B1(n_174),
.B2(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_18),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_154),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_18),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_18),
.C(n_1),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_199),
.C(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_18),
.C(n_1),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_169),
.B1(n_161),
.B2(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_151),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_223),
.B1(n_201),
.B2(n_181),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_150),
.B(n_175),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_205),
.C(n_209),
.Y(n_233)
);

XNOR2x2_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_165),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_146),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_212),
.C(n_214),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_158),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_163),
.B1(n_166),
.B2(n_168),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_196),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_236),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_192),
.B1(n_179),
.B2(n_189),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_235),
.B1(n_241),
.B2(n_242),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_192),
.B1(n_176),
.B2(n_200),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_207),
.C(n_212),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_207),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_176),
.B1(n_186),
.B2(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_197),
.B1(n_199),
.B2(n_188),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_216),
.B(n_213),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_247),
.B(n_253),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_251),
.C(n_231),
.Y(n_262)
);

OAI322xp33_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_217),
.A3(n_213),
.B1(n_210),
.B2(n_216),
.C1(n_209),
.C2(n_206),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_204),
.B1(n_223),
.B2(n_2),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_235),
.B1(n_234),
.B2(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_12),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_244),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_0),
.B(n_1),
.Y(n_254)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_226),
.B(n_11),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_8),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_266),
.C(n_8),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_254),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_267),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_239),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_233),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_241),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_253),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_276),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_256),
.B1(n_250),
.B2(n_242),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_277),
.C(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_251),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_246),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_262),
.C(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_287),
.C(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_6),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_265),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_279),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_9),
.C(n_3),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_291),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.C(n_292),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_284),
.B(n_5),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_284),
.B(n_5),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_295),
.B1(n_293),
.B2(n_6),
.Y(n_297)
);

AOI31xp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_6),
.A3(n_4),
.B(n_5),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_4),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_5),
.C(n_6),
.Y(n_300)
);


endmodule