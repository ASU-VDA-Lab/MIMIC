module real_jpeg_25151_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_0),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_0),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_0),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_0),
.B(n_17),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_0),
.B(n_53),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_0),
.B(n_34),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_28),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_0),
.B(n_202),
.Y(n_258)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_2),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_2),
.B(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_2),
.B(n_53),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_34),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_3),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_3),
.B(n_84),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_3),
.B(n_50),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_3),
.B(n_53),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_3),
.B(n_34),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_3),
.B(n_28),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_4),
.B(n_17),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_99),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_4),
.B(n_84),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_4),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_4),
.B(n_53),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_4),
.B(n_34),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_6),
.B(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_84),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_50),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_53),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_6),
.B(n_34),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_6),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_6),
.B(n_202),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_28),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_8),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_8),
.B(n_99),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_8),
.B(n_84),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_8),
.B(n_50),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_8),
.B(n_53),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_8),
.B(n_34),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_10),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_10),
.B(n_84),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_13),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_84),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_13),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_13),
.B(n_34),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_13),
.B(n_28),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_13),
.B(n_24),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_14),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_14),
.B(n_50),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_14),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_28),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_16),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_16),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_16),
.B(n_34),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_28),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_16),
.B(n_202),
.Y(n_241)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_17),
.Y(n_145)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_64),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_41),
.B2(n_42),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_25),
.Y(n_202)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_25),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_27),
.B(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_27),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_27),
.B(n_250),
.Y(n_344)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_29),
.B(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_29),
.B(n_238),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_61),
.C(n_62),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_43),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_43),
.B(n_389),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.CI(n_54),
.CON(n_43),
.SN(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.C(n_52),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_46),
.A2(n_47),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_48),
.A2(n_318),
.B1(n_319),
.B2(n_346),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_48),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_SL g376 ( 
.A(n_48),
.B(n_319),
.C(n_344),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_48),
.A2(n_52),
.B1(n_57),
.B2(n_346),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_49),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_49),
.B(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_58),
.C(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_53),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_59),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_61),
.B(n_62),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_388),
.C(n_390),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_383),
.C(n_384),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_365),
.C(n_366),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_336),
.C(n_337),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_311),
.C(n_312),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_279),
.C(n_280),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_243),
.C(n_244),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_208),
.C(n_209),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_175),
.C(n_176),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_150),
.C(n_151),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_110),
.C(n_122),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_91),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_77),
.B(n_86),
.C(n_91),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.C(n_82),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_79),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_87),
.B(n_89),
.C(n_90),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_92),
.B(n_102),
.C(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_99),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_109),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_121),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_115),
.B1(n_121),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_146),
.C(n_147),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.C(n_136),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_129),
.C(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_141),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_139),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_145),
.B(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_164),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_165),
.C(n_174),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_159),
.C(n_160),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_158),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_160),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.CI(n_163),
.CON(n_160),
.SN(n_160)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_174),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_172),
.B2(n_173),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_180),
.C(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_187),
.C(n_190),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_182),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.CI(n_185),
.CON(n_182),
.SN(n_182)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_184),
.C(n_185),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_199),
.C(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B1(n_206),
.B2(n_207),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_197),
.B(n_198),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_197),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_233),
.C(n_234),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_228)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_229),
.B2(n_242),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_230),
.C(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_214),
.C(n_222),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_218),
.C(n_221),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_226),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_235),
.B(n_275),
.C(n_276),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.CI(n_241),
.CON(n_235),
.SN(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_277),
.B2(n_278),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_245),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_269),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_269),
.C(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_256),
.C(n_257),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_248),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.CI(n_253),
.CON(n_248),
.SN(n_248)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_268),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_258),
.Y(n_268)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_266),
.B2(n_267),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_262),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_267),
.C(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_261),
.B(n_286),
.C(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_283),
.C(n_310),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_297),
.B2(n_310),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_292),
.C(n_293),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_290),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_SL g350 ( 
.A(n_289),
.B(n_316),
.C(n_319),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_293),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.CI(n_296),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_297),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.CI(n_300),
.CON(n_297),
.SN(n_297)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_299),
.C(n_300),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_309),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_304),
.C(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_304),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_306),
.A2(n_307),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_333),
.C(n_334),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_335),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_326),
.C(n_335),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_321),
.C(n_322),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_322),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.CI(n_325),
.CON(n_322),
.SN(n_322)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_329),
.C(n_330),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_332),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_340),
.C(n_352),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_351),
.B2(n_352),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_347),
.B2(n_348),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_349),
.C(n_350),
.Y(n_368)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_355),
.C(n_358),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_358),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_361),
.C(n_364),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_362),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_363),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_380),
.B1(n_381),
.B2(n_382),
.Y(n_366)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_369),
.C(n_382),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_376),
.C(n_377),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_385),
.C(n_387),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.CI(n_374),
.CON(n_371),
.SN(n_371)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_378),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_380),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);


endmodule