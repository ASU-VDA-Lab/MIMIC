module fake_jpeg_18343_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_55),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_58),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_44),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_35),
.B1(n_45),
.B2(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_1),
.Y(n_78)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_41),
.B1(n_38),
.B2(n_3),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_78),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_4),
.C(n_5),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_68),
.C(n_79),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_10),
.C(n_11),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_90),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_12),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_5),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_94),
.B(n_95),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_88),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_92),
.B1(n_84),
.B2(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_92),
.B1(n_81),
.B2(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_22),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_106),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_24),
.Y(n_109)
);


endmodule