module fake_jpeg_21010_n_148 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_17),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_25),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_67),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_57),
.B1(n_66),
.B2(n_74),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_48),
.B1(n_61),
.B2(n_74),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_72),
.B1(n_67),
.B2(n_52),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_79),
.B1(n_53),
.B2(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_49),
.B1(n_56),
.B2(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_68),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.C(n_102),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_69),
.B1(n_54),
.B2(n_63),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_101),
.B1(n_103),
.B2(n_0),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_79),
.B1(n_58),
.B2(n_72),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_62),
.B1(n_50),
.B2(n_60),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_88),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_111),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_26),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_117),
.B(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_22),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_27),
.B(n_42),
.C(n_41),
.D(n_40),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_123),
.B1(n_127),
.B2(n_113),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_30),
.C(n_35),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_129),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_31),
.B(n_11),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.C(n_135),
.Y(n_136)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_117),
.B1(n_120),
.B2(n_125),
.C(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_131),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_126),
.C(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_34),
.C(n_13),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_14),
.B(n_33),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g148 ( 
.A(n_147),
.Y(n_148)
);


endmodule