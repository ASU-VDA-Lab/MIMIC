module real_jpeg_24873_n_16 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_1),
.A2(n_43),
.B(n_130),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_1),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_1),
.B(n_32),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_132),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_1),
.B(n_52),
.C(n_57),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_1),
.B(n_65),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_1),
.A2(n_108),
.B1(n_225),
.B2(n_232),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_33),
.B1(n_36),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_25),
.B1(n_77),
.B2(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_123),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_123),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_6),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_33),
.B1(n_36),
.B2(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_7),
.A2(n_43),
.B1(n_60),
.B2(n_77),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_27),
.B1(n_77),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_10),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_33),
.B1(n_36),
.B2(n_135),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_135),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_135),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_11),
.A2(n_28),
.B1(n_56),
.B2(n_57),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_11),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_33),
.B1(n_36),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_13),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_125),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_125),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_13),
.A2(n_25),
.B1(n_42),
.B2(n_125),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_14),
.A2(n_33),
.B1(n_36),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_14),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_14),
.A2(n_27),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_72),
.Y(n_115)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_15),
.Y(n_153)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_15),
.Y(n_226)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_15),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_78),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_20),
.A2(n_21),
.B1(n_73),
.B2(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_44),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_46),
.C(n_61),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B1(n_32),
.B2(n_40),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_24),
.A2(n_31),
.B(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_26),
.B(n_35),
.C(n_36),
.Y(n_147)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_30),
.A2(n_40),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_30),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_30),
.A2(n_32),
.B1(n_134),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_30),
.A2(n_32),
.B1(n_142),
.B2(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_30),
.A2(n_270),
.B(n_292),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_30),
.A2(n_88),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_76),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_31),
.A2(n_128),
.B1(n_129),
.B2(n_133),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_31),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_33),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_33),
.A2(n_37),
.B(n_131),
.C(n_147),
.Y(n_146)
);

HAxp5_ASAP7_75t_SL g177 ( 
.A(n_33),
.B(n_132),
.CON(n_177),
.SN(n_177)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_36),
.A2(n_51),
.A3(n_66),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_39),
.B(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_73),
.C(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_45),
.A2(n_46),
.B1(n_79),
.B2(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_55),
.B(n_58),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_48),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_48),
.A2(n_59),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_48),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_48),
.A2(n_186),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_48),
.A2(n_185),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_48),
.A2(n_184),
.B1(n_185),
.B2(n_205),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_48),
.A2(n_185),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_48),
.A2(n_119),
.B(n_264),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_51),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_50),
.B(n_67),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_51),
.B(n_207),
.Y(n_206)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_55),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_55),
.B(n_58),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_55),
.B(n_132),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_56),
.B(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_121),
.B(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_65),
.B(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_64),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_65),
.A2(n_69),
.B1(n_168),
.B2(n_177),
.Y(n_182)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_68),
.A2(n_126),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_73),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_73),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_78),
.B(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_79),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_81),
.A2(n_121),
.B1(n_126),
.B2(n_296),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_83),
.A2(n_121),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_322),
.A3(n_332),
.B1(n_335),
.B2(n_336),
.C(n_339),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_301),
.B(n_321),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_278),
.B(n_300),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_169),
.B(n_254),
.C(n_277),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_154),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_154),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_138),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_116),
.B1(n_136),
.B2(n_137),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_101),
.B(n_137),
.C(n_138),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_102),
.B(n_107),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_103),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_104),
.B(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_114),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_108),
.A2(n_114),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_108),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_108),
.A2(n_222),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_108),
.A2(n_180),
.B(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_113),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_109),
.B(n_115),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_109),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_111),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_127),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_132),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_275)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_155),
.B(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_158),
.B(n_160),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_164),
.B1(n_165),
.B2(n_191),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_161),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_163),
.B(n_216),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_249),
.B(n_253),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_199),
.B(n_248),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_187),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_174),
.B(n_187),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.C(n_183),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_175),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_182),
.B(n_183),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_195),
.C(n_198),
.Y(n_250)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_197),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_243),
.B(n_247),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_218),
.B(n_242),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_228),
.B(n_241),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_227),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_227),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_235),
.B(n_240),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_275),
.B2(n_276),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_266),
.C(n_276),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_265),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_265),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_262),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_274),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_271),
.C(n_274),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_279),
.B(n_280),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_299),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_287),
.B1(n_297),
.B2(n_298),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_298),
.C(n_299),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_285),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_286),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_315),
.B(n_316),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_291),
.C(n_294),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_303),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_319),
.B2(n_320),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_311),
.B1(n_317),
.B2(n_318),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_318),
.C(n_320),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_309),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_309),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_324),
.C(n_329),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_310),
.B(n_324),
.CI(n_329),
.CON(n_334),
.SN(n_334)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_334),
.Y(n_338)
);


endmodule