module fake_jpeg_2211_n_490 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_490);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_490;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_56),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_84),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_64),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_66),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_90),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_15),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_29),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_91),
.Y(n_148)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_13),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_14),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_95),
.B(n_109),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_12),
.B(n_11),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_98),
.B(n_0),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_18),
.B(n_11),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_53),
.B(n_0),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_117),
.Y(n_156)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_49),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_54),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_47),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_62),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_26),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_122),
.B(n_124),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_57),
.B(n_54),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_123),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_63),
.B(n_26),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_57),
.A2(n_49),
.B1(n_48),
.B2(n_54),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_137),
.B1(n_92),
.B2(n_100),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_62),
.A2(n_119),
.B1(n_49),
.B2(n_48),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_37),
.B1(n_21),
.B2(n_42),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_143),
.A2(n_152),
.B1(n_159),
.B2(n_193),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_71),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_147),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_67),
.A2(n_37),
.B1(n_21),
.B2(n_31),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_158),
.B(n_139),
.C(n_136),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_69),
.A2(n_31),
.B1(n_40),
.B2(n_42),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_163),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_73),
.Y(n_163)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_169),
.Y(n_255)
);

INVx6_ASAP7_75t_SL g173 ( 
.A(n_91),
.Y(n_173)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

NAND2x1_ASAP7_75t_L g174 ( 
.A(n_104),
.B(n_54),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_174),
.B(n_136),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_93),
.B(n_27),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_96),
.B(n_27),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_107),
.B(n_25),
.C(n_41),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_78),
.A2(n_25),
.B1(n_41),
.B2(n_33),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_81),
.B(n_33),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_55),
.B(n_28),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_86),
.B(n_28),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_146),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_58),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_201),
.A2(n_144),
.B1(n_169),
.B2(n_191),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_176),
.B1(n_45),
.B2(n_148),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_202),
.A2(n_205),
.B1(n_249),
.B2(n_253),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_129),
.A2(n_99),
.B1(n_102),
.B2(n_97),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_204),
.A2(n_224),
.B1(n_239),
.B2(n_244),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_207),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_120),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_208),
.B(n_211),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_130),
.B(n_75),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

OAI211xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_103),
.B(n_47),
.C(n_75),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_126),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_236),
.Y(n_283)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_152),
.A2(n_45),
.B1(n_101),
.B2(n_47),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_103),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_228),
.A2(n_229),
.B(n_233),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_174),
.A2(n_30),
.B(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_128),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_232),
.A2(n_254),
.B1(n_257),
.B2(n_265),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_123),
.B(n_9),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_134),
.B(n_3),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_159),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_178),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_241),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_164),
.Y(n_241)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_128),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_246),
.Y(n_309)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_164),
.A2(n_4),
.B(n_6),
.C(n_8),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_248),
.A2(n_250),
.B(n_205),
.C(n_202),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_191),
.A2(n_8),
.B1(n_9),
.B2(n_145),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_137),
.A2(n_9),
.B1(n_153),
.B2(n_138),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_156),
.B(n_125),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_258),
.Y(n_300)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_140),
.Y(n_252)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_145),
.A2(n_144),
.B1(n_149),
.B2(n_166),
.Y(n_254)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_172),
.Y(n_256)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_142),
.A2(n_167),
.B1(n_172),
.B2(n_189),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_127),
.B(n_161),
.Y(n_258)
);

NAND2xp67_ASAP7_75t_SL g259 ( 
.A(n_189),
.B(n_197),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_194),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_263),
.Y(n_307)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_182),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_267),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_138),
.A2(n_153),
.B1(n_182),
.B2(n_171),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_132),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_269),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_141),
.A2(n_170),
.B(n_200),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_139),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_207),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_139),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_270),
.B(n_275),
.C(n_284),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_141),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_272),
.B(n_297),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_154),
.B1(n_175),
.B2(n_170),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_274),
.A2(n_278),
.B1(n_279),
.B2(n_288),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_203),
.B(n_155),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_213),
.A2(n_154),
.B1(n_175),
.B2(n_171),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_287),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_221),
.A2(n_200),
.B1(n_215),
.B2(n_229),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_231),
.A2(n_224),
.B1(n_204),
.B2(n_232),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_233),
.A2(n_244),
.B1(n_209),
.B2(n_239),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_286),
.A2(n_302),
.B(n_276),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_205),
.A2(n_250),
.B1(n_233),
.B2(n_249),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_233),
.B(n_206),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_227),
.A2(n_228),
.B1(n_259),
.B2(n_216),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_308),
.A2(n_271),
.B1(n_286),
.B2(n_307),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_243),
.B1(n_223),
.B2(n_219),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_313),
.B1(n_256),
.B2(n_255),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_206),
.A2(n_257),
.B1(n_254),
.B2(n_248),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_210),
.B(n_212),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_305),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_290),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_323),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_266),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_292),
.A2(n_234),
.B(n_242),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_321),
.A2(n_324),
.B(n_355),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_214),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_297),
.A2(n_242),
.B(n_250),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_346),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_331),
.Y(n_360)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_271),
.A2(n_264),
.B1(n_252),
.B2(n_262),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_328),
.A2(n_329),
.B1(n_303),
.B2(n_309),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_279),
.A2(n_289),
.B1(n_278),
.B2(n_288),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_332),
.B1(n_293),
.B2(n_301),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_255),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_237),
.B1(n_310),
.B2(n_272),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_270),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_340),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_325),
.Y(n_385)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_306),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_347),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_302),
.C(n_282),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_344),
.Y(n_369)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_284),
.B(n_291),
.C(n_285),
.Y(n_344)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

AO22x1_ASAP7_75t_SL g346 ( 
.A1(n_276),
.A2(n_274),
.B1(n_304),
.B2(n_295),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_281),
.B(n_282),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_276),
.A2(n_308),
.A3(n_296),
.B1(n_316),
.B2(n_291),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_353),
.Y(n_368)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

OA22x2_ASAP7_75t_SL g350 ( 
.A1(n_316),
.A2(n_281),
.B1(n_285),
.B2(n_318),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_350),
.Y(n_357)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_349),
.Y(n_384)
);

AOI21xp33_ASAP7_75t_L g355 ( 
.A1(n_312),
.A2(n_309),
.B(n_298),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g359 ( 
.A1(n_327),
.A2(n_293),
.B1(n_301),
.B2(n_317),
.Y(n_359)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_312),
.B(n_317),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_363),
.A2(n_364),
.B1(n_370),
.B2(n_374),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_330),
.A2(n_273),
.B1(n_305),
.B2(n_303),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_322),
.A2(n_332),
.B1(n_334),
.B2(n_338),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_322),
.A2(n_329),
.B1(n_343),
.B2(n_346),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_375),
.A2(n_382),
.B1(n_341),
.B2(n_344),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_379),
.A2(n_385),
.B1(n_354),
.B2(n_345),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g380 ( 
.A1(n_343),
.A2(n_353),
.A3(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_368),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_346),
.A2(n_324),
.B1(n_335),
.B2(n_351),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_321),
.A2(n_333),
.B(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_383),
.B(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_384),
.Y(n_388)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_390),
.A2(n_393),
.B1(n_400),
.B2(n_407),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_369),
.C(n_383),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_404),
.C(n_401),
.Y(n_414)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_375),
.A2(n_328),
.B1(n_350),
.B2(n_352),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_357),
.A2(n_339),
.B1(n_342),
.B2(n_336),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_397),
.Y(n_423)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_401),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_372),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_374),
.A2(n_364),
.B1(n_356),
.B2(n_382),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_369),
.B(n_368),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_365),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_402),
.B(n_406),
.Y(n_427)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_358),
.C(n_367),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_357),
.A2(n_358),
.B1(n_356),
.B2(n_367),
.Y(n_405)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_378),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_385),
.B1(n_363),
.B2(n_379),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_360),
.A2(n_380),
.B1(n_366),
.B2(n_373),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_409),
.B(n_359),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_376),
.B1(n_361),
.B2(n_372),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_376),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_410),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_413),
.B(n_387),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_418),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_359),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_416),
.B(n_421),
.C(n_425),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_359),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_361),
.C(n_359),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_394),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_424),
.B(n_386),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_404),
.Y(n_425)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_428),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_409),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_389),
.C(n_393),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_428),
.A2(n_400),
.B(n_407),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_432),
.A2(n_440),
.B(n_445),
.Y(n_452)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_411),
.Y(n_433)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_413),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_446),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_430),
.A2(n_423),
.B1(n_389),
.B2(n_419),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_438),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_442),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_430),
.A2(n_392),
.B(n_395),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_412),
.C(n_416),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_422),
.C(n_444),
.Y(n_453)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_427),
.B(n_396),
.Y(n_443)
);

OAI322xp33_ASAP7_75t_L g450 ( 
.A1(n_443),
.A2(n_426),
.A3(n_420),
.B1(n_422),
.B2(n_412),
.C1(n_411),
.C2(n_421),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_429),
.A2(n_403),
.B(n_418),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_423),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_431),
.A2(n_417),
.B(n_425),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_448),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_449),
.B(n_438),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_456),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_458),
.C(n_449),
.Y(n_467)
);

BUFx12_ASAP7_75t_L g456 ( 
.A(n_440),
.Y(n_456)
);

NOR2x1_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_446),
.Y(n_457)
);

AOI221xp5_ASAP7_75t_L g465 ( 
.A1(n_457),
.A2(n_432),
.B1(n_433),
.B2(n_436),
.C(n_454),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_444),
.C(n_441),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_458),
.B(n_435),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_434),
.C(n_445),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_460),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_437),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_467),
.C(n_447),
.Y(n_475)
);

XNOR2x1_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_457),
.Y(n_474)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_465),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_454),
.B(n_452),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_452),
.Y(n_469)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_457),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_474),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_459),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_479),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_462),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_462),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_474),
.Y(n_483)
);

NOR3xp33_ASAP7_75t_SL g481 ( 
.A(n_478),
.B(n_470),
.C(n_471),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_477),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_477),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_484),
.A2(n_485),
.B(n_482),
.Y(n_486)
);

A2O1A1O1Ixp25_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_447),
.B(n_455),
.C(n_456),
.D(n_463),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_455),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_488),
.B(n_456),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_SL g490 ( 
.A(n_489),
.B(n_456),
.Y(n_490)
);


endmodule