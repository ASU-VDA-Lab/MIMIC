module fake_netlist_1_12118_n_969 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_969);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_969;
wire n_117;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_185;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_627;
wire n_532;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_786;
wire n_228;
wire n_724;
wire n_599;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_961;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_822;
wire n_706;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_948;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_962;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_967;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_695;
wire n_650;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g112 ( .A(n_2), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_44), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_2), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_84), .B(n_57), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_37), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_19), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_89), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_87), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_47), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_24), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_8), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_73), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_103), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_109), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_20), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_5), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_51), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_10), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_52), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_111), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_7), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_21), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_72), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_85), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_77), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
BUFx10_ASAP7_75t_L g142 ( .A(n_42), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_13), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_22), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_43), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_106), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_29), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_45), .Y(n_151) );
CKINVDCx14_ASAP7_75t_R g152 ( .A(n_105), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_133), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_156) );
OAI22xp33_ASAP7_75t_SL g157 ( .A1(n_119), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_113), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_113), .B(n_4), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_141), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_114), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_129), .B(n_5), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_120), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_115), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_128), .B(n_6), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_124), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_126), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx8_ASAP7_75t_L g180 ( .A(n_161), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_165), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_159), .B(n_121), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_165), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_169), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_169), .Y(n_190) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_168), .A2(n_117), .B(n_147), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
AO22x2_ASAP7_75t_L g196 ( .A1(n_161), .A2(n_148), .B1(n_149), .B2(n_146), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_171), .B(n_142), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_163), .B(n_145), .C(n_151), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_163), .Y(n_203) );
NAND2xp33_ASAP7_75t_R g204 ( .A(n_153), .B(n_116), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_160), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_173), .B(n_142), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_164), .B(n_142), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g212 ( .A(n_164), .B(n_132), .C(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
NOR2x1p5_ASAP7_75t_L g214 ( .A(n_178), .B(n_116), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_178), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_176), .B(n_118), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_170), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_170), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
AO22x2_ASAP7_75t_L g223 ( .A1(n_175), .A2(n_112), .B1(n_134), .B2(n_143), .Y(n_223) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_179), .A2(n_152), .B(n_139), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_172), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_175), .B(n_118), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_172), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_172), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_167), .B(n_130), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_172), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_167), .B(n_125), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_156), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_177), .B(n_125), .Y(n_234) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_174), .A2(n_139), .B(n_135), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_177), .Y(n_237) );
AND2x6_ASAP7_75t_L g238 ( .A(n_177), .B(n_123), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_203), .B(n_132), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_203), .B(n_135), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_229), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_232), .B(n_167), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_193), .B(n_157), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_193), .B(n_166), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_193), .B(n_166), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_193), .B(n_162), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_199), .B(n_162), .Y(n_247) );
INVxp67_ASAP7_75t_SL g248 ( .A(n_184), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_180), .A2(n_177), .B(n_131), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_190), .B(n_130), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_209), .B(n_131), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_196), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_180), .B(n_150), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_211), .B(n_23), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_196), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_217), .B(n_25), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_180), .B(n_26), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_180), .B(n_27), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_180), .B(n_6), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_221), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_199), .B(n_7), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_221), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_191), .B(n_8), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_191), .B(n_9), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_200), .B(n_28), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_191), .B(n_9), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_235), .B(n_10), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_235), .B(n_11), .Y(n_269) );
NAND2xp33_ASAP7_75t_L g270 ( .A(n_196), .B(n_30), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_200), .B(n_31), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_204), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_272) );
O2A1O1Ixp5_ASAP7_75t_L g273 ( .A1(n_224), .A2(n_67), .B(n_108), .C(n_107), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_226), .B(n_64), .Y(n_275) );
NOR2x1p5_ASAP7_75t_L g276 ( .A(n_187), .B(n_14), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_235), .B(n_14), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_212), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_184), .B(n_15), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_212), .B(n_66), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_234), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_224), .B(n_15), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_183), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_208), .B(n_68), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_225), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_223), .B(n_16), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_215), .B(n_16), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_188), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_208), .B(n_69), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_214), .B(n_17), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_223), .B(n_17), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g294 ( .A(n_181), .B(n_18), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_181), .B(n_70), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_223), .B(n_238), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_223), .B(n_18), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_181), .B(n_71), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_238), .B(n_19), .Y(n_299) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_238), .B(n_20), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_214), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_241), .B(n_238), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_246), .A2(n_218), .B(n_237), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_252), .A2(n_233), .B1(n_238), .B2(n_236), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_286), .A2(n_181), .B(n_207), .C(n_185), .Y(n_305) );
CKINVDCx14_ASAP7_75t_R g306 ( .A(n_279), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_248), .B(n_238), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_274), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_283), .B(n_238), .Y(n_309) );
AOI33xp33_ASAP7_75t_L g310 ( .A1(n_301), .A2(n_237), .A3(n_236), .B1(n_216), .B2(n_218), .B3(n_219), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_255), .B(n_185), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_256), .B(n_185), .Y(n_312) );
INVxp33_ASAP7_75t_SL g313 ( .A(n_253), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_244), .A2(n_216), .B(n_219), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_239), .B(n_185), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_245), .A2(n_222), .B(n_220), .Y(n_316) );
CKINVDCx8_ASAP7_75t_R g317 ( .A(n_257), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_274), .Y(n_318) );
OR2x6_ASAP7_75t_L g319 ( .A(n_247), .B(n_207), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_270), .B(n_222), .C(n_220), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_240), .A2(n_231), .B(n_230), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_278), .A2(n_273), .B(n_264), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
OAI321xp33_ASAP7_75t_L g324 ( .A1(n_293), .A2(n_195), .A3(n_213), .B1(n_182), .B2(n_202), .C(n_194), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_247), .B(n_207), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_265), .A2(n_207), .B(n_230), .C(n_231), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_242), .A2(n_231), .B(n_230), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_297), .A2(n_228), .B(n_227), .C(n_213), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_267), .A2(n_195), .B(n_228), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_243), .B(n_227), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_251), .B(n_32), .Y(n_332) );
OR2x6_ASAP7_75t_L g333 ( .A(n_291), .B(n_182), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_249), .A2(n_210), .B(n_206), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_250), .B(n_34), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_300), .B(n_201), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_276), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_262), .B(n_182), .C(n_194), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_268), .A2(n_210), .B(n_206), .C(n_186), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_281), .A2(n_186), .B(n_192), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_296), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_269), .A2(n_197), .B1(n_192), .B2(n_198), .Y(n_344) );
AOI21x1_ASAP7_75t_L g345 ( .A1(n_280), .A2(n_197), .B(n_198), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_287), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_261), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_337), .A2(n_272), .B1(n_277), .B2(n_282), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_313), .B(n_260), .Y(n_352) );
AOI21x1_ASAP7_75t_SL g353 ( .A1(n_302), .A2(n_299), .B(n_280), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_319), .Y(n_355) );
OR2x6_ASAP7_75t_L g356 ( .A(n_337), .B(n_258), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_307), .B(n_257), .Y(n_357) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_322), .A2(n_275), .B(n_254), .C(n_284), .Y(n_358) );
CKINVDCx11_ASAP7_75t_R g359 ( .A(n_317), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_343), .B(n_254), .Y(n_360) );
OAI22x1_ASAP7_75t_L g361 ( .A1(n_338), .A2(n_271), .B1(n_266), .B2(n_289), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_322), .A2(n_259), .B(n_271), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_275), .B(n_284), .C(n_266), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_335), .A2(n_295), .B(n_294), .C(n_289), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_309), .B(n_295), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_333), .B(n_292), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_326), .A2(n_292), .B(n_285), .Y(n_369) );
INVx3_ASAP7_75t_SL g370 ( .A(n_337), .Y(n_370) );
OAI21x1_ASAP7_75t_SL g371 ( .A1(n_304), .A2(n_285), .B(n_263), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_318), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_306), .A2(n_263), .B1(n_298), .B2(n_202), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_346), .B(n_205), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_327), .A2(n_288), .B(n_205), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_333), .B(n_288), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_333), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_336), .B(n_205), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_345), .A2(n_202), .B(n_194), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_362), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_376), .B(n_342), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_365), .A2(n_340), .B(n_330), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_359), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_367), .A2(n_315), .B1(n_339), .B2(n_318), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_354), .B(n_308), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_376), .Y(n_387) );
CKINVDCx6p67_ASAP7_75t_R g388 ( .A(n_370), .Y(n_388) );
OAI21x1_ASAP7_75t_SL g389 ( .A1(n_371), .A2(n_330), .B(n_305), .Y(n_389) );
NOR2x1_ASAP7_75t_SL g390 ( .A(n_377), .B(n_348), .Y(n_390) );
XOR2xp5_ASAP7_75t_L g391 ( .A(n_352), .B(n_325), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_363), .A2(n_320), .B(n_324), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_350), .Y(n_393) );
AO31x2_ASAP7_75t_L g394 ( .A1(n_358), .A2(n_321), .A3(n_334), .B(n_342), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_353), .A2(n_329), .B(n_344), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_353), .A2(n_341), .B(n_314), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_347), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_379), .A2(n_316), .B(n_303), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_378), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g400 ( .A(n_354), .B(n_348), .Y(n_400) );
BUFx4f_ASAP7_75t_SL g401 ( .A(n_355), .Y(n_401) );
NAND2x1_ASAP7_75t_L g402 ( .A(n_356), .B(n_348), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_351), .B(n_328), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_369), .A2(n_312), .B(n_311), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_351), .B(n_201), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_372), .B(n_201), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_324), .B(n_201), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_357), .Y(n_410) );
OAI21x1_ASAP7_75t_L g411 ( .A1(n_366), .A2(n_201), .B(n_189), .Y(n_411) );
INVx6_ASAP7_75t_L g412 ( .A(n_356), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_411), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_411), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_394), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_394), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_388), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_410), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_410), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_404), .B(n_358), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_388), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_397), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_387), .Y(n_431) );
OAI222xp33_ASAP7_75t_L g432 ( .A1(n_403), .A2(n_356), .B1(n_360), .B2(n_373), .C1(n_361), .C2(n_359), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_404), .B(n_365), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_409), .Y(n_437) );
OAI21x1_ASAP7_75t_L g438 ( .A1(n_409), .A2(n_364), .B(n_189), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
OR2x2_ASAP7_75t_SL g440 ( .A(n_412), .B(n_383), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_407), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_396), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_387), .B(n_364), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_387), .B(n_35), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_412), .B(n_189), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_391), .Y(n_447) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_389), .A2(n_189), .B(n_188), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_401), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_387), .B(n_189), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_382), .B(n_188), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_395), .A2(n_188), .B(n_38), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_395), .A2(n_188), .B(n_39), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_398), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_386), .B(n_36), .Y(n_459) );
NAND2xp33_ASAP7_75t_R g460 ( .A(n_384), .B(n_40), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_398), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_385), .A2(n_41), .B(n_46), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_386), .B(n_48), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_400), .Y(n_464) );
OR2x6_ASAP7_75t_L g465 ( .A(n_412), .B(n_49), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_389), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_392), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_384), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_412), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_424), .B(n_386), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_413), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_440), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_439), .B(n_381), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_390), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_467), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_422), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_465), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_425), .B(n_390), .Y(n_483) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_438), .A2(n_405), .B(n_408), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_422), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_415), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_430), .Y(n_488) );
AOI221x1_ASAP7_75t_SL g489 ( .A1(n_439), .A2(n_50), .B1(n_53), .B2(n_54), .C(n_55), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_436), .B(n_392), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_434), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_428), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_433), .B(n_405), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_431), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_425), .B(n_392), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_465), .A2(n_392), .B1(n_58), .B2(n_60), .Y(n_498) );
AO31x2_ASAP7_75t_L g499 ( .A1(n_418), .A2(n_56), .A3(n_61), .B(n_62), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_427), .B(n_63), .Y(n_500) );
AND2x4_ASAP7_75t_SL g501 ( .A(n_429), .B(n_74), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_428), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_418), .B(n_75), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_447), .B(n_110), .Y(n_505) );
INVx4_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_455), .B(n_76), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_466), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_418), .Y(n_512) );
AND2x4_ASAP7_75t_SL g513 ( .A(n_429), .B(n_82), .Y(n_513) );
INVx4_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_426), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_459), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_459), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_440), .B(n_83), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_463), .Y(n_520) );
OAI321xp33_ASAP7_75t_L g521 ( .A1(n_462), .A2(n_86), .A3(n_88), .B1(n_91), .B2(n_92), .C(n_93), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_467), .Y(n_522) );
AND2x4_ASAP7_75t_SL g523 ( .A(n_465), .B(n_94), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_419), .B(n_95), .Y(n_524) );
INVx5_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_467), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_463), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_442), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_469), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_469), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_453), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_431), .B(n_104), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_453), .B(n_96), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_419), .B(n_97), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_420), .B(n_98), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_458), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_442), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_442), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_420), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_420), .B(n_100), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_423), .B(n_101), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_423), .B(n_102), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_423), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_435), .B(n_441), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_435), .B(n_441), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_435), .B(n_458), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_431), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_433), .B(n_450), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_446), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_464), .B(n_431), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_444), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_444), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_464), .B(n_450), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_431), .B(n_450), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_444), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_433), .B(n_450), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_431), .B(n_433), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_431), .B(n_448), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_448), .B(n_457), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_457), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_457), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_461), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_446), .Y(n_563) );
AND3x1_ASAP7_75t_L g564 ( .A(n_449), .B(n_460), .C(n_468), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_461), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_448), .B(n_461), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_446), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_525), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_492), .B(n_448), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_506), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_491), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_492), .B(n_414), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_481), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_472), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_558), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_472), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_480), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_479), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_470), .B(n_446), .Y(n_579) );
OR2x6_ASAP7_75t_L g580 ( .A(n_506), .B(n_445), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_488), .B(n_449), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_480), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_479), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_558), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_485), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_522), .Y(n_586) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_481), .B(n_432), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_548), .B(n_414), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_470), .B(n_445), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_493), .B(n_414), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_477), .B(n_445), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_485), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_477), .B(n_445), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_487), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_487), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_526), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_562), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_493), .B(n_416), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_505), .B(n_432), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_471), .B(n_452), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_471), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_473), .Y(n_604) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_473), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_474), .B(n_452), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_474), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_478), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_507), .B(n_486), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_478), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_546), .B(n_416), .Y(n_612) );
AND2x4_ASAP7_75t_SL g613 ( .A(n_506), .B(n_416), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_531), .B(n_451), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_546), .B(n_438), .Y(n_615) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_486), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_503), .B(n_438), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_476), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_503), .B(n_437), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_547), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_508), .B(n_437), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_494), .B(n_462), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_536), .B(n_451), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_483), .B(n_454), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_494), .B(n_451), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_559), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_483), .B(n_456), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_502), .B(n_454), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_502), .B(n_437), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_565), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_550), .B(n_517), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_550), .B(n_454), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_508), .B(n_454), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_518), .B(n_456), .Y(n_635) );
BUFx2_ASAP7_75t_L g636 ( .A(n_496), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_520), .B(n_456), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_529), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_530), .B(n_456), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_548), .B(n_514), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_527), .B(n_544), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_511), .B(n_515), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_512), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_525), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_509), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_512), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_544), .B(n_545), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_516), .Y(n_649) );
NAND2x1_ASAP7_75t_L g650 ( .A(n_514), .B(n_482), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_496), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_509), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_514), .B(n_519), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_553), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_545), .B(n_490), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_482), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_490), .B(n_500), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_516), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_553), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_548), .B(n_557), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_539), .B(n_543), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_500), .B(n_539), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_525), .B(n_482), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_549), .B(n_567), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_543), .B(n_566), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_489), .B(n_567), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_549), .B(n_563), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_554), .B(n_557), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_554), .B(n_475), .Y(n_669) );
INVxp33_ASAP7_75t_L g670 ( .A(n_519), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_560), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_560), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_475), .B(n_525), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_525), .B(n_524), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_504), .B(n_534), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_497), .B(n_534), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_504), .B(n_535), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_542), .B(n_556), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_556), .B(n_495), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_521), .B(n_498), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_566), .B(n_495), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_523), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_561), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_561), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_528), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_528), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_524), .B(n_535), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_495), .B(n_537), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_542), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_537), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_538), .B(n_551), .Y(n_691) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_523), .Y(n_692) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_540), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_571), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_574), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_576), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_616), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_618), .B(n_538), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_577), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_654), .B(n_555), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_603), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_582), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_585), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_603), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_594), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_659), .B(n_555), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_668), .B(n_541), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_648), .B(n_541), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_596), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_597), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_575), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_605), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_638), .Y(n_713) );
NAND2x1p5_ASAP7_75t_L g714 ( .A(n_682), .B(n_564), .Y(n_714) );
INVx3_ASAP7_75t_L g715 ( .A(n_645), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_646), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_648), .B(n_540), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_652), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_665), .B(n_552), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_575), .Y(n_720) );
INVxp67_ASAP7_75t_L g721 ( .A(n_584), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_605), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_665), .B(n_552), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_642), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_643), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_661), .B(n_551), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_578), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_604), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_608), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_609), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_578), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_583), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_661), .B(n_484), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_611), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_584), .B(n_484), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_683), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_669), .B(n_501), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_627), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_587), .B(n_510), .C(n_532), .D(n_533), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_627), .B(n_640), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_640), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_581), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_636), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_655), .B(n_484), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_572), .B(n_484), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_681), .B(n_501), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_681), .B(n_513), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_621), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_641), .B(n_513), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_579), .B(n_499), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_651), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_664), .B(n_499), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_657), .B(n_499), .Y(n_753) );
OR2x2_ASAP7_75t_L g754 ( .A(n_662), .B(n_499), .Y(n_754) );
BUFx2_ASAP7_75t_L g755 ( .A(n_573), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_572), .B(n_499), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_682), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_680), .A2(n_666), .B(n_670), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_591), .B(n_600), .Y(n_759) );
INVx1_ASAP7_75t_SL g760 ( .A(n_673), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_632), .B(n_593), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_591), .B(n_600), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_685), .Y(n_763) );
OR2x2_ASAP7_75t_L g764 ( .A(n_678), .B(n_667), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_660), .B(n_676), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_660), .B(n_644), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_644), .Y(n_767) );
INVxp67_ASAP7_75t_L g768 ( .A(n_685), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_647), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_569), .B(n_620), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_569), .B(n_620), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_647), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_660), .B(n_649), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_649), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_583), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_595), .B(n_589), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_622), .B(n_658), .Y(n_777) );
OR2x2_ASAP7_75t_L g778 ( .A(n_658), .B(n_606), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_622), .B(n_617), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_679), .B(n_675), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_586), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_617), .B(n_684), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_679), .B(n_677), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_641), .B(n_679), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_674), .B(n_641), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_610), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_671), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_586), .Y(n_788) );
BUFx2_ASAP7_75t_L g789 ( .A(n_692), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_688), .B(n_612), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_688), .B(n_612), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_670), .B(n_693), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_602), .B(n_592), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_590), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_653), .B(n_610), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_656), .B(n_570), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_671), .B(n_684), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_590), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_656), .B(n_570), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_592), .B(n_598), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_672), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_672), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_598), .B(n_689), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_630), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_656), .B(n_570), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_738), .B(n_615), .Y(n_806) );
INVx2_ASAP7_75t_SL g807 ( .A(n_697), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_740), .B(n_687), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_694), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_713), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_789), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_780), .B(n_613), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_740), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_741), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_759), .B(n_615), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_786), .B(n_601), .Y(n_816) );
INVx2_ASAP7_75t_SL g817 ( .A(n_757), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_758), .A2(n_601), .B1(n_580), .B2(n_663), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_695), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_696), .Y(n_820) );
INVx1_ASAP7_75t_SL g821 ( .A(n_760), .Y(n_821) );
INVxp67_ASAP7_75t_L g822 ( .A(n_748), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_783), .B(n_613), .Y(n_823) );
AOI211xp5_ASAP7_75t_L g824 ( .A1(n_758), .A2(n_663), .B(n_568), .C(n_645), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_724), .B(n_623), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_699), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_742), .B(n_568), .Y(n_827) );
A2O1A1Ixp33_ASAP7_75t_L g828 ( .A1(n_795), .A2(n_650), .B(n_645), .C(n_635), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_804), .B(n_635), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_722), .B(n_629), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_702), .Y(n_831) );
INVx1_ASAP7_75t_SL g832 ( .A(n_760), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_703), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_714), .A2(n_580), .B1(n_645), .B2(n_624), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_705), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_744), .B(n_629), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_725), .B(n_637), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_790), .B(n_580), .Y(n_838) );
OR2x2_ASAP7_75t_L g839 ( .A(n_759), .B(n_619), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_709), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_784), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_744), .B(n_599), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_710), .Y(n_843) );
CKINVDCx16_ASAP7_75t_R g844 ( .A(n_749), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_763), .Y(n_845) );
INVxp67_ASAP7_75t_L g846 ( .A(n_755), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_762), .B(n_619), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_762), .B(n_631), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_791), .B(n_588), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_716), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_769), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_714), .B(n_626), .Y(n_852) );
NOR2x1p5_ASAP7_75t_L g853 ( .A(n_749), .B(n_614), .Y(n_853) );
OR2x2_ASAP7_75t_L g854 ( .A(n_770), .B(n_599), .Y(n_854) );
OR2x2_ASAP7_75t_L g855 ( .A(n_770), .B(n_607), .Y(n_855) );
OR2x2_ASAP7_75t_L g856 ( .A(n_771), .B(n_607), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_718), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_768), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_736), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_761), .B(n_588), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_728), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_785), .B(n_588), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_729), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_782), .B(n_690), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_784), .B(n_625), .Y(n_865) );
INVx1_ASAP7_75t_SL g866 ( .A(n_711), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_768), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_782), .B(n_631), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_743), .B(n_628), .Y(n_869) );
AND2x4_ASAP7_75t_L g870 ( .A(n_796), .B(n_633), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_720), .B(n_691), .Y(n_871) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_721), .A2(n_639), .B(n_634), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_776), .B(n_691), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_750), .A2(n_691), .B1(n_686), .B2(n_690), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_751), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_813), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_844), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_814), .Y(n_878) );
OAI31xp33_ASAP7_75t_L g879 ( .A1(n_811), .A2(n_737), .A3(n_721), .B(n_746), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_836), .B(n_779), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_818), .A2(n_792), .B1(n_747), .B2(n_765), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g882 ( .A1(n_824), .A2(n_739), .B1(n_752), .B2(n_735), .C(n_753), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_841), .B(n_764), .Y(n_883) );
AOI31xp33_ASAP7_75t_L g884 ( .A1(n_824), .A2(n_773), .A3(n_766), .B(n_799), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_809), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_858), .Y(n_886) );
INVx3_ASAP7_75t_L g887 ( .A(n_811), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_810), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_819), .Y(n_889) );
INVxp33_ASAP7_75t_L g890 ( .A(n_852), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_866), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_820), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_816), .B(n_739), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_853), .A2(n_771), .B1(n_779), .B2(n_723), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_815), .B(n_723), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_826), .Y(n_896) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_866), .Y(n_897) );
AOI21xp33_ASAP7_75t_L g898 ( .A1(n_834), .A2(n_698), .B(n_754), .Y(n_898) );
OAI21xp33_ASAP7_75t_L g899 ( .A1(n_836), .A2(n_777), .B(n_719), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_831), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_833), .Y(n_901) );
OAI332xp33_ASAP7_75t_L g902 ( .A1(n_825), .A2(n_756), .A3(n_733), .B1(n_719), .B2(n_777), .B3(n_778), .C1(n_745), .C2(n_698), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_822), .A2(n_707), .B1(n_717), .B2(n_708), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g904 ( .A(n_828), .B(n_706), .C(n_700), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_846), .A2(n_733), .B1(n_726), .B2(n_730), .C(n_734), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_835), .Y(n_906) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_830), .B(n_700), .C(n_706), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_840), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g909 ( .A1(n_821), .A2(n_715), .B1(n_756), .B2(n_745), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_830), .B(n_701), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_862), .B(n_805), .Y(n_911) );
AOI21xp33_ASAP7_75t_SL g912 ( .A1(n_817), .A2(n_715), .B(n_793), .Y(n_912) );
AOI21xp33_ASAP7_75t_L g913 ( .A1(n_875), .A2(n_803), .B(n_704), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_910), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g915 ( .A(n_893), .B(n_874), .C(n_827), .D(n_869), .Y(n_915) );
OAI21xp33_ASAP7_75t_L g916 ( .A1(n_893), .A2(n_829), .B(n_821), .Y(n_916) );
AOI21xp33_ASAP7_75t_L g917 ( .A1(n_890), .A2(n_807), .B(n_867), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_897), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_902), .B(n_845), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_897), .Y(n_920) );
NOR2xp33_ASAP7_75t_SL g921 ( .A(n_877), .B(n_832), .Y(n_921) );
O2A1O1Ixp33_ASAP7_75t_L g922 ( .A1(n_884), .A2(n_832), .B(n_850), .C(n_843), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_877), .A2(n_812), .B(n_823), .C(n_838), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_876), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_890), .A2(n_870), .B1(n_808), .B2(n_865), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_894), .A2(n_857), .B1(n_859), .B2(n_861), .C(n_863), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g927 ( .A1(n_879), .A2(n_871), .B1(n_864), .B2(n_868), .C(n_842), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_905), .B(n_851), .Y(n_928) );
AOI321xp33_ASAP7_75t_L g929 ( .A1(n_882), .A2(n_872), .A3(n_806), .B1(n_837), .B2(n_870), .C(n_842), .Y(n_929) );
OAI321xp33_ASAP7_75t_L g930 ( .A1(n_909), .A2(n_868), .A3(n_864), .B1(n_847), .B2(n_839), .C(n_848), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_912), .A2(n_860), .B1(n_873), .B2(n_856), .Y(n_931) );
AOI21xp33_ASAP7_75t_L g932 ( .A1(n_909), .A2(n_712), .B(n_855), .Y(n_932) );
AOI21xp33_ASAP7_75t_SL g933 ( .A1(n_887), .A2(n_854), .B(n_849), .Y(n_933) );
INVx1_ASAP7_75t_SL g934 ( .A(n_887), .Y(n_934) );
AOI211xp5_ASAP7_75t_L g935 ( .A1(n_922), .A2(n_898), .B(n_904), .C(n_913), .Y(n_935) );
NAND4xp25_ASAP7_75t_L g936 ( .A(n_929), .B(n_881), .C(n_878), .D(n_903), .Y(n_936) );
OAI211xp5_ASAP7_75t_L g937 ( .A1(n_922), .A2(n_899), .B(n_891), .C(n_903), .Y(n_937) );
AOI221x1_ASAP7_75t_L g938 ( .A1(n_916), .A2(n_892), .B1(n_908), .B2(n_888), .C(n_906), .Y(n_938) );
NOR2xp67_ASAP7_75t_L g939 ( .A(n_930), .B(n_907), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_914), .Y(n_940) );
AOI311xp33_ASAP7_75t_L g941 ( .A1(n_927), .A2(n_889), .A3(n_885), .B(n_901), .C(n_900), .Y(n_941) );
NAND4xp75_ASAP7_75t_L g942 ( .A(n_919), .B(n_883), .C(n_880), .D(n_896), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_933), .A2(n_895), .B(n_911), .C(n_886), .Y(n_943) );
AOI211x1_ASAP7_75t_SL g944 ( .A1(n_917), .A2(n_886), .B(n_726), .C(n_797), .Y(n_944) );
AOI21xp33_ASAP7_75t_SL g945 ( .A1(n_931), .A2(n_797), .B(n_802), .Y(n_945) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_936), .B(n_921), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_943), .B(n_934), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_940), .Y(n_948) );
NOR2x1_ASAP7_75t_L g949 ( .A(n_942), .B(n_915), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g950 ( .A(n_937), .B(n_928), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_944), .B(n_926), .Y(n_951) );
OAI322xp33_ASAP7_75t_L g952 ( .A1(n_950), .A2(n_945), .A3(n_918), .B1(n_920), .B2(n_941), .C1(n_939), .C2(n_924), .Y(n_952) );
NOR2x1_ASAP7_75t_L g953 ( .A(n_949), .B(n_937), .Y(n_953) );
NAND3x1_ASAP7_75t_SL g954 ( .A(n_947), .B(n_935), .C(n_938), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_946), .B(n_925), .Y(n_955) );
NOR2xp67_ASAP7_75t_L g956 ( .A(n_955), .B(n_948), .Y(n_956) );
AND3x2_ASAP7_75t_L g957 ( .A(n_954), .B(n_951), .C(n_923), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_953), .B(n_932), .Y(n_958) );
XOR2xp5_ASAP7_75t_L g959 ( .A(n_958), .B(n_952), .Y(n_959) );
AOI22xp5_ASAP7_75t_SL g960 ( .A1(n_957), .A2(n_801), .B1(n_787), .B2(n_774), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_959), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_960), .A2(n_956), .B1(n_772), .B2(n_767), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_961), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_962), .B(n_781), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_963), .B(n_775), .Y(n_965) );
AOI222xp33_ASAP7_75t_L g966 ( .A1(n_965), .A2(n_964), .B1(n_727), .B2(n_731), .C1(n_732), .C2(n_788), .Y(n_966) );
AO21x2_ASAP7_75t_L g967 ( .A1(n_966), .A2(n_964), .B(n_794), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_967), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_968), .A2(n_798), .B1(n_800), .B2(n_686), .Y(n_969) );
endmodule