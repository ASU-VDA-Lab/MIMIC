module fake_ibex_359_n_2416 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2416);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2416;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_422;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_399;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_398;
wire n_2377;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_864;
wire n_608;
wire n_412;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2390;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_458;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_2358;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2252;
wire n_1982;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_444;
wire n_1761;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_2395;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2251;
wire n_722;
wire n_2012;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_415;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_424;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_924;
wire n_2331;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_401;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_866;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_408;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_1506;
wire n_559;
wire n_425;

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_53),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_327),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_119),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_54),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_109),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_42),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_293),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_346),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_18),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_202),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_26),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_349),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_48),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_6),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_47),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_57),
.Y(n_415)
);

BUFx8_ASAP7_75t_SL g416 ( 
.A(n_333),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_104),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_46),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_104),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_102),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_350),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_374),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_155),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_308),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_302),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_251),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_336),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_382),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_252),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_260),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_228),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_50),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_295),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_179),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_213),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_241),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_16),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_190),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_378),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_397),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_297),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_40),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_116),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_36),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_230),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_127),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_38),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_110),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_117),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_115),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_99),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_247),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_335),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_188),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_329),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_395),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_223),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_181),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_23),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_307),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_168),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_161),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_29),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_249),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_330),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_86),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_52),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_87),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_31),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_238),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_37),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_290),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_70),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_100),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_334),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_216),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_314),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_245),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_292),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_119),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_154),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_9),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_123),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_248),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_78),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_64),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_149),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_98),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_13),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_207),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_384),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_146),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_366),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_233),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_1),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_362),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_133),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_95),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_265),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_385),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_321),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_19),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_376),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_347),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_143),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_367),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_261),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_9),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_115),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_206),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_380),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_0),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_54),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_135),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_51),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_211),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_278),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_64),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_205),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_317),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_324),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_118),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_51),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_162),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_27),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_23),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_152),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_217),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_105),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_58),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_1),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_162),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_319),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_74),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_129),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_66),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_130),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_157),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_95),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_38),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_4),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_147),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_246),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_117),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_5),
.Y(n_548)
);

BUFx8_ASAP7_75t_SL g549 ( 
.A(n_268),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_361),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_19),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_345),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_56),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_171),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_235),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_218),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_214),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_369),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_164),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_355),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_141),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_168),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_166),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_185),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_33),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_316),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_194),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_221),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_305),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_348),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_176),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_291),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_210),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_364),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_341),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_301),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_109),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_61),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_147),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_118),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_129),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_250),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_78),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_368),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_337),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_232),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_83),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_152),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_320),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_53),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_0),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_275),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_7),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_42),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_56),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_288),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_88),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_338),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_318),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_283),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_381),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_31),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_81),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_197),
.Y(n_604)
);

CKINVDCx14_ASAP7_75t_R g605 ( 
.A(n_79),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_74),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_27),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_138),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_289),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_121),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_138),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_93),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_201),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_309),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_363),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_328),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_88),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_105),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_294),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_92),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_331),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_272),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_8),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_170),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_231),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_255),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_68),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_68),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_343),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_57),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_344),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_63),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_171),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_225),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_183),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_310),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_339),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_323),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_140),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_102),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_83),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_300),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_178),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_99),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_130),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_322),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_365),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_121),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_340),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_126),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_342),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_372),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_12),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_40),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_282),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_156),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_35),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_287),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_46),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_50),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_332),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_69),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_125),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_325),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_195),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_196),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_326),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_354),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_17),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_63),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_18),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_143),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_311),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_286),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_198),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_352),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_182),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_150),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_112),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_91),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_75),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_356),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_22),
.Y(n_683)
);

INVxp33_ASAP7_75t_SL g684 ( 
.A(n_398),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_402),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_605),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_441),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_542),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_554),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_445),
.B(n_636),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_554),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_416),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_549),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_415),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_597),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_445),
.B(n_2),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_597),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_558),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_421),
.B(n_177),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_432),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_417),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_432),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_R g704 ( 
.A(n_474),
.B(n_499),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_508),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_508),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_581),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_581),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_400),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_400),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_410),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_410),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_459),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_459),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_412),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_437),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_468),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_443),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_468),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_462),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_610),
.B(n_501),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_501),
.B(n_2),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_660),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_660),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_670),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_406),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_670),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_401),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_403),
.Y(n_729)
);

CKINVDCx16_ASAP7_75t_R g730 ( 
.A(n_470),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_636),
.B(n_3),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_503),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_507),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_504),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_412),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_407),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_463),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_513),
.Y(n_738)
);

INVxp67_ASAP7_75t_SL g739 ( 
.A(n_414),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_522),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_419),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_446),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_448),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_473),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_488),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_570),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_487),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_470),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_413),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_507),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_500),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_604),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_614),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_511),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_521),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_413),
.B(n_3),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_526),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_616),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_510),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_408),
.B(n_4),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_409),
.B(n_5),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_539),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_R g763 ( 
.A(n_435),
.B(n_180),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_530),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_541),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_675),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_544),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_425),
.B(n_6),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_538),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_545),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_563),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_565),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_571),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_577),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_579),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_418),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_587),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_438),
.B(n_439),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_580),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_588),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_418),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_590),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_420),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_632),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_606),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_611),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_612),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_618),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_399),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_623),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_399),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_630),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_633),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_639),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_653),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_510),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_404),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_404),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_640),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_644),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_648),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_663),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_466),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_405),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_525),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_525),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_466),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_672),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_683),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_466),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_481),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_481),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_420),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_525),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_726),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_690),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_715),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_696),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_691),
.B(n_423),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_733),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_803),
.B(n_423),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_733),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_698),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_750),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_689),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_732),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_807),
.B(n_657),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_810),
.B(n_657),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_734),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_692),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_701),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_750),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_703),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_759),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_811),
.B(n_659),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_738),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_740),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_812),
.B(n_659),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_705),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_731),
.B(n_651),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_809),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_746),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_R g843 ( 
.A(n_711),
.B(n_662),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_759),
.Y(n_844)
);

AND2x6_ASAP7_75t_L g845 ( 
.A(n_697),
.B(n_460),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_706),
.B(n_651),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_707),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_708),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_723),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_699),
.B(n_739),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_686),
.B(n_470),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_749),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_796),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_728),
.B(n_514),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_796),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_729),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_747),
.B(n_662),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_736),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_741),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_684),
.B(n_789),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_684),
.B(n_669),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_709),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_711),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_710),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_752),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_753),
.Y(n_866)
);

INVx6_ASAP7_75t_L g867 ( 
.A(n_730),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_713),
.Y(n_868)
);

OA21x2_ASAP7_75t_L g869 ( 
.A1(n_806),
.A2(n_436),
.B(n_434),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_809),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_742),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_758),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_714),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_748),
.B(n_528),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_717),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_743),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_766),
.Y(n_877)
);

CKINVDCx11_ASAP7_75t_R g878 ( 
.A(n_695),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_695),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_712),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_719),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_791),
.B(n_669),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_702),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_744),
.A2(n_456),
.B(n_453),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_751),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_712),
.B(n_528),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_755),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_797),
.B(n_405),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_762),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_693),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_724),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_798),
.B(n_804),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_694),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_765),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_704),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_767),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_778),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_725),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_727),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_R g900 ( 
.A(n_687),
.B(n_411),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_735),
.B(n_528),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_687),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_814),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_735),
.B(n_680),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_770),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_776),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_771),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_773),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_774),
.B(n_458),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_702),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_779),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_780),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_776),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_785),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_786),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_781),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_790),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_781),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_792),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_783),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_783),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_794),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_716),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_685),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_813),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_813),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_685),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_799),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_801),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_754),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_782),
.B(n_680),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_716),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_787),
.B(n_671),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_760),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_793),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_718),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_800),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_761),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_756),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_700),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_688),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_768),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_721),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_688),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_722),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_805),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_718),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_720),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_763),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_720),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_737),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_737),
.B(n_671),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_745),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_745),
.B(n_678),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_757),
.Y(n_956)
);

CKINVDCx6p67_ASAP7_75t_R g957 ( 
.A(n_757),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_R g958 ( 
.A(n_764),
.B(n_678),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_764),
.A2(n_681),
.B1(n_683),
.B2(n_679),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_769),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_769),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_772),
.B(n_679),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_772),
.B(n_681),
.Y(n_963)
);

OA21x2_ASAP7_75t_L g964 ( 
.A1(n_775),
.A2(n_480),
.B(n_471),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_775),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_777),
.Y(n_966)
);

AND2x6_ASAP7_75t_L g967 ( 
.A(n_777),
.B(n_460),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_784),
.B(n_411),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_784),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_795),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_795),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_802),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_802),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_808),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_808),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_690),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_733),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_803),
.B(n_496),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_726),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_690),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_686),
.B(n_680),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_726),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_690),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_733),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_690),
.B(n_422),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_726),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_690),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_809),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_726),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_733),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_733),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_696),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_733),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_726),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_726),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_690),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_690),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_711),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_690),
.B(n_422),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_726),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_726),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_690),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_690),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_803),
.B(n_525),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_686),
.B(n_481),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_731),
.B(n_524),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_SL g1007 ( 
.A(n_730),
.B(n_424),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_690),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_693),
.B(n_424),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_733),
.Y(n_1010)
);

OA21x2_ASAP7_75t_L g1011 ( 
.A1(n_731),
.A2(n_552),
.B(n_550),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_690),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_789),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_715),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_715),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_690),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_803),
.B(n_525),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_733),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_733),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_690),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_726),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_726),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_992),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_947),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_1004),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_1004),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_940),
.B(n_426),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_947),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_884),
.B(n_935),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_911),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_1017),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_820),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_992),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_880),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_820),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_867),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_852),
.B(n_442),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_820),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_985),
.B(n_426),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_867),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1017),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_935),
.B(n_555),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_819),
.B(n_497),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_867),
.B(n_594),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_818),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_863),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_1007),
.B(n_427),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_823),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_998),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_1014),
.Y(n_1050)
);

AO22x2_ASAP7_75t_L g1051 ( 
.A1(n_857),
.A2(n_551),
.B1(n_595),
.B2(n_484),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_861),
.B(n_628),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_1014),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_820),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_903),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_953),
.B(n_444),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_1013),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_824),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_824),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_881),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_932),
.B(n_447),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_878),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1015),
.B(n_874),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_823),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_999),
.B(n_427),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_849),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_1015),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_839),
.Y(n_1068)
);

INVx6_ASAP7_75t_L g1069 ( 
.A(n_864),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_1013),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_931),
.B(n_497),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_816),
.A2(n_450),
.B1(n_451),
.B2(n_449),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_957),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_976),
.B(n_461),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_857),
.B(n_467),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_824),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_839),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_935),
.B(n_939),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_881),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_875),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_875),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_851),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_962),
.B(n_963),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_825),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_943),
.B(n_428),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_864),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_824),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_843),
.B(n_428),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_943),
.B(n_429),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_856),
.B(n_429),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_832),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_980),
.B(n_469),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_830),
.Y(n_1093)
);

AO22x2_ASAP7_75t_L g1094 ( 
.A1(n_934),
.A2(n_557),
.B1(n_560),
.B2(n_556),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_895),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_832),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_936),
.A2(n_608),
.B1(n_594),
.B2(n_572),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_862),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_862),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_903),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_935),
.B(n_939),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_858),
.B(n_430),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_897),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_934),
.B(n_817),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_832),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_859),
.B(n_430),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_868),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_983),
.B(n_987),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_832),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_868),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_996),
.B(n_475),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_869),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_997),
.B(n_476),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_913),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_864),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_991),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1002),
.B(n_482),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_873),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_991),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_873),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_898),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_938),
.B(n_497),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_821),
.B(n_629),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_898),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_831),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_991),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_991),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_993),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_L g1129 ( 
.A(n_845),
.B(n_682),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_833),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_913),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_847),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_993),
.Y(n_1133)
);

NAND2xp33_ASAP7_75t_L g1134 ( 
.A(n_845),
.B(n_682),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_848),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_919),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1003),
.B(n_483),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_853),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_967),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_L g1140 ( 
.A(n_845),
.B(n_939),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_911),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_958),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_864),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1008),
.A2(n_489),
.B1(n_490),
.B2(n_485),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_L g1145 ( 
.A(n_843),
.B(n_494),
.C(n_491),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_939),
.B(n_574),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_920),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_869),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_827),
.B(n_629),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_891),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_920),
.B(n_585),
.Y(n_1151)
);

AND2x6_ASAP7_75t_L g1152 ( 
.A(n_886),
.B(n_495),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_923),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_919),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_993),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_871),
.B(n_431),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_967),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1012),
.B(n_498),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_967),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_L g1160 ( 
.A(n_845),
.B(n_433),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_923),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_929),
.B(n_599),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_828),
.B(n_629),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1016),
.B(n_505),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_929),
.B(n_600),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1020),
.B(n_512),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_891),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_993),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_876),
.B(n_433),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_841),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_850),
.B(n_901),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_981),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_891),
.Y(n_1173)
);

AND2x2_ASAP7_75t_SL g1174 ( 
.A(n_964),
.B(n_594),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_966),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_869),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_891),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1010),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_835),
.B(n_631),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_885),
.B(n_658),
.Y(n_1180)
);

AND2x2_ASAP7_75t_SL g1181 ( 
.A(n_964),
.B(n_888),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1011),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1010),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_899),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_899),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_887),
.B(n_601),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_899),
.Y(n_1187)
);

AND2x6_ASAP7_75t_L g1188 ( 
.A(n_904),
.B(n_850),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_889),
.B(n_658),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_967),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_899),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_916),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_822),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_822),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1010),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1005),
.B(n_515),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_834),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_900),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1011),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_978),
.B(n_894),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1010),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1011),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_834),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_900),
.B(n_516),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_844),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_896),
.B(n_609),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_844),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_955),
.A2(n_625),
.B1(n_635),
.B2(n_615),
.Y(n_1208)
);

INVx4_ASAP7_75t_SL g1209 ( 
.A(n_845),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_855),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_860),
.B(n_517),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_906),
.B(n_917),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_855),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_905),
.B(n_661),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_977),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_964),
.B(n_907),
.Y(n_1216)
);

AND2x2_ASAP7_75t_SL g1217 ( 
.A(n_892),
.B(n_594),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_977),
.Y(n_1218)
);

INVx8_ASAP7_75t_L g1219 ( 
.A(n_967),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_984),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_921),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_984),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_990),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_870),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_908),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_922),
.Y(n_1226)
);

AND2x2_ASAP7_75t_SL g1227 ( 
.A(n_955),
.B(n_594),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_912),
.B(n_661),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_914),
.B(n_664),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_990),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_915),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_918),
.B(n_664),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_838),
.B(n_518),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1018),
.Y(n_1234)
);

AND2x6_ASAP7_75t_L g1235 ( 
.A(n_978),
.B(n_495),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_956),
.B(n_961),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1006),
.B(n_631),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_930),
.B(n_665),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1018),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1019),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_926),
.B(n_527),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_854),
.B(n_1006),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_840),
.B(n_631),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_946),
.B(n_529),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1019),
.Y(n_1245)
);

AND2x6_ASAP7_75t_L g1246 ( 
.A(n_909),
.B(n_586),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_846),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_846),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_840),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_909),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_927),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_854),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_944),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_950),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1009),
.B(n_532),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_944),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_958),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_882),
.A2(n_534),
.B1(n_535),
.B2(n_533),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_950),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1009),
.B(n_537),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_941),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_968),
.B(n_665),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_902),
.B(n_540),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_959),
.B(n_543),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_956),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_956),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1225),
.B(n_1231),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1225),
.B(n_1231),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1233),
.B(n_547),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1252),
.B(n_548),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1055),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1053),
.B(n_925),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1233),
.B(n_553),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1034),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1050),
.B(n_559),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1050),
.B(n_561),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1055),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1136),
.B(n_815),
.Y(n_1278)
);

AND2x6_ASAP7_75t_SL g1279 ( 
.A(n_1170),
.B(n_951),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1044),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1067),
.B(n_666),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1047),
.B(n_666),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1114),
.B(n_1022),
.Y(n_1283)
);

NAND2x1_ASAP7_75t_L g1284 ( 
.A(n_1044),
.B(n_1069),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1083),
.B(n_969),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1181),
.A2(n_608),
.B1(n_622),
.B2(n_586),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1057),
.B(n_960),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1199),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1170),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1057),
.B(n_673),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1062),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1250),
.B(n_562),
.Y(n_1292)
);

AND2x6_ASAP7_75t_SL g1293 ( 
.A(n_1062),
.B(n_970),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1181),
.A2(n_608),
.B1(n_622),
.B2(n_637),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1030),
.A2(n_829),
.B1(n_836),
.B2(n_826),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1070),
.B(n_673),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1066),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1100),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1045),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1070),
.B(n_960),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1030),
.B(n_578),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1051),
.A2(n_988),
.B1(n_956),
.B2(n_973),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1203),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1049),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1046),
.Y(n_1305)
);

O2A1O1Ixp5_ASAP7_75t_L g1306 ( 
.A1(n_1029),
.A2(n_667),
.B(n_647),
.C(n_566),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1027),
.B(n_1085),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1089),
.B(n_583),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1084),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1221),
.B(n_837),
.Y(n_1310)
);

BUFx8_ASAP7_75t_L g1311 ( 
.A(n_1226),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1203),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1174),
.A2(n_1182),
.B1(n_1199),
.B2(n_1200),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1088),
.B(n_674),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1088),
.B(n_674),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1044),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1171),
.B(n_971),
.Y(n_1317)
);

AND2x6_ASAP7_75t_SL g1318 ( 
.A(n_1212),
.B(n_879),
.Y(n_1318)
);

BUFx4_ASAP7_75t_L g1319 ( 
.A(n_1073),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1154),
.B(n_1021),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1131),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1175),
.B(n_972),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1242),
.A2(n_591),
.B(n_602),
.C(n_593),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1108),
.B(n_603),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1139),
.B(n_608),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1131),
.B(n_842),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1029),
.A2(n_621),
.B(n_531),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1171),
.B(n_1082),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1211),
.B(n_1093),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1174),
.A2(n_608),
.B1(n_617),
.B2(n_607),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1063),
.B(n_865),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1259),
.B(n_676),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1236),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1259),
.B(n_676),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1125),
.B(n_620),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1130),
.B(n_624),
.Y(n_1336)
);

NOR3xp33_ASAP7_75t_SL g1337 ( 
.A(n_1142),
.B(n_942),
.C(n_928),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1132),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1135),
.B(n_1200),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1192),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_L g1342 ( 
.A(n_1182),
.B(n_677),
.Y(n_1342)
);

OR2x6_ASAP7_75t_L g1343 ( 
.A(n_1219),
.B(n_961),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1200),
.B(n_627),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1200),
.B(n_641),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1221),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1056),
.B(n_645),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1104),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1123),
.B(n_650),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1219),
.B(n_961),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1060),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1259),
.B(n_677),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1036),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1052),
.B(n_972),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1037),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1078),
.A2(n_649),
.B(n_642),
.Y(n_1356)
);

OR2x6_ASAP7_75t_L g1357 ( 
.A(n_1219),
.B(n_961),
.Y(n_1357)
);

NOR3xp33_ASAP7_75t_L g1358 ( 
.A(n_1145),
.B(n_1001),
.C(n_872),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1227),
.A2(n_1061),
.B1(n_1188),
.B2(n_1208),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1123),
.B(n_654),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1200),
.B(n_656),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1112),
.Y(n_1362)
);

AND2x6_ASAP7_75t_L g1363 ( 
.A(n_1112),
.B(n_566),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1203),
.Y(n_1364)
);

NOR2xp67_ASAP7_75t_L g1365 ( 
.A(n_1251),
.B(n_1103),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1240),
.Y(n_1366)
);

INVx5_ASAP7_75t_L g1367 ( 
.A(n_1202),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1188),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1148),
.A2(n_975),
.B1(n_973),
.B2(n_626),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1148),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1227),
.A2(n_877),
.B1(n_979),
.B2(n_866),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1240),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1217),
.A2(n_982),
.B1(n_989),
.B2(n_986),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1251),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1149),
.B(n_994),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1039),
.B(n_995),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1196),
.B(n_945),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1224),
.A2(n_910),
.B1(n_924),
.B2(n_883),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1065),
.B(n_1000),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1090),
.B(n_440),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1102),
.B(n_452),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1078),
.A2(n_455),
.B(n_454),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1176),
.A2(n_1216),
.B1(n_1217),
.B2(n_1246),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1061),
.B(n_973),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1176),
.A2(n_975),
.B1(n_973),
.B2(n_626),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1106),
.B(n_457),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_1103),
.B(n_890),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1259),
.B(n_464),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1156),
.B(n_465),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1216),
.A2(n_933),
.B(n_948),
.C(n_937),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1257),
.B(n_893),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1198),
.B(n_472),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1060),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1025),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1236),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1101),
.A2(n_1140),
.B(n_1134),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1169),
.B(n_477),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1025),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1180),
.B(n_478),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1079),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1079),
.B(n_479),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1189),
.B(n_486),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1188),
.A2(n_975),
.B1(n_952),
.B2(n_954),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1149),
.B(n_975),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1261),
.B(n_492),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1261),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1026),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1188),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1214),
.B(n_493),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1246),
.A2(n_626),
.B1(n_668),
.B2(n_566),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1026),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1074),
.B(n_949),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1246),
.A2(n_626),
.B1(n_668),
.B2(n_566),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1261),
.B(n_502),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1196),
.B(n_1172),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1261),
.B(n_506),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1163),
.B(n_509),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_SL g1418 ( 
.A(n_1097),
.B(n_520),
.C(n_519),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1246),
.A2(n_626),
.B1(n_668),
.B2(n_566),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1204),
.B(n_523),
.Y(n_1421)
);

O2A1O1Ixp5_ASAP7_75t_L g1422 ( 
.A1(n_1101),
.A2(n_1146),
.B(n_1042),
.C(n_1151),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1163),
.B(n_536),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1139),
.B(n_546),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1179),
.B(n_564),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1031),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1232),
.B(n_567),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1031),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1157),
.B(n_568),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1179),
.B(n_569),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1188),
.A2(n_974),
.B1(n_965),
.B2(n_575),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1236),
.B(n_668),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_L g1433 ( 
.A(n_1202),
.B(n_573),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1040),
.B(n_668),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1262),
.B(n_576),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1210),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1138),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1074),
.B(n_7),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1043),
.B(n_582),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1092),
.B(n_8),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1202),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1210),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1095),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1041),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1092),
.B(n_1111),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1215),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1238),
.B(n_584),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1202),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1208),
.A2(n_592),
.B1(n_596),
.B2(n_589),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_SL g1450 ( 
.A1(n_1043),
.A2(n_1237),
.B(n_1243),
.C(n_1122),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1080),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1157),
.B(n_598),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1159),
.B(n_655),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1265),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1215),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1140),
.A2(n_619),
.B(n_613),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1095),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1024),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1113),
.B(n_634),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1257),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1072),
.A2(n_13),
.B(n_10),
.C(n_11),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1266),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1263),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1237),
.B(n_638),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1111),
.B(n_14),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1137),
.B(n_643),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1081),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1158),
.B(n_646),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1263),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1243),
.B(n_652),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1223),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1239),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1117),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1159),
.B(n_15),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1023),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1246),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1117),
.B(n_20),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_R g1478 ( 
.A(n_1129),
.B(n_1134),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1166),
.B(n_21),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1235),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1033),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1164),
.B(n_24),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1051),
.Y(n_1483)
);

NOR3xp33_ASAP7_75t_L g1484 ( 
.A(n_1264),
.B(n_25),
.C(n_26),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1141),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1071),
.B(n_28),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1186),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1147),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1239),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1152),
.B(n_1071),
.Y(n_1490)
);

BUFx12f_ASAP7_75t_L g1491 ( 
.A(n_1164),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1256),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1051),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1153),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1129),
.B(n_30),
.C(n_32),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_R g1496 ( 
.A(n_1160),
.B(n_32),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1152),
.B(n_33),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1249),
.A2(n_186),
.B(n_184),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1190),
.B(n_34),
.Y(n_1499)
);

NOR2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1255),
.B(n_1260),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1152),
.B(n_35),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1152),
.B(n_36),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1190),
.B(n_37),
.Y(n_1503)
);

O2A1O1Ixp5_ASAP7_75t_L g1504 ( 
.A1(n_1042),
.A2(n_43),
.B(n_39),
.C(n_41),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1241),
.B(n_39),
.Y(n_1505)
);

NOR2x2_ASAP7_75t_L g1506 ( 
.A(n_1094),
.B(n_41),
.Y(n_1506)
);

AND2x6_ASAP7_75t_SL g1507 ( 
.A(n_1244),
.B(n_43),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1161),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1122),
.B(n_44),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1048),
.Y(n_1510)
);

NAND2xp33_ASAP7_75t_L g1511 ( 
.A(n_1235),
.B(n_187),
.Y(n_1511)
);

INVx4_ASAP7_75t_L g1512 ( 
.A(n_1024),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1194),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1256),
.B(n_44),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1064),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1028),
.B(n_45),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1144),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1254),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1396),
.A2(n_1035),
.B(n_1032),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1274),
.B(n_1075),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1311),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1297),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1311),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_SL g1524 ( 
.A(n_1302),
.B(n_1097),
.C(n_1146),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1304),
.B(n_1258),
.Y(n_1525)
);

AO22x1_ASAP7_75t_L g1526 ( 
.A1(n_1289),
.A2(n_1235),
.B1(n_1244),
.B2(n_1094),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1321),
.B(n_1209),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1267),
.B(n_1094),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1299),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1309),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1338),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1278),
.B(n_1028),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1272),
.B(n_1253),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1268),
.B(n_1098),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1305),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1437),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1307),
.A2(n_1254),
.B(n_1107),
.C(n_1110),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1329),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1340),
.Y(n_1539)
);

CKINVDCx8_ASAP7_75t_R g1540 ( 
.A(n_1279),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1436),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1359),
.A2(n_1118),
.B1(n_1120),
.B2(n_1099),
.Y(n_1542)
);

NOR3xp33_ASAP7_75t_SL g1543 ( 
.A(n_1373),
.B(n_1206),
.C(n_1186),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1291),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1492),
.Y(n_1545)
);

AND2x6_ASAP7_75t_SL g1546 ( 
.A(n_1319),
.B(n_1247),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1346),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1442),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1285),
.A2(n_1160),
.B1(n_1235),
.B2(n_1077),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_SL g1550 ( 
.A(n_1302),
.B(n_1496),
.C(n_1484),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1444),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1446),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1420),
.B(n_1121),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1346),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1313),
.A2(n_1514),
.B1(n_1383),
.B2(n_1370),
.Y(n_1555)
);

BUFx4f_ASAP7_75t_L g1556 ( 
.A(n_1463),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1348),
.B(n_1124),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1288),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1432),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1326),
.B(n_1348),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1280),
.B(n_1116),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1280),
.B(n_1209),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1445),
.B(n_1354),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1455),
.Y(n_1564)
);

NAND2x2_ASAP7_75t_L g1565 ( 
.A(n_1457),
.B(n_1500),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1374),
.B(n_1365),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1514),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1510),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1515),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1484),
.A2(n_1206),
.B1(n_1162),
.B2(n_1165),
.C(n_1151),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1443),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1331),
.B(n_1194),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1374),
.B(n_1209),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1362),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1451),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1310),
.B(n_1295),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1491),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1458),
.Y(n_1578)
);

NOR3xp33_ASAP7_75t_SL g1579 ( 
.A(n_1378),
.B(n_1165),
.C(n_1162),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1467),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1362),
.B(n_1248),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1283),
.B(n_1320),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1471),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1370),
.B(n_1248),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1432),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1472),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1368),
.B(n_1068),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1293),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1485),
.B(n_1245),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1488),
.B(n_1494),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1318),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1353),
.B(n_1245),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1483),
.A2(n_1222),
.B1(n_1220),
.B2(n_1197),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1475),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1355),
.B(n_1220),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1287),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1347),
.B(n_1328),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_R g1598 ( 
.A(n_1322),
.B(n_1235),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1349),
.B(n_1127),
.C(n_1116),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1368),
.B(n_1222),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_R g1601 ( 
.A(n_1517),
.B(n_1193),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1337),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1489),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1271),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1432),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1508),
.B(n_1205),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1481),
.B(n_1207),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1458),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1512),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1333),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1408),
.B(n_1116),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1347),
.B(n_1213),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1301),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1395),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1408),
.B(n_1116),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1412),
.B(n_1218),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1479),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1288),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1493),
.A2(n_1234),
.B1(n_1230),
.B2(n_1069),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1512),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1438),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1328),
.B(n_1127),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1371),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1387),
.B(n_1391),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1288),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1486),
.B(n_1167),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_L g1627 ( 
.A(n_1377),
.B(n_1493),
.C(n_1461),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1317),
.A2(n_1069),
.B1(n_1115),
.B2(n_1086),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1384),
.B(n_1127),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_R g1630 ( 
.A(n_1507),
.B(n_1086),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1288),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1269),
.B(n_1127),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1269),
.B(n_1115),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1277),
.Y(n_1634)
);

AND3x1_ASAP7_75t_L g1635 ( 
.A(n_1337),
.B(n_1150),
.C(n_1143),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1440),
.Y(n_1636)
);

AND3x1_ASAP7_75t_SL g1637 ( 
.A(n_1506),
.B(n_45),
.C(n_47),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1486),
.B(n_1450),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_L g1639 ( 
.A(n_1363),
.B(n_1038),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1465),
.B(n_1143),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1287),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1473),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1316),
.B(n_1038),
.Y(n_1643)
);

OR2x2_ASAP7_75t_SL g1644 ( 
.A(n_1376),
.B(n_48),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1300),
.B(n_1469),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1335),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1336),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1300),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_R g1649 ( 
.A(n_1418),
.B(n_1150),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1394),
.Y(n_1650)
);

INVx5_ASAP7_75t_L g1651 ( 
.A(n_1363),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1434),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1339),
.B(n_1173),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1398),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1367),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1407),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1411),
.Y(n_1657)
);

NAND2xp33_ASAP7_75t_SL g1658 ( 
.A(n_1478),
.B(n_1038),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1367),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_SL g1660 ( 
.A(n_1390),
.B(n_1184),
.C(n_1177),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1298),
.B(n_1185),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1298),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1434),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1441),
.A2(n_1422),
.B(n_1306),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1367),
.B(n_1187),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1505),
.B(n_1191),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1426),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1428),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1518),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1363),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1462),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1292),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1516),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1448),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1367),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1324),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1379),
.B(n_1032),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1415),
.A2(n_1054),
.B1(n_1058),
.B2(n_1035),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1434),
.B(n_1038),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1270),
.Y(n_1680)
);

OR2x4_ASAP7_75t_L g1681 ( 
.A(n_1375),
.B(n_1059),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1351),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1406),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1275),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1375),
.B(n_1054),
.Y(n_1685)
);

NOR3xp33_ASAP7_75t_SL g1686 ( 
.A(n_1404),
.B(n_49),
.C(n_52),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1448),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1276),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1404),
.B(n_1058),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1349),
.B(n_49),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1509),
.B(n_1076),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_SL g1692 ( 
.A(n_1477),
.B(n_55),
.C(n_58),
.Y(n_1692)
);

BUFx4f_ASAP7_75t_L g1693 ( 
.A(n_1343),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1343),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1360),
.B(n_1076),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1449),
.B(n_1059),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_SL g1697 ( 
.A(n_1482),
.B(n_55),
.C(n_59),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1363),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1273),
.B(n_59),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1363),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1360),
.B(n_60),
.Y(n_1701)
);

OR2x6_ASAP7_75t_L g1702 ( 
.A(n_1343),
.B(n_1059),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1513),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1350),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1351),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1350),
.B(n_1059),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1313),
.A2(n_1383),
.B1(n_1294),
.B2(n_1286),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1441),
.B(n_1087),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1487),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1448),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1490),
.B(n_1087),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1350),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1448),
.Y(n_1713)
);

INVx5_ASAP7_75t_L g1714 ( 
.A(n_1357),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1308),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1284),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1421),
.B(n_1091),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1513),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1460),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1400),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1459),
.B(n_60),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1323),
.B(n_1096),
.Y(n_1722)
);

NAND2x2_ASAP7_75t_L g1723 ( 
.A(n_1466),
.B(n_1468),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1431),
.B(n_61),
.Y(n_1724)
);

NAND2x1p5_ASAP7_75t_L g1725 ( 
.A(n_1393),
.B(n_1133),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1357),
.Y(n_1726)
);

INVxp33_ASAP7_75t_L g1727 ( 
.A(n_1358),
.Y(n_1727)
);

NOR3xp33_ASAP7_75t_SL g1728 ( 
.A(n_1314),
.B(n_1315),
.C(n_1439),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1435),
.B(n_1105),
.Y(n_1729)
);

NOR3xp33_ASAP7_75t_SL g1730 ( 
.A(n_1439),
.B(n_62),
.C(n_65),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1435),
.B(n_1109),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1325),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1357),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1405),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1403),
.B(n_1133),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_R g1736 ( 
.A(n_1418),
.B(n_62),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1281),
.B(n_1109),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1400),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1325),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1504),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1504),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1344),
.B(n_1133),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1303),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1342),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1497),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1312),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1358),
.B(n_1119),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1341),
.Y(n_1748)
);

AO22x1_ASAP7_75t_L g1749 ( 
.A1(n_1417),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1417),
.B(n_67),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1364),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1454),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1464),
.B(n_1119),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1401),
.B(n_1126),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1501),
.Y(n_1755)
);

AND2x4_ASAP7_75t_SL g1756 ( 
.A(n_1476),
.B(n_1133),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1290),
.B(n_1126),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1414),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1416),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1366),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1502),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1372),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1296),
.B(n_1128),
.Y(n_1763)
);

AND2x4_ASAP7_75t_SL g1764 ( 
.A(n_1476),
.B(n_1155),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_SL g1765 ( 
.A(n_1480),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1388),
.B(n_1168),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1470),
.B(n_1178),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1306),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1474),
.B(n_1178),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1345),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1332),
.B(n_1183),
.Y(n_1771)
);

OR2x2_ASAP7_75t_SL g1772 ( 
.A(n_1495),
.B(n_69),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1535),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1538),
.B(n_1423),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1535),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1550),
.A2(n_1480),
.B(n_1330),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1563),
.B(n_1380),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1560),
.B(n_1423),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1519),
.A2(n_1498),
.B(n_1286),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1659),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_L g1781 ( 
.A1(n_1664),
.A2(n_1327),
.B(n_1499),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1655),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1531),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1740),
.A2(n_1330),
.B(n_1410),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1664),
.A2(n_1503),
.B(n_1413),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1601),
.B(n_1369),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1638),
.A2(n_1511),
.B(n_1433),
.Y(n_1787)
);

OAI22x1_ASAP7_75t_L g1788 ( 
.A1(n_1591),
.A2(n_1425),
.B1(n_1430),
.B2(n_1282),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1638),
.A2(n_1385),
.B(n_1369),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1550),
.A2(n_1430),
.B(n_1425),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1713),
.A2(n_1413),
.B(n_1410),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1534),
.A2(n_1356),
.B(n_1361),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1534),
.A2(n_1352),
.B(n_1334),
.Y(n_1793)
);

AO21x1_ASAP7_75t_L g1794 ( 
.A1(n_1707),
.A2(n_1429),
.B(n_1424),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1585),
.B(n_1385),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1616),
.B(n_1597),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1526),
.B(n_1392),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1625),
.A2(n_1419),
.B(n_1201),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1544),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1553),
.A2(n_1453),
.B(n_1452),
.Y(n_1800)
);

AOI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1741),
.A2(n_1456),
.B(n_1382),
.Y(n_1801)
);

AO31x2_ASAP7_75t_L g1802 ( 
.A1(n_1707),
.A2(n_1201),
.A3(n_1195),
.B(n_1470),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1642),
.B(n_1381),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1582),
.B(n_1386),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1566),
.B(n_1672),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1553),
.B(n_1389),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1676),
.B(n_1447),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1725),
.A2(n_1399),
.B(n_1397),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1680),
.B(n_1402),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1522),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1558),
.Y(n_1811)
);

OA22x2_ASAP7_75t_L g1812 ( 
.A1(n_1576),
.A2(n_1427),
.B1(n_1409),
.B2(n_72),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1722),
.A2(n_191),
.B(n_189),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1558),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1556),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1537),
.A2(n_70),
.B(n_71),
.Y(n_1816)
);

NAND2x1p5_ASAP7_75t_L g1817 ( 
.A(n_1693),
.B(n_71),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1525),
.B(n_72),
.Y(n_1818)
);

AO22x2_ASAP7_75t_L g1819 ( 
.A1(n_1542),
.A2(n_77),
.B1(n_73),
.B2(n_76),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1556),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1571),
.B(n_73),
.Y(n_1821)
);

NOR4xp25_ASAP7_75t_L g1822 ( 
.A(n_1528),
.B(n_79),
.C(n_76),
.D(n_77),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1529),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1521),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1709),
.A2(n_80),
.B(n_81),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1613),
.A2(n_80),
.B(n_82),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1585),
.B(n_82),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1722),
.A2(n_193),
.B(n_192),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1530),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1577),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1646),
.B(n_84),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1691),
.A2(n_200),
.B(n_199),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1768),
.A2(n_204),
.B(n_203),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1523),
.Y(n_1834)
);

O2A1O1Ixp5_ASAP7_75t_L g1835 ( 
.A1(n_1658),
.A2(n_1696),
.B(n_1735),
.C(n_1727),
.Y(n_1835)
);

AO31x2_ASAP7_75t_L g1836 ( 
.A1(n_1555),
.A2(n_1542),
.A3(n_1719),
.B(n_1528),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1742),
.A2(n_209),
.B(n_208),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1695),
.A2(n_84),
.B(n_85),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1631),
.A2(n_215),
.B(n_212),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1520),
.B(n_85),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1647),
.B(n_86),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1631),
.A2(n_222),
.B(n_220),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1715),
.B(n_87),
.Y(n_1843)
);

A2O1A1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1570),
.A2(n_89),
.B(n_90),
.C(n_91),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1708),
.A2(n_226),
.B(n_224),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1708),
.A2(n_229),
.B(n_227),
.Y(n_1846)
);

A2O1A1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1570),
.A2(n_1677),
.B(n_1673),
.C(n_1684),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1681),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1765),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1765),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1572),
.B(n_1688),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1711),
.A2(n_236),
.B(n_234),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1536),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1681),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1539),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1700),
.A2(n_239),
.B(n_237),
.Y(n_1856)
);

AO22x2_ASAP7_75t_L g1857 ( 
.A1(n_1555),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1557),
.B(n_97),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1557),
.B(n_98),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1568),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1627),
.B(n_100),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1590),
.A2(n_101),
.B1(n_103),
.B2(n_106),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1675),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1711),
.A2(n_242),
.B(n_240),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1695),
.A2(n_101),
.B(n_103),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1561),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1729),
.A2(n_244),
.B(n_243),
.Y(n_1867)
);

NAND2xp33_ASAP7_75t_L g1868 ( 
.A(n_1598),
.B(n_106),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1729),
.A2(n_254),
.B(n_253),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1590),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1693),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1569),
.Y(n_1872)
);

OAI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1762),
.A2(n_257),
.B(n_256),
.Y(n_1873)
);

AO21x1_ASAP7_75t_L g1874 ( 
.A1(n_1574),
.A2(n_107),
.B(n_108),
.Y(n_1874)
);

HAxp5_ASAP7_75t_L g1875 ( 
.A(n_1637),
.B(n_111),
.CON(n_1875),
.SN(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1753),
.A2(n_111),
.B(n_112),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1627),
.B(n_113),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1575),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1762),
.A2(n_259),
.B(n_258),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1580),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1731),
.A2(n_1767),
.B(n_1753),
.Y(n_1881)
);

NAND2xp33_ASAP7_75t_L g1882 ( 
.A(n_1732),
.B(n_113),
.Y(n_1882)
);

NOR4xp25_ASAP7_75t_L g1883 ( 
.A(n_1524),
.B(n_114),
.C(n_116),
.D(n_120),
.Y(n_1883)
);

NAND3xp33_ASAP7_75t_SL g1884 ( 
.A(n_1623),
.B(n_114),
.C(n_120),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1767),
.A2(n_122),
.B(n_123),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1612),
.B(n_1551),
.Y(n_1886)
);

BUFx2_ASAP7_75t_L g1887 ( 
.A(n_1641),
.Y(n_1887)
);

NAND2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1714),
.B(n_122),
.Y(n_1888)
);

AOI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1745),
.A2(n_280),
.B(n_394),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1685),
.A2(n_124),
.B(n_125),
.C(n_126),
.Y(n_1890)
);

OAI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1643),
.A2(n_1562),
.B(n_1581),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1731),
.A2(n_124),
.B(n_127),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1610),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1606),
.A2(n_1644),
.B1(n_1574),
.B2(n_1744),
.Y(n_1894)
);

AO21x1_ASAP7_75t_L g1895 ( 
.A1(n_1593),
.A2(n_128),
.B(n_131),
.Y(n_1895)
);

OAI21x1_ASAP7_75t_L g1896 ( 
.A1(n_1581),
.A2(n_284),
.B(n_393),
.Y(n_1896)
);

OAI21x1_ASAP7_75t_L g1897 ( 
.A1(n_1584),
.A2(n_281),
.B(n_391),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1617),
.B(n_128),
.Y(n_1898)
);

O2A1O1Ixp5_ASAP7_75t_L g1899 ( 
.A1(n_1744),
.A2(n_285),
.B(n_390),
.C(n_389),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1686),
.A2(n_277),
.B(n_388),
.Y(n_1900)
);

AO31x2_ASAP7_75t_L g1901 ( 
.A1(n_1567),
.A2(n_131),
.A3(n_132),
.B(n_133),
.Y(n_1901)
);

O2A1O1Ixp5_ASAP7_75t_L g1902 ( 
.A1(n_1700),
.A2(n_279),
.B(n_386),
.C(n_383),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1533),
.B(n_132),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1594),
.B(n_134),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1621),
.B(n_134),
.Y(n_1905)
);

AOI211x1_ASAP7_75t_L g1906 ( 
.A1(n_1749),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1714),
.B(n_136),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1743),
.A2(n_1751),
.B(n_1748),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1686),
.A2(n_296),
.B(n_379),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1566),
.B(n_137),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1541),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1579),
.B(n_139),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1626),
.A2(n_139),
.B(n_140),
.Y(n_1913)
);

O2A1O1Ixp5_ASAP7_75t_L g1914 ( 
.A1(n_1532),
.A2(n_298),
.B(n_377),
.C(n_373),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1636),
.B(n_141),
.Y(n_1915)
);

AOI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1745),
.A2(n_276),
.B(n_371),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1561),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1626),
.A2(n_142),
.B(n_144),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1579),
.B(n_142),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1606),
.A2(n_1589),
.B1(n_1607),
.B2(n_1605),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1639),
.A2(n_1679),
.B(n_1589),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1607),
.B(n_144),
.Y(n_1922)
);

NAND2x1p5_ASAP7_75t_L g1923 ( 
.A(n_1714),
.B(n_145),
.Y(n_1923)
);

AO31x2_ASAP7_75t_L g1924 ( 
.A1(n_1689),
.A2(n_145),
.A3(n_146),
.B(n_148),
.Y(n_1924)
);

AOI31xp67_ASAP7_75t_L g1925 ( 
.A1(n_1747),
.A2(n_396),
.A3(n_274),
.B(n_299),
.Y(n_1925)
);

AO31x2_ASAP7_75t_L g1926 ( 
.A1(n_1689),
.A2(n_148),
.A3(n_149),
.B(n_150),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1595),
.B(n_151),
.Y(n_1927)
);

AO31x2_ASAP7_75t_L g1928 ( 
.A1(n_1653),
.A2(n_151),
.A3(n_153),
.B(n_154),
.Y(n_1928)
);

AO32x2_ASAP7_75t_L g1929 ( 
.A1(n_1596),
.A2(n_153),
.A3(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1654),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1679),
.A2(n_304),
.B(n_360),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1558),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1679),
.A2(n_303),
.B(n_359),
.Y(n_1933)
);

AO31x2_ASAP7_75t_L g1934 ( 
.A1(n_1653),
.A2(n_158),
.A3(n_159),
.B(n_160),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1645),
.B(n_158),
.Y(n_1935)
);

INVxp67_ASAP7_75t_SL g1936 ( 
.A(n_1559),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1559),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_1937)
);

AO21x1_ASAP7_75t_L g1938 ( 
.A1(n_1756),
.A2(n_163),
.B(n_164),
.Y(n_1938)
);

NAND2xp33_ASAP7_75t_L g1939 ( 
.A(n_1732),
.B(n_163),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1605),
.A2(n_1549),
.B1(n_1703),
.B2(n_1750),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1666),
.A2(n_306),
.B(n_358),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_SL g1942 ( 
.A1(n_1547),
.A2(n_1554),
.B(n_1619),
.Y(n_1942)
);

BUFx10_ASAP7_75t_L g1943 ( 
.A(n_1546),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1656),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1714),
.B(n_165),
.Y(n_1945)
);

A2O1A1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1730),
.A2(n_165),
.B(n_166),
.C(n_167),
.Y(n_1946)
);

AND2x2_ASAP7_75t_SL g1947 ( 
.A(n_1652),
.B(n_167),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1661),
.A2(n_1662),
.B(n_1682),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1736),
.B(n_169),
.Y(n_1949)
);

BUFx12f_ASAP7_75t_L g1950 ( 
.A(n_1588),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1648),
.B(n_169),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1666),
.A2(n_312),
.B(n_357),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1703),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1710),
.A2(n_313),
.B(n_353),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1721),
.B(n_172),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1624),
.B(n_173),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1661),
.A2(n_315),
.B(n_351),
.Y(n_1957)
);

AO21x2_ASAP7_75t_L g1958 ( 
.A1(n_1779),
.A2(n_1524),
.B(n_1543),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1920),
.A2(n_1790),
.B(n_1894),
.C(n_1776),
.Y(n_1959)
);

OAI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1798),
.A2(n_1662),
.B(n_1599),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1908),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1948),
.A2(n_1705),
.B(n_1682),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1833),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_SL g1964 ( 
.A1(n_1947),
.A2(n_1724),
.B1(n_1701),
.B2(n_1690),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_L g1965 ( 
.A(n_1824),
.B(n_1602),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1810),
.Y(n_1966)
);

A2O1A1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1920),
.A2(n_1730),
.B(n_1692),
.C(n_1697),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1796),
.B(n_1614),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1811),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1773),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1787),
.A2(n_1552),
.B(n_1548),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_SL g1972 ( 
.A1(n_1894),
.A2(n_1942),
.B(n_1825),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1823),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1881),
.A2(n_1710),
.B(n_1687),
.Y(n_1974)
);

OAI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1845),
.A2(n_1583),
.B(n_1564),
.Y(n_1975)
);

OA21x2_ASAP7_75t_L g1976 ( 
.A1(n_1781),
.A2(n_1543),
.B(n_1692),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1815),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1860),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1833),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1799),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1834),
.Y(n_1981)
);

OAI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1846),
.A2(n_1603),
.B(n_1586),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1866),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1849),
.A2(n_1723),
.B1(n_1704),
.B2(n_1624),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1925),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1851),
.B(n_1645),
.Y(n_1986)
);

AOI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1940),
.A2(n_1663),
.B(n_1761),
.Y(n_1987)
);

OA21x2_ASAP7_75t_L g1988 ( 
.A1(n_1785),
.A2(n_1697),
.B(n_1755),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1886),
.B(n_1660),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1820),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1805),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1817),
.A2(n_1540),
.B1(n_1565),
.B2(n_1720),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1847),
.A2(n_1699),
.B(n_1660),
.Y(n_1993)
);

OAI21x1_ASAP7_75t_SL g1994 ( 
.A1(n_1825),
.A2(n_1718),
.B(n_1698),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1817),
.A2(n_1720),
.B1(n_1772),
.B2(n_1738),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1896),
.A2(n_1635),
.B(n_1678),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1897),
.A2(n_1592),
.B(n_1669),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1822),
.A2(n_1630),
.B1(n_1668),
.B2(n_1657),
.C(n_1667),
.Y(n_1998)
);

BUFx12f_ASAP7_75t_L g1999 ( 
.A(n_1943),
.Y(n_1999)
);

OA21x2_ASAP7_75t_L g2000 ( 
.A1(n_1784),
.A2(n_1755),
.B(n_1747),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1911),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1829),
.Y(n_2002)
);

OAI21x1_ASAP7_75t_L g2003 ( 
.A1(n_1921),
.A2(n_1604),
.B(n_1634),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1775),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1872),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1790),
.A2(n_1728),
.B(n_1633),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1878),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1840),
.B(n_1752),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1776),
.A2(n_1728),
.B(n_1737),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1778),
.A2(n_1632),
.B1(n_1770),
.B2(n_1734),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_SL g2011 ( 
.A1(n_1913),
.A2(n_1698),
.B(n_1670),
.Y(n_2011)
);

OAI21x1_ASAP7_75t_L g2012 ( 
.A1(n_1852),
.A2(n_1608),
.B(n_1609),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1880),
.Y(n_2013)
);

AO31x2_ASAP7_75t_L g2014 ( 
.A1(n_1940),
.A2(n_1650),
.A3(n_1545),
.B(n_1671),
.Y(n_2014)
);

OA21x2_ASAP7_75t_L g2015 ( 
.A1(n_1784),
.A2(n_1816),
.B(n_1791),
.Y(n_2015)
);

AOI21xp33_ASAP7_75t_L g2016 ( 
.A1(n_1788),
.A2(n_1726),
.B(n_1769),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_L g2017 ( 
.A(n_1906),
.B(n_1759),
.C(n_1758),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1853),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1855),
.Y(n_2019)
);

OAI21x1_ASAP7_75t_L g2020 ( 
.A1(n_1864),
.A2(n_1578),
.B(n_1609),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1777),
.B(n_1622),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1783),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1883),
.B(n_1651),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1884),
.A2(n_1738),
.B1(n_1694),
.B2(n_1733),
.Y(n_2024)
);

NAND2xp33_ASAP7_75t_SL g2025 ( 
.A(n_1849),
.B(n_1850),
.Y(n_2025)
);

CKINVDCx8_ASAP7_75t_R g2026 ( 
.A(n_1871),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_1946),
.B(n_1628),
.C(n_1716),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1866),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1850),
.A2(n_1706),
.B1(n_1702),
.B2(n_1670),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1812),
.A2(n_1712),
.B1(n_1587),
.B2(n_1769),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1830),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1807),
.B(n_1809),
.Y(n_2032)
);

OAI21x1_ASAP7_75t_L g2033 ( 
.A1(n_1957),
.A2(n_1608),
.B(n_1620),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1811),
.Y(n_2034)
);

BUFx2_ASAP7_75t_SL g2035 ( 
.A(n_1805),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1792),
.A2(n_1868),
.B(n_1789),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1893),
.Y(n_2037)
);

OAI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1889),
.A2(n_1674),
.B(n_1640),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1910),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1916),
.A2(n_1629),
.B(n_1670),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_1910),
.Y(n_2041)
);

OAI21x1_ASAP7_75t_L g2042 ( 
.A1(n_1891),
.A2(n_1618),
.B(n_1670),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1857),
.A2(n_1587),
.B1(n_1769),
.B2(n_1716),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_1857),
.A2(n_1716),
.B1(n_1600),
.B2(n_1706),
.Y(n_2044)
);

OAI21x1_ASAP7_75t_L g2045 ( 
.A1(n_1873),
.A2(n_1879),
.B(n_1837),
.Y(n_2045)
);

AO21x2_ASAP7_75t_L g2046 ( 
.A1(n_1789),
.A2(n_1816),
.B(n_1883),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1811),
.Y(n_2047)
);

OAI21x1_ASAP7_75t_L g2048 ( 
.A1(n_1839),
.A2(n_1651),
.B(n_1698),
.Y(n_2048)
);

OAI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1842),
.A2(n_1651),
.B(n_1698),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1930),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1814),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1944),
.Y(n_2052)
);

NAND2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1917),
.B(n_1659),
.Y(n_2053)
);

A2O1A1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1913),
.A2(n_1764),
.B(n_1651),
.C(n_1573),
.Y(n_2054)
);

AO21x2_ASAP7_75t_L g2055 ( 
.A1(n_1861),
.A2(n_1877),
.B(n_1794),
.Y(n_2055)
);

OAI21x1_ASAP7_75t_L g2056 ( 
.A1(n_1801),
.A2(n_1618),
.B(n_1739),
.Y(n_2056)
);

INVx4_ASAP7_75t_L g2057 ( 
.A(n_1917),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1922),
.A2(n_1888),
.B1(n_1923),
.B2(n_1806),
.Y(n_2058)
);

O2A1O1Ixp33_ASAP7_75t_L g2059 ( 
.A1(n_1774),
.A2(n_1717),
.B(n_1702),
.C(n_1706),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1888),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_SL g2061 ( 
.A1(n_1923),
.A2(n_1702),
.B(n_1732),
.Y(n_2061)
);

OA21x2_ASAP7_75t_L g2062 ( 
.A1(n_1835),
.A2(n_1771),
.B(n_1766),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_SL g2063 ( 
.A(n_1943),
.B(n_1573),
.Y(n_2063)
);

OAI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1818),
.A2(n_1757),
.B(n_1763),
.Y(n_2064)
);

AO21x2_ASAP7_75t_L g2065 ( 
.A1(n_1892),
.A2(n_1649),
.B(n_1771),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1819),
.A2(n_1600),
.B1(n_1717),
.B2(n_1527),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1780),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1964),
.A2(n_1819),
.B1(n_1870),
.B2(n_1862),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1984),
.A2(n_1870),
.B1(n_1862),
.B2(n_1937),
.Y(n_2069)
);

OAI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1995),
.A2(n_1937),
.B1(n_1953),
.B2(n_1918),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2025),
.A2(n_1912),
.B1(n_1919),
.B2(n_1895),
.Y(n_2071)
);

NAND2x1p5_ASAP7_75t_L g2072 ( 
.A(n_2060),
.B(n_1780),
.Y(n_2072)
);

INVx5_ASAP7_75t_L g2073 ( 
.A(n_2060),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2067),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2032),
.B(n_1966),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1970),
.B(n_2004),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_1999),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2025),
.A2(n_1949),
.B1(n_1956),
.B2(n_1803),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_R g2079 ( 
.A(n_1990),
.B(n_1956),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2001),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_2057),
.B(n_1848),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1968),
.B(n_1875),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_2031),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2008),
.B(n_1935),
.Y(n_2084)
);

OR2x6_ASAP7_75t_L g2085 ( 
.A(n_2061),
.B(n_1854),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1973),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1978),
.Y(n_2087)
);

OAI21x1_ASAP7_75t_L g2088 ( 
.A1(n_2056),
.A2(n_1899),
.B(n_1902),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2005),
.B(n_1822),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_L g2090 ( 
.A(n_1965),
.B(n_1953),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_2057),
.Y(n_2091)
);

CKINVDCx11_ASAP7_75t_R g2092 ( 
.A(n_1999),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_1990),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2007),
.Y(n_2094)
);

CKINVDCx20_ASAP7_75t_R g2095 ( 
.A(n_1981),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1986),
.B(n_1903),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_2058),
.B(n_1938),
.Y(n_2097)
);

NAND2xp33_ASAP7_75t_R g2098 ( 
.A(n_1980),
.B(n_1821),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2001),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_1989),
.A2(n_1874),
.B1(n_1826),
.B2(n_1918),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2021),
.B(n_1782),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2010),
.A2(n_2041),
.B1(n_1998),
.B2(n_2024),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1981),
.Y(n_2103)
);

CKINVDCx11_ASAP7_75t_R g2104 ( 
.A(n_2026),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2013),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1969),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2050),
.B(n_1922),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2039),
.A2(n_1826),
.B1(n_1885),
.B2(n_1838),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2035),
.B(n_1782),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2052),
.B(n_1836),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_2009),
.A2(n_1865),
.B1(n_1838),
.B2(n_1876),
.Y(n_2111)
);

AND2x6_ASAP7_75t_SL g2112 ( 
.A(n_1980),
.B(n_1950),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2022),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_1977),
.Y(n_2114)
);

OAI22xp5_ASAP7_75t_SL g2115 ( 
.A1(n_2030),
.A2(n_1797),
.B1(n_1887),
.B2(n_1865),
.Y(n_2115)
);

INVx11_ASAP7_75t_L g2116 ( 
.A(n_2063),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2002),
.Y(n_2117)
);

INVx3_ASAP7_75t_L g2118 ( 
.A(n_2057),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_2006),
.A2(n_1885),
.B1(n_1876),
.B2(n_1786),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2018),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1992),
.B(n_1804),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2053),
.Y(n_2122)
);

NAND2xp33_ASAP7_75t_R g2123 ( 
.A(n_1988),
.B(n_1900),
.Y(n_2123)
);

OR2x2_ASAP7_75t_SL g2124 ( 
.A(n_1976),
.B(n_1900),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2014),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_2053),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2002),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_1991),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2019),
.B(n_1863),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_2037),
.B(n_1863),
.Y(n_2130)
);

AO31x2_ASAP7_75t_L g2131 ( 
.A1(n_2036),
.A2(n_1844),
.A3(n_1828),
.B(n_1813),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2066),
.A2(n_1827),
.B1(n_1797),
.B2(n_1892),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2024),
.A2(n_1951),
.B1(n_1955),
.B2(n_1859),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_2066),
.A2(n_1797),
.B1(n_1945),
.B2(n_1907),
.Y(n_2134)
);

NAND2xp33_ASAP7_75t_R g2135 ( 
.A(n_1988),
.B(n_1909),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_1972),
.A2(n_1927),
.B1(n_1909),
.B2(n_1858),
.Y(n_2136)
);

BUFx2_ASAP7_75t_L g2137 ( 
.A(n_1983),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_1959),
.B(n_1936),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_1983),
.B(n_1843),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_2028),
.Y(n_2140)
);

HB1xp67_ASAP7_75t_L g2141 ( 
.A(n_2014),
.Y(n_2141)
);

OAI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2029),
.A2(n_1831),
.B1(n_1841),
.B2(n_1898),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2017),
.Y(n_2143)
);

INVx4_ASAP7_75t_SL g2144 ( 
.A(n_2014),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_SL g2145 ( 
.A1(n_1993),
.A2(n_2065),
.B1(n_1988),
.B2(n_1976),
.Y(n_2145)
);

AOI221xp5_ASAP7_75t_L g2146 ( 
.A1(n_1959),
.A2(n_1905),
.B1(n_1915),
.B2(n_1890),
.C(n_1904),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_1963),
.A2(n_1939),
.B(n_1882),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2086),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_SL g2149 ( 
.A1(n_2068),
.A2(n_2065),
.B1(n_1994),
.B2(n_2011),
.Y(n_2149)
);

AOI33xp33_ASAP7_75t_L g2150 ( 
.A1(n_2082),
.A2(n_2070),
.A3(n_2071),
.B1(n_2119),
.B2(n_2111),
.B3(n_2096),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2069),
.A2(n_2030),
.B1(n_2044),
.B2(n_2043),
.Y(n_2151)
);

OAI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2078),
.A2(n_1987),
.B1(n_2064),
.B2(n_2027),
.Y(n_2152)
);

OAI211xp5_ASAP7_75t_SL g2153 ( 
.A1(n_2102),
.A2(n_1967),
.B(n_2016),
.C(n_2044),
.Y(n_2153)
);

OAI211xp5_ASAP7_75t_L g2154 ( 
.A1(n_2090),
.A2(n_1967),
.B(n_2043),
.C(n_2059),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2084),
.B(n_2014),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_2070),
.A2(n_2055),
.B1(n_2023),
.B2(n_1976),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_2093),
.B(n_2028),
.Y(n_2157)
);

INVx5_ASAP7_75t_SL g2158 ( 
.A(n_2116),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2074),
.Y(n_2159)
);

OAI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_2079),
.A2(n_2023),
.B1(n_2000),
.B2(n_2015),
.Y(n_2160)
);

INVx2_ASAP7_75t_SL g2161 ( 
.A(n_2103),
.Y(n_2161)
);

AOI22xp33_ASAP7_75t_L g2162 ( 
.A1(n_2115),
.A2(n_2055),
.B1(n_2046),
.B2(n_1958),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_SL g2163 ( 
.A1(n_2091),
.A2(n_2046),
.B1(n_2062),
.B2(n_2000),
.Y(n_2163)
);

OAI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2132),
.A2(n_2054),
.B1(n_1795),
.B2(n_2062),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2121),
.A2(n_1958),
.B1(n_2062),
.B2(n_2015),
.Y(n_2165)
);

AOI221xp5_ASAP7_75t_L g2166 ( 
.A1(n_2089),
.A2(n_2108),
.B1(n_2142),
.B2(n_2071),
.C(n_2146),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2119),
.A2(n_2054),
.B1(n_2034),
.B2(n_2051),
.Y(n_2167)
);

INVxp67_ASAP7_75t_L g2168 ( 
.A(n_2083),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2147),
.A2(n_2108),
.B(n_2097),
.Y(n_2169)
);

BUFx4f_ASAP7_75t_SL g2170 ( 
.A(n_2095),
.Y(n_2170)
);

AOI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2138),
.A2(n_2015),
.B1(n_2000),
.B2(n_1793),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2117),
.Y(n_2172)
);

NOR2xp67_ASAP7_75t_L g2173 ( 
.A(n_2091),
.B(n_174),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_2138),
.A2(n_1808),
.B1(n_1800),
.B2(n_1763),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2111),
.A2(n_2051),
.B1(n_2034),
.B2(n_2047),
.Y(n_2175)
);

CKINVDCx6p67_ASAP7_75t_R g2176 ( 
.A(n_2104),
.Y(n_2176)
);

CKINVDCx20_ASAP7_75t_R g2177 ( 
.A(n_2092),
.Y(n_2177)
);

AOI22xp33_ASAP7_75t_L g2178 ( 
.A1(n_2146),
.A2(n_1757),
.B1(n_1754),
.B2(n_1766),
.Y(n_2178)
);

INVxp67_ASAP7_75t_L g2179 ( 
.A(n_2098),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_SL g2180 ( 
.A1(n_2118),
.A2(n_1969),
.B1(n_2047),
.B2(n_1996),
.Y(n_2180)
);

OAI211xp5_ASAP7_75t_L g2181 ( 
.A1(n_2145),
.A2(n_2134),
.B(n_2133),
.C(n_2100),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_2112),
.Y(n_2182)
);

AND2x4_ASAP7_75t_L g2183 ( 
.A(n_2118),
.B(n_1836),
.Y(n_2183)
);

OA21x2_ASAP7_75t_L g2184 ( 
.A1(n_2136),
.A2(n_2056),
.B(n_1985),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2120),
.B(n_1836),
.Y(n_2185)
);

OAI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2073),
.A2(n_1739),
.B1(n_1961),
.B2(n_1929),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2142),
.A2(n_1754),
.B1(n_1527),
.B2(n_1974),
.Y(n_2187)
);

OA21x2_ASAP7_75t_L g2188 ( 
.A1(n_2136),
.A2(n_1985),
.B(n_2038),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2107),
.A2(n_2075),
.B1(n_2139),
.B2(n_2094),
.C(n_2105),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2101),
.A2(n_1683),
.B1(n_1615),
.B2(n_1611),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2100),
.A2(n_1931),
.B1(n_1933),
.B2(n_1856),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2127),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2074),
.A2(n_1952),
.B1(n_1941),
.B2(n_1869),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2073),
.A2(n_2085),
.B1(n_2126),
.B2(n_2122),
.Y(n_2194)
);

AO31x2_ASAP7_75t_L g2195 ( 
.A1(n_2143),
.A2(n_1963),
.A3(n_1979),
.B(n_1961),
.Y(n_2195)
);

AOI221xp5_ASAP7_75t_L g2196 ( 
.A1(n_2087),
.A2(n_1867),
.B1(n_1832),
.B2(n_1914),
.C(n_1954),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2189),
.B(n_2076),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2148),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_2183),
.B(n_2144),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2159),
.B(n_2110),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2195),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2195),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2172),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2192),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2183),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2185),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2195),
.Y(n_2207)
);

INVxp67_ASAP7_75t_SL g2208 ( 
.A(n_2159),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2155),
.B(n_2125),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2166),
.B(n_2150),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2195),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2168),
.B(n_2113),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2184),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_2161),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2171),
.B(n_2125),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2184),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2184),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2175),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2167),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2151),
.B(n_2181),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_2194),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2156),
.B(n_2141),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2169),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2149),
.B(n_2129),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_2220),
.A2(n_2153),
.B1(n_2179),
.B2(n_2152),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2223),
.A2(n_2152),
.B(n_2186),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_2199),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_2210),
.A2(n_2158),
.B1(n_2164),
.B2(n_2160),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2198),
.Y(n_2229)
);

AOI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2197),
.A2(n_2160),
.B1(n_2154),
.B2(n_2162),
.C(n_2130),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_2214),
.Y(n_2231)
);

NAND5xp2_ASAP7_75t_SL g2232 ( 
.A(n_2215),
.B(n_2182),
.C(n_2077),
.D(n_2176),
.E(n_2158),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2198),
.Y(n_2233)
);

OAI31xp33_ASAP7_75t_SL g2234 ( 
.A1(n_2208),
.A2(n_2186),
.A3(n_2157),
.B(n_2081),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2209),
.B(n_2141),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2200),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2200),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2219),
.B(n_2206),
.Y(n_2238)
);

OAI31xp33_ASAP7_75t_L g2239 ( 
.A1(n_2221),
.A2(n_2191),
.A3(n_2114),
.B(n_2109),
.Y(n_2239)
);

OAI222xp33_ASAP7_75t_L g2240 ( 
.A1(n_2221),
.A2(n_2145),
.B1(n_2170),
.B2(n_2177),
.C1(n_2163),
.C2(n_2085),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2212),
.Y(n_2241)
);

NAND4xp25_ASAP7_75t_L g2242 ( 
.A(n_2224),
.B(n_2187),
.C(n_2174),
.D(n_2173),
.Y(n_2242)
);

OR2x6_ASAP7_75t_L g2243 ( 
.A(n_2199),
.B(n_2085),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2209),
.B(n_2080),
.Y(n_2244)
);

OAI21x1_ASAP7_75t_L g2245 ( 
.A1(n_2213),
.A2(n_2165),
.B(n_2188),
.Y(n_2245)
);

AO21x2_ASAP7_75t_L g2246 ( 
.A1(n_2223),
.A2(n_2147),
.B(n_2038),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2214),
.A2(n_2158),
.B1(n_2190),
.B2(n_2170),
.Y(n_2247)
);

AOI22xp33_ASAP7_75t_L g2248 ( 
.A1(n_2219),
.A2(n_2128),
.B1(n_2178),
.B2(n_2137),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2236),
.Y(n_2249)
);

NAND3xp33_ASAP7_75t_SL g2250 ( 
.A(n_2225),
.B(n_2072),
.C(n_2180),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2227),
.B(n_2199),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2237),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2227),
.B(n_2205),
.Y(n_2253)
);

NOR2xp67_ASAP7_75t_L g2254 ( 
.A(n_2227),
.B(n_2226),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2229),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2233),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2238),
.Y(n_2257)
);

INVx4_ASAP7_75t_L g2258 ( 
.A(n_2243),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2241),
.B(n_2206),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2235),
.B(n_2218),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2245),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_2231),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2245),
.B(n_2205),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2240),
.A2(n_2199),
.B(n_2081),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2246),
.B(n_2215),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2246),
.B(n_2218),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2230),
.B(n_2203),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_2243),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2246),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2243),
.B(n_2213),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2243),
.B(n_2216),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2244),
.B(n_2216),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_2228),
.B(n_2217),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2228),
.B(n_2217),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2259),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2263),
.B(n_2234),
.Y(n_2276)
);

INVxp67_ASAP7_75t_L g2277 ( 
.A(n_2262),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2259),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2261),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2267),
.B(n_2225),
.Y(n_2280)
);

AND2x4_ASAP7_75t_SL g2281 ( 
.A(n_2258),
.B(n_2126),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2267),
.B(n_2239),
.Y(n_2282)
);

NAND2x1p5_ASAP7_75t_L g2283 ( 
.A(n_2258),
.B(n_2214),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2261),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_2260),
.B(n_2222),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2261),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2263),
.B(n_2222),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2259),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2275),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2283),
.B(n_2277),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2283),
.B(n_2258),
.Y(n_2291)
);

NOR2xp67_ASAP7_75t_L g2292 ( 
.A(n_2276),
.B(n_2258),
.Y(n_2292)
);

NOR3xp33_ASAP7_75t_L g2293 ( 
.A(n_2280),
.B(n_2250),
.C(n_2258),
.Y(n_2293)
);

AOI32xp33_ASAP7_75t_L g2294 ( 
.A1(n_2276),
.A2(n_2274),
.A3(n_2273),
.B1(n_2268),
.B2(n_2265),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2278),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2285),
.B(n_2260),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2281),
.B(n_2268),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2288),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2282),
.B(n_2257),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2285),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2279),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2287),
.B(n_2266),
.Y(n_2302)
);

NOR2x1_ASAP7_75t_L g2303 ( 
.A(n_2287),
.B(n_2250),
.Y(n_2303)
);

OR2x2_ASAP7_75t_L g2304 ( 
.A(n_2283),
.B(n_2266),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2300),
.Y(n_2305)
);

OAI32xp33_ASAP7_75t_L g2306 ( 
.A1(n_2293),
.A2(n_2268),
.A3(n_2262),
.B1(n_2274),
.B2(n_2247),
.Y(n_2306)
);

AOI221xp5_ASAP7_75t_L g2307 ( 
.A1(n_2294),
.A2(n_2266),
.B1(n_2265),
.B2(n_2232),
.C(n_2273),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_L g2308 ( 
.A1(n_2293),
.A2(n_2299),
.B1(n_2303),
.B2(n_2292),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2299),
.A2(n_2265),
.B1(n_2273),
.B2(n_2274),
.C(n_2263),
.Y(n_2309)
);

AOI21xp33_ASAP7_75t_SL g2310 ( 
.A1(n_2291),
.A2(n_2273),
.B(n_2251),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2296),
.Y(n_2311)
);

OAI221xp5_ASAP7_75t_L g2312 ( 
.A1(n_2304),
.A2(n_2254),
.B1(n_2264),
.B2(n_2268),
.C(n_2262),
.Y(n_2312)
);

AOI222xp33_ASAP7_75t_SL g2313 ( 
.A1(n_2289),
.A2(n_2286),
.B1(n_2284),
.B2(n_2279),
.C1(n_2257),
.C2(n_2252),
.Y(n_2313)
);

NAND3xp33_ASAP7_75t_L g2314 ( 
.A(n_2290),
.B(n_2254),
.C(n_2284),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2295),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2297),
.A2(n_2264),
.B(n_2281),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2311),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2305),
.B(n_2302),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2308),
.A2(n_2297),
.B1(n_2298),
.B2(n_2262),
.Y(n_2319)
);

AOI221x1_ASAP7_75t_L g2320 ( 
.A1(n_2316),
.A2(n_2301),
.B1(n_2286),
.B2(n_2273),
.C(n_2269),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2315),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2306),
.B(n_2249),
.Y(n_2322)
);

AOI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2307),
.A2(n_2242),
.B1(n_2301),
.B2(n_2248),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2314),
.Y(n_2324)
);

AOI322xp5_ASAP7_75t_L g2325 ( 
.A1(n_2308),
.A2(n_2251),
.A3(n_2253),
.B1(n_2249),
.B2(n_2252),
.C1(n_2248),
.C2(n_2270),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2312),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2313),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2326),
.B(n_2310),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2317),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2318),
.Y(n_2330)
);

OR2x2_ASAP7_75t_L g2331 ( 
.A(n_2324),
.B(n_2255),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2327),
.B(n_2309),
.Y(n_2332)
);

INVxp33_ASAP7_75t_L g2333 ( 
.A(n_2319),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2321),
.Y(n_2334)
);

NAND3xp33_ASAP7_75t_L g2335 ( 
.A(n_2323),
.B(n_2269),
.C(n_2255),
.Y(n_2335)
);

INVx1_ASAP7_75t_SL g2336 ( 
.A(n_2323),
.Y(n_2336)
);

XNOR2xp5_ASAP7_75t_L g2337 ( 
.A(n_2320),
.B(n_2251),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2322),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2325),
.B(n_2256),
.Y(n_2339)
);

OAI221xp5_ASAP7_75t_L g2340 ( 
.A1(n_2323),
.A2(n_2269),
.B1(n_2271),
.B2(n_2270),
.C(n_2253),
.Y(n_2340)
);

XOR2x2_ASAP7_75t_L g2341 ( 
.A(n_2336),
.B(n_2251),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2333),
.B(n_2251),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2330),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2336),
.A2(n_2269),
.B(n_2256),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2332),
.B(n_2253),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2329),
.Y(n_2346)
);

NOR3xp33_ASAP7_75t_SL g2347 ( 
.A(n_2338),
.B(n_2135),
.C(n_2123),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2328),
.A2(n_2271),
.B(n_2270),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2334),
.B(n_2271),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_L g2350 ( 
.A(n_2335),
.B(n_2073),
.C(n_2196),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2331),
.B(n_2272),
.Y(n_2351)
);

AOI221xp5_ASAP7_75t_L g2352 ( 
.A1(n_2346),
.A2(n_2340),
.B1(n_2339),
.B2(n_2337),
.C(n_2272),
.Y(n_2352)
);

AOI221xp5_ASAP7_75t_L g2353 ( 
.A1(n_2343),
.A2(n_2339),
.B1(n_2272),
.B2(n_2140),
.C(n_2211),
.Y(n_2353)
);

AOI222xp33_ASAP7_75t_L g2354 ( 
.A1(n_2341),
.A2(n_2211),
.B1(n_2073),
.B2(n_2217),
.C1(n_2144),
.C2(n_2201),
.Y(n_2354)
);

AOI221xp5_ASAP7_75t_L g2355 ( 
.A1(n_2345),
.A2(n_2140),
.B1(n_2193),
.B2(n_2203),
.C(n_2204),
.Y(n_2355)
);

A2O1A1Ixp33_ASAP7_75t_L g2356 ( 
.A1(n_2342),
.A2(n_2204),
.B(n_2202),
.C(n_2201),
.Y(n_2356)
);

AOI222xp33_ASAP7_75t_L g2357 ( 
.A1(n_2349),
.A2(n_2350),
.B1(n_2351),
.B2(n_2344),
.C1(n_2347),
.C2(n_2348),
.Y(n_2357)
);

AOI221xp5_ASAP7_75t_L g2358 ( 
.A1(n_2346),
.A2(n_2202),
.B1(n_2201),
.B2(n_2207),
.C(n_2072),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2346),
.B(n_1969),
.Y(n_2359)
);

AOI221xp5_ASAP7_75t_SL g2360 ( 
.A1(n_2343),
.A2(n_2124),
.B1(n_2202),
.B2(n_2207),
.C(n_1929),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2359),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2357),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2356),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2352),
.B(n_2353),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2360),
.B(n_1615),
.C(n_1611),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2355),
.B(n_2358),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_2354),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2357),
.A2(n_2106),
.B1(n_1969),
.B2(n_2188),
.Y(n_2368)
);

INVxp33_ASAP7_75t_L g2369 ( 
.A(n_2359),
.Y(n_2369)
);

AND4x1_ASAP7_75t_L g2370 ( 
.A(n_2362),
.B(n_174),
.C(n_175),
.D(n_176),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2364),
.B(n_175),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2361),
.B(n_2144),
.Y(n_2372)
);

NOR2x1p5_ASAP7_75t_L g2373 ( 
.A(n_2367),
.B(n_2106),
.Y(n_2373)
);

OR2x2_ASAP7_75t_L g2374 ( 
.A(n_2363),
.B(n_2368),
.Y(n_2374)
);

OAI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2368),
.A2(n_2188),
.B1(n_2099),
.B2(n_2106),
.Y(n_2375)
);

AOI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2369),
.A2(n_1814),
.B1(n_1932),
.B2(n_1929),
.C(n_1739),
.Y(n_2376)
);

XNOR2x1_ASAP7_75t_L g2377 ( 
.A(n_2365),
.B(n_262),
.Y(n_2377)
);

AOI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_2366),
.A2(n_1814),
.B1(n_1932),
.B2(n_1665),
.Y(n_2378)
);

AOI322xp5_ASAP7_75t_L g2379 ( 
.A1(n_2362),
.A2(n_1901),
.A3(n_1926),
.B1(n_1924),
.B2(n_1928),
.C1(n_1934),
.C2(n_1979),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2371),
.A2(n_1932),
.B1(n_2040),
.B2(n_1665),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2373),
.A2(n_1996),
.B1(n_1962),
.B2(n_2040),
.Y(n_2381)
);

AOI21xp33_ASAP7_75t_L g2382 ( 
.A1(n_2374),
.A2(n_263),
.B(n_264),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_SL g2383 ( 
.A1(n_2370),
.A2(n_1926),
.B1(n_1924),
.B2(n_1934),
.Y(n_2383)
);

AOI22xp5_ASAP7_75t_L g2384 ( 
.A1(n_2377),
.A2(n_2033),
.B1(n_2048),
.B2(n_2049),
.Y(n_2384)
);

NAND3xp33_ASAP7_75t_SL g2385 ( 
.A(n_2378),
.B(n_1926),
.C(n_1924),
.Y(n_2385)
);

AOI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_2372),
.A2(n_2033),
.B1(n_2048),
.B2(n_2049),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_2375),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2376),
.Y(n_2388)
);

NAND3xp33_ASAP7_75t_SL g2389 ( 
.A(n_2379),
.B(n_1934),
.C(n_1928),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_2388),
.B(n_1901),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2387),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2382),
.B(n_2380),
.Y(n_2392)
);

XNOR2xp5_ASAP7_75t_L g2393 ( 
.A(n_2383),
.B(n_266),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2389),
.A2(n_1997),
.B1(n_2012),
.B2(n_2020),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2384),
.A2(n_1618),
.B1(n_1901),
.B2(n_1928),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2385),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2386),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_2391),
.Y(n_2398)
);

OAI211xp5_ASAP7_75t_L g2399 ( 
.A1(n_2396),
.A2(n_2381),
.B(n_269),
.C(n_270),
.Y(n_2399)
);

OAI21xp5_ASAP7_75t_L g2400 ( 
.A1(n_2393),
.A2(n_1997),
.B(n_2012),
.Y(n_2400)
);

NAND3xp33_ASAP7_75t_L g2401 ( 
.A(n_2392),
.B(n_1760),
.C(n_1746),
.Y(n_2401)
);

INVx1_ASAP7_75t_SL g2402 ( 
.A(n_2397),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2390),
.Y(n_2403)
);

XNOR2xp5_ASAP7_75t_L g2404 ( 
.A(n_2402),
.B(n_2395),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2398),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2401),
.Y(n_2406)
);

AOI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2399),
.A2(n_2403),
.B1(n_2400),
.B2(n_2394),
.Y(n_2407)
);

BUFx4f_ASAP7_75t_SL g2408 ( 
.A(n_2405),
.Y(n_2408)
);

NAND2xp33_ASAP7_75t_SL g2409 ( 
.A(n_2404),
.B(n_1760),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2407),
.Y(n_2410)
);

XNOR2xp5_ASAP7_75t_L g2411 ( 
.A(n_2410),
.B(n_2406),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2408),
.B(n_267),
.Y(n_2412)
);

AOI222xp33_ASAP7_75t_L g2413 ( 
.A1(n_2411),
.A2(n_2409),
.B1(n_1746),
.B2(n_1760),
.C1(n_2020),
.C2(n_2088),
.Y(n_2413)
);

AOI222xp33_ASAP7_75t_L g2414 ( 
.A1(n_2413),
.A2(n_2412),
.B1(n_2045),
.B2(n_2003),
.C1(n_1982),
.C2(n_1975),
.Y(n_2414)
);

OAI221xp5_ASAP7_75t_R g2415 ( 
.A1(n_2414),
.A2(n_2131),
.B1(n_1802),
.B2(n_271),
.C(n_273),
.Y(n_2415)
);

AOI211xp5_ASAP7_75t_L g2416 ( 
.A1(n_2415),
.A2(n_2042),
.B(n_1971),
.C(n_1960),
.Y(n_2416)
);


endmodule