module fake_jpeg_4000_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_18),
.B1(n_28),
.B2(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_17),
.C(n_19),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_67),
.C(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_20),
.B1(n_33),
.B2(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_25),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_18),
.C(n_28),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_74),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_27),
.B1(n_32),
.B2(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_77),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_90),
.B1(n_93),
.B2(n_20),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_31),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_31),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_92),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_20),
.B1(n_33),
.B2(n_21),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_97),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_66),
.B1(n_53),
.B2(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_78),
.B1(n_82),
.B2(n_89),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_105),
.Y(n_144)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_44),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_60),
.B1(n_62),
.B2(n_51),
.Y(n_129)
);

AND2x4_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_39),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_68),
.B1(n_63),
.B2(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_93),
.B(n_74),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_22),
.B(n_26),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_74),
.B1(n_76),
.B2(n_86),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_49),
.B1(n_53),
.B2(n_45),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_47),
.B1(n_65),
.B2(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_87),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_109),
.B1(n_104),
.B2(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_145),
.B1(n_118),
.B2(n_119),
.Y(n_166)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_21),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_13),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_116),
.B1(n_83),
.B2(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_124),
.C(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_152),
.C(n_153),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_42),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_108),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_127),
.B(n_135),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_160),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_163),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_23),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_169),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_64),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_142),
.C(n_129),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_81),
.B(n_80),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_21),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_170),
.B(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_22),
.B1(n_26),
.B2(n_59),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_83),
.A3(n_89),
.B1(n_42),
.B2(n_50),
.C1(n_59),
.C2(n_33),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_133),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_173),
.B1(n_126),
.B2(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_106),
.B(n_50),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_130),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_186),
.B(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_180),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_190),
.B(n_16),
.Y(n_222)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_157),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_197),
.C(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_132),
.B1(n_130),
.B2(n_105),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_132),
.B1(n_117),
.B2(n_114),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_22),
.B1(n_26),
.B2(n_99),
.Y(n_223)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_139),
.B1(n_128),
.B2(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_151),
.B(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_128),
.C(n_12),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_163),
.C(n_161),
.Y(n_203)
);

XOR2x2_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_11),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_173),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_16),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_131),
.B1(n_26),
.B2(n_22),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_205),
.C(n_206),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_153),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_149),
.C(n_148),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_162),
.C(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_209),
.C(n_210),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_169),
.C(n_161),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_158),
.C(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_188),
.C(n_182),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.C(n_177),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_173),
.C(n_170),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_219),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_151),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_224),
.Y(n_229)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_184),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_193),
.B(n_178),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_196),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_232),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_190),
.B(n_199),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_242),
.B1(n_214),
.B2(n_217),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_204),
.C(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_238),
.C(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_175),
.C(n_194),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_198),
.B(n_200),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_210),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_115),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_157),
.C(n_113),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_0),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_229),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_220),
.C(n_213),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_257),
.C(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_215),
.C(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_2),
.C(n_3),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_238),
.B1(n_240),
.B2(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_275),
.B(n_253),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_276),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_232),
.B1(n_228),
.B2(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_248),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_278),
.C(n_253),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_241),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_277),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_226),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_285),
.C(n_272),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_284),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_249),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_286),
.B(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_259),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_9),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_269),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_9),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_10),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_9),
.B(n_12),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_8),
.B(n_11),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_299),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_15),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_291),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_297),
.B(n_298),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_300),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_4),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_10),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_288),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_280),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_307),
.A2(n_309),
.B(n_301),
.C(n_5),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_4),
.B(n_5),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_15),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_311),
.B(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_304),
.C(n_302),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_314),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_312),
.B(n_308),
.C(n_315),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_6),
.C(n_7),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_6),
.B1(n_7),
.B2(n_313),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_6),
.Y(n_320)
);


endmodule