module fake_netlist_1_6688_n_915 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_39, n_915);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_39;
output n_915;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g225 ( .A(n_43), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_105), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_54), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_60), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_67), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_138), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_217), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_100), .Y(n_234) );
INVxp33_ASAP7_75t_SL g235 ( .A(n_27), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_31), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_149), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_75), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_153), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_65), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_127), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_110), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_50), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_117), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_15), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_7), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_196), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_128), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_22), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_147), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_126), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g252 ( .A(n_216), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_72), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_152), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_63), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_181), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_56), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_36), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_135), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_143), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_18), .Y(n_261) );
INVxp33_ASAP7_75t_SL g262 ( .A(n_144), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_104), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_31), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_133), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_95), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_167), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_85), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_89), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_209), .B(n_132), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_198), .B(n_67), .Y(n_272) );
CKINVDCx16_ASAP7_75t_R g273 ( .A(n_72), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_45), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_139), .Y(n_275) );
CKINVDCx14_ASAP7_75t_R g276 ( .A(n_187), .Y(n_276) );
CKINVDCx16_ASAP7_75t_R g277 ( .A(n_66), .Y(n_277) );
BUFx2_ASAP7_75t_SL g278 ( .A(n_111), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_204), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_13), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_26), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_131), .Y(n_282) );
INVxp33_ASAP7_75t_L g283 ( .A(n_164), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_130), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_78), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_52), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_30), .Y(n_287) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_188), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_80), .Y(n_289) );
CKINVDCx16_ASAP7_75t_R g290 ( .A(n_68), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_118), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_218), .B(n_34), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_220), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_91), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_151), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_157), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_215), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_15), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_163), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_50), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_98), .Y(n_301) );
INVxp33_ASAP7_75t_SL g302 ( .A(n_65), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_9), .Y(n_303) );
INVxp33_ASAP7_75t_L g304 ( .A(n_44), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_185), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_81), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_186), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_120), .Y(n_308) );
CKINVDCx16_ASAP7_75t_R g309 ( .A(n_109), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_192), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_46), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g312 ( .A(n_175), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_71), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_90), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_222), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_55), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_173), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_5), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_79), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_61), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_115), .Y(n_321) );
INVxp33_ASAP7_75t_L g322 ( .A(n_178), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_146), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_161), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_77), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_189), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_205), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_199), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_124), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_207), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_180), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_99), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_158), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_86), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_73), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_169), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_184), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_34), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_62), .Y(n_339) );
INVxp33_ASAP7_75t_SL g340 ( .A(n_148), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_76), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_141), .Y(n_342) );
INVxp33_ASAP7_75t_SL g343 ( .A(n_123), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_59), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_197), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_125), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_108), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_232), .B(n_0), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_269), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_280), .Y(n_350) );
INVx4_ASAP7_75t_L g351 ( .A(n_272), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_269), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_280), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_253), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_253), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_304), .B(n_0), .Y(n_356) );
AND2x6_ASAP7_75t_L g357 ( .A(n_319), .B(n_74), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_269), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_269), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_272), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_279), .B(n_1), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_325), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_237), .B(n_1), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_344), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_301), .B(n_2), .Y(n_366) );
NAND2xp33_ASAP7_75t_L g367 ( .A(n_283), .B(n_224), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_309), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_272), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_321), .B(n_2), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_344), .B(n_319), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_278), .B(n_3), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_283), .B(n_3), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_226), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_312), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_246), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_304), .B(n_264), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_273), .B(n_4), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_228), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_277), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_345), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_375), .B(n_233), .C(n_231), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_351), .B(n_285), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_356), .A2(n_227), .B1(n_229), .B2(n_225), .Y(n_386) );
BUFx10_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_360), .B(n_230), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_351), .B(n_322), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_351), .B(n_322), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_378), .B(n_240), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_360), .B(n_236), .Y(n_393) );
XOR2xp5_ASAP7_75t_L g394 ( .A(n_381), .B(n_255), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_360), .B(n_240), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_360), .B(n_234), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_377), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_369), .B(n_258), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_349), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_349), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_369), .B(n_243), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_349), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_377), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_358), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_380), .B(n_244), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_380), .B(n_252), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_372), .B(n_252), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_358), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_372), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_352), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_372), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_354), .B(n_244), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_359), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_357), .Y(n_420) );
NAND3x1_ASAP7_75t_L g421 ( .A(n_379), .B(n_249), .C(n_245), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_373), .B(n_261), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_354), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_422), .A2(n_373), .B1(n_357), .B2(n_365), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_422), .B(n_373), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_410), .B(n_384), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_392), .B(n_290), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_386), .A2(n_373), .B1(n_242), .B2(n_330), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_410), .B(n_374), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_391), .B(n_348), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_423), .Y(n_435) );
AO21x1_ASAP7_75t_L g436 ( .A1(n_397), .A2(n_422), .B(n_418), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_394), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_422), .B(n_362), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_389), .B(n_366), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_423), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_397), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_413), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_423), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_408), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_411), .B(n_371), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_411), .B(n_373), .Y(n_447) );
OAI21xp33_ASAP7_75t_SL g448 ( .A1(n_395), .A2(n_365), .B(n_355), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_388), .B(n_364), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_401), .A2(n_255), .B1(n_300), .B2(n_257), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_415), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_408), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_387), .Y(n_453) );
INVx5_ASAP7_75t_L g454 ( .A(n_387), .Y(n_454) );
OR2x2_ASAP7_75t_SL g455 ( .A(n_403), .B(n_257), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_399), .B(n_382), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_388), .B(n_355), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_421), .A2(n_302), .B1(n_235), .B2(n_242), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_383), .A2(n_357), .B(n_367), .Y(n_462) );
OR2x6_ASAP7_75t_L g463 ( .A(n_401), .B(n_381), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_390), .B(n_238), .Y(n_464) );
INVx4_ASAP7_75t_L g465 ( .A(n_390), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_388), .B(n_350), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_409), .B(n_258), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_383), .B(n_353), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_397), .A2(n_330), .B1(n_333), .B2(n_324), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_390), .B(n_239), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_393), .Y(n_472) );
INVx4_ASAP7_75t_L g473 ( .A(n_393), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_419), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_418), .A2(n_338), .B1(n_286), .B2(n_320), .C(n_311), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_404), .B(n_353), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_394), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_420), .B(n_241), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_404), .B(n_247), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_404), .B(n_259), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_398), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_398), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_420), .B(n_262), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_407), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_407), .A2(n_271), .B(n_268), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_402), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_402), .B(n_300), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_402), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_406), .B(n_259), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_406), .Y(n_493) );
AND2x2_ASAP7_75t_SL g494 ( .A(n_385), .B(n_246), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_385), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_414), .A2(n_343), .B1(n_340), .B2(n_274), .Y(n_496) );
INVx4_ASAP7_75t_L g497 ( .A(n_454), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_426), .A2(n_343), .B1(n_287), .B2(n_298), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_428), .B(n_281), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_435), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_470), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_437), .A2(n_276), .B1(n_293), .B2(n_289), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_441), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_440), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_434), .A2(n_284), .B(n_270), .Y(n_507) );
NOR2xp33_ASAP7_75t_SL g508 ( .A(n_494), .B(n_357), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_427), .A2(n_337), .B(n_288), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_454), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_447), .A2(n_357), .B1(n_303), .B2(n_316), .Y(n_511) );
BUFx12f_ASAP7_75t_L g512 ( .A(n_455), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_468), .B(n_313), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_490), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_454), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_429), .B(n_318), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_443), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_479), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_443), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_463), .A2(n_296), .B1(n_310), .B2(n_307), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_424), .A2(n_339), .B1(n_292), .B2(n_250), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_438), .B(n_439), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_425), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_425), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_494), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_473), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_448), .A2(n_254), .B(n_256), .C(n_251), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_436), .B(n_357), .Y(n_531) );
INVx3_ASAP7_75t_SL g532 ( .A(n_463), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_449), .A2(n_357), .B1(n_263), .B2(n_265), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_480), .B(n_6), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_465), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_465), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_433), .B(n_357), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_444), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_446), .B(n_260), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_456), .B(n_248), .Y(n_541) );
CKINVDCx11_ASAP7_75t_R g542 ( .A(n_437), .Y(n_542) );
INVx4_ASAP7_75t_L g543 ( .A(n_453), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_424), .A2(n_275), .B(n_282), .C(n_267), .Y(n_544) );
OR2x6_ASAP7_75t_L g545 ( .A(n_474), .B(n_246), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_460), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_442), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_451), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_458), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_464), .A2(n_294), .B(n_291), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_464), .A2(n_297), .B(n_295), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_478), .A2(n_306), .B(n_314), .C(n_305), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_430), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_469), .A2(n_323), .B1(n_326), .B2(n_317), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_486), .A2(n_331), .B1(n_334), .B2(n_329), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_431), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_471), .A2(n_336), .B(n_335), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_486), .A2(n_496), .B1(n_482), .B2(n_483), .Y(n_558) );
INVx3_ASAP7_75t_L g559 ( .A(n_432), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_485), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_445), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_488), .A2(n_346), .B(n_347), .C(n_342), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_487), .B(n_308), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_452), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_459), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_459), .Y(n_566) );
OR2x6_ASAP7_75t_L g567 ( .A(n_462), .B(n_266), .Y(n_567) );
INVx5_ASAP7_75t_L g568 ( .A(n_461), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_467), .A2(n_299), .B(n_315), .C(n_268), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_484), .A2(n_341), .B1(n_315), .B2(n_327), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_475), .Y(n_571) );
INVx5_ASAP7_75t_L g572 ( .A(n_475), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_476), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_481), .A2(n_328), .B(n_299), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_477), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_492), .Y(n_576) );
CKINVDCx16_ASAP7_75t_R g577 ( .A(n_484), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_491), .Y(n_578) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_493), .Y(n_579) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_495), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_489), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_489), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_495), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_434), .A2(n_332), .B(n_417), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_470), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_472), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_426), .A2(n_359), .B1(n_363), .B2(n_325), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_577), .A2(n_359), .B1(n_363), .B2(n_361), .Y(n_588) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_531), .A2(n_363), .B(n_417), .Y(n_589) );
BUFx3_ASAP7_75t_L g590 ( .A(n_516), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_502), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_505), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_571), .Y(n_594) );
AO21x2_ASAP7_75t_L g595 ( .A1(n_531), .A2(n_361), .B(n_352), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_542), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_585), .A2(n_361), .B1(n_370), .B2(n_352), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_546), .A2(n_352), .B1(n_361), .B2(n_370), .C(n_10), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_560), .Y(n_600) );
OA21x2_ASAP7_75t_L g601 ( .A1(n_584), .A2(n_370), .B(n_361), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_497), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_512), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_538), .A2(n_396), .B(n_385), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_561), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_561), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_524), .A2(n_400), .B(n_396), .C(n_385), .Y(n_607) );
AO22x2_ASAP7_75t_L g608 ( .A1(n_523), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_499), .A2(n_400), .B1(n_396), .B2(n_385), .C(n_13), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_524), .A2(n_400), .B(n_396), .C(n_12), .Y(n_610) );
AO31x2_ASAP7_75t_L g611 ( .A1(n_569), .A2(n_8), .A3(n_11), .B(n_12), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_564), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_574), .A2(n_83), .B(n_82), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_565), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_566), .Y(n_615) );
INVx6_ASAP7_75t_L g616 ( .A(n_516), .Y(n_616) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_574), .A2(n_87), .B(n_84), .Y(n_617) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_523), .A2(n_11), .A3(n_14), .B(n_16), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_545), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_514), .A2(n_400), .B1(n_396), .B2(n_19), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_567), .A2(n_400), .B(n_396), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_567), .A2(n_400), .B(n_88), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_532), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_586), .Y(n_624) );
INVx5_ASAP7_75t_L g625 ( .A(n_497), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_575), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_517), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_503), .B(n_20), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_568), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_526), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_510), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_579), .Y(n_632) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_559), .A2(n_93), .B(n_92), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g634 ( .A(n_528), .B(n_94), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_558), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_579), .Y(n_636) );
OR2x6_ASAP7_75t_SL g637 ( .A(n_534), .B(n_25), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_510), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g639 ( .A1(n_545), .A2(n_26), .B(n_27), .Y(n_639) );
CKINVDCx16_ASAP7_75t_R g640 ( .A(n_504), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_498), .B(n_28), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_515), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_558), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_552), .A2(n_29), .B(n_32), .C(n_33), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_525), .Y(n_646) );
AO21x2_ASAP7_75t_L g647 ( .A1(n_530), .A2(n_97), .B(n_96), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_519), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_513), .A2(n_33), .B1(n_35), .B2(n_36), .Y(n_649) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_525), .Y(n_650) );
OR2x6_ASAP7_75t_L g651 ( .A(n_545), .B(n_35), .Y(n_651) );
OAI222xp33_ASAP7_75t_L g652 ( .A1(n_498), .A2(n_37), .B1(n_38), .B2(n_39), .C1(n_40), .C2(n_41), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_582), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_520), .B(n_540), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_528), .B(n_38), .Y(n_655) );
OAI21x1_ASAP7_75t_SL g656 ( .A1(n_543), .A2(n_39), .B(n_40), .Y(n_656) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_562), .A2(n_102), .B(n_101), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_547), .Y(n_658) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_553), .A2(n_145), .B(n_221), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_548), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_549), .Y(n_661) );
OAI21x1_ASAP7_75t_SL g662 ( .A1(n_543), .A2(n_42), .B(n_43), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_525), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_500), .Y(n_664) );
OA21x2_ASAP7_75t_L g665 ( .A1(n_544), .A2(n_150), .B(n_219), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_551), .A2(n_154), .B(n_214), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_527), .Y(n_667) );
OA21x2_ASAP7_75t_L g668 ( .A1(n_533), .A2(n_142), .B(n_213), .Y(n_668) );
OAI21x1_ASAP7_75t_L g669 ( .A1(n_581), .A2(n_140), .B(n_212), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_515), .Y(n_670) );
OAI21x1_ASAP7_75t_L g671 ( .A1(n_556), .A2(n_137), .B(n_211), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_529), .Y(n_672) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_527), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_508), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_674) );
OAI21x1_ASAP7_75t_L g675 ( .A1(n_506), .A2(n_155), .B(n_208), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_555), .A2(n_51), .B(n_52), .C(n_53), .Y(n_676) );
AOI21x1_ASAP7_75t_L g677 ( .A1(n_567), .A2(n_159), .B(n_206), .Y(n_677) );
OAI21x1_ASAP7_75t_L g678 ( .A1(n_518), .A2(n_539), .B(n_521), .Y(n_678) );
AO32x2_ASAP7_75t_L g679 ( .A1(n_554), .A2(n_57), .A3(n_58), .B1(n_59), .B2(n_60), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_568), .Y(n_680) );
AO21x2_ASAP7_75t_L g681 ( .A1(n_550), .A2(n_165), .B(n_203), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_537), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_572), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_507), .A2(n_509), .B(n_557), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_578), .A2(n_162), .B(n_202), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_541), .B(n_62), .Y(n_686) );
INVx6_ASAP7_75t_L g687 ( .A(n_572), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_527), .Y(n_688) );
INVx8_ASAP7_75t_L g689 ( .A(n_572), .Y(n_689) );
BUFx4f_ASAP7_75t_L g690 ( .A(n_528), .Y(n_690) );
OAI21x1_ASAP7_75t_L g691 ( .A1(n_587), .A2(n_168), .B(n_201), .Y(n_691) );
OAI21x1_ASAP7_75t_L g692 ( .A1(n_587), .A2(n_166), .B(n_200), .Y(n_692) );
AO21x2_ASAP7_75t_L g693 ( .A1(n_607), .A2(n_554), .B(n_509), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_651), .A2(n_576), .B1(n_570), .B2(n_511), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_684), .A2(n_563), .B(n_508), .C(n_535), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_592), .B(n_536), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_629), .Y(n_697) );
INVx3_ASAP7_75t_L g698 ( .A(n_689), .Y(n_698) );
AO21x2_ASAP7_75t_L g699 ( .A1(n_595), .A2(n_583), .B(n_580), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_655), .A2(n_64), .B1(n_66), .B2(n_69), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_652), .A2(n_69), .B(n_70), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_639), .A2(n_103), .B(n_106), .C(n_107), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_608), .A2(n_112), .B1(n_113), .B2(n_114), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_604), .A2(n_116), .B(n_119), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_594), .B(n_121), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_626), .B(n_122), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_676), .A2(n_129), .B(n_134), .C(n_136), .Y(n_707) );
AO22x2_ASAP7_75t_L g708 ( .A1(n_628), .A2(n_156), .B1(n_160), .B2(n_170), .Y(n_708) );
AO31x2_ASAP7_75t_L g709 ( .A1(n_610), .A2(n_171), .A3(n_172), .B(n_174), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_686), .A2(n_176), .B1(n_177), .B2(n_179), .C(n_182), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_641), .A2(n_190), .B1(n_191), .B2(n_194), .C(n_195), .Y(n_711) );
AO21x2_ASAP7_75t_L g712 ( .A1(n_595), .A2(n_223), .B(n_610), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_689), .Y(n_713) );
OAI211xp5_ASAP7_75t_L g714 ( .A1(n_635), .A2(n_644), .B(n_627), .C(n_649), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_640), .B(n_593), .Y(n_715) );
OAI221xp5_ASAP7_75t_SL g716 ( .A1(n_627), .A2(n_649), .B1(n_619), .B2(n_645), .C(n_630), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_608), .A2(n_624), .B1(n_661), .B2(n_660), .C(n_658), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_620), .A2(n_609), .B(n_599), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_625), .B(n_632), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_672), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_629), .A2(n_680), .B1(n_683), .B2(n_642), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_637), .B(n_636), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_682), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_678), .A2(n_598), .B(n_622), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_596), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_648), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_687), .B(n_616), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g728 ( .A1(n_674), .A2(n_631), .B(n_670), .C(n_638), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_601), .A2(n_589), .B(n_653), .Y(n_729) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_602), .B(n_590), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_687), .A2(n_638), .B1(n_631), .B2(n_670), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_656), .A2(n_662), .B1(n_603), .B2(n_623), .C(n_588), .Y(n_732) );
INVx2_ASAP7_75t_SL g733 ( .A(n_625), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_612), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_614), .B(n_615), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_653), .A2(n_614), .B(n_664), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_634), .A2(n_664), .B(n_643), .C(n_691), .Y(n_737) );
AOI21x1_ASAP7_75t_L g738 ( .A1(n_677), .A2(n_668), .B(n_665), .Y(n_738) );
AOI21xp33_ASAP7_75t_SL g739 ( .A1(n_647), .A2(n_657), .B(n_668), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_634), .A2(n_657), .B(n_665), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_690), .B(n_679), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_597), .A2(n_605), .B(n_606), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_647), .A2(n_690), .B1(n_591), .B2(n_616), .Y(n_743) );
AO21x2_ASAP7_75t_L g744 ( .A1(n_685), .A2(n_659), .B(n_675), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_616), .A2(n_591), .B1(n_667), .B2(n_646), .Y(n_745) );
INVx4_ASAP7_75t_L g746 ( .A(n_650), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_646), .A2(n_667), .B1(n_688), .B2(n_673), .Y(n_747) );
BUFx3_ASAP7_75t_L g748 ( .A(n_688), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_650), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_681), .A2(n_692), .B1(n_679), .B2(n_671), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_650), .A2(n_663), .B1(n_673), .B2(n_666), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_650), .B(n_663), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_663), .A2(n_673), .B1(n_618), .B2(n_611), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_613), .A2(n_617), .B1(n_633), .B2(n_669), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_618), .A2(n_577), .B1(n_501), .B2(n_470), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g756 ( .A1(n_639), .A2(n_450), .B(n_394), .C(n_522), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_600), .Y(n_757) );
BUFx3_ASAP7_75t_L g758 ( .A(n_689), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_607), .A2(n_604), .B(n_621), .Y(n_759) );
INVx3_ASAP7_75t_L g760 ( .A(n_689), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g761 ( .A1(n_654), .A2(n_544), .B(n_558), .Y(n_761) );
AO21x2_ASAP7_75t_L g762 ( .A1(n_739), .A2(n_740), .B(n_759), .Y(n_762) );
BUFx3_ASAP7_75t_L g763 ( .A(n_713), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_735), .Y(n_764) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_746), .Y(n_765) );
AND2x4_ASAP7_75t_SL g766 ( .A(n_713), .B(n_698), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_757), .B(n_756), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_734), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_697), .B(n_696), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_726), .B(n_720), .Y(n_770) );
INVx3_ASAP7_75t_L g771 ( .A(n_713), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_723), .B(n_708), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_699), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_708), .B(n_761), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_753), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_708), .B(n_701), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_699), .Y(n_777) );
INVxp67_ASAP7_75t_L g778 ( .A(n_715), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_717), .B(n_736), .Y(n_779) );
BUFx2_ASAP7_75t_L g780 ( .A(n_749), .Y(n_780) );
BUFx2_ASAP7_75t_L g781 ( .A(n_746), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_755), .B(n_758), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_709), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_725), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_733), .B(n_693), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_709), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_709), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_698), .B(n_760), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_709), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_741), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_722), .B(n_714), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_693), .B(n_721), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_719), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_729), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_729), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_719), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_703), .B(n_705), .Y(n_797) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_728), .B(n_702), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_744), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_716), .A2(n_714), .B1(n_700), .B2(n_732), .C(n_718), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_730), .B(n_727), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_727), .Y(n_802) );
OR2x6_ASAP7_75t_L g803 ( .A(n_727), .B(n_694), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_742), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_742), .Y(n_805) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_706), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_744), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_748), .B(n_745), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_738), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_752), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_712), .Y(n_811) );
INVx3_ASAP7_75t_SL g812 ( .A(n_747), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_712), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_737), .B(n_724), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_711), .Y(n_815) );
INVxp67_ASAP7_75t_L g816 ( .A(n_707), .Y(n_816) );
INVx5_ASAP7_75t_L g817 ( .A(n_731), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_750), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_750), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_710), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_695), .B(n_743), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_776), .B(n_751), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_785), .B(n_704), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_770), .Y(n_824) );
INVx4_ASAP7_75t_L g825 ( .A(n_781), .Y(n_825) );
AOI221xp5_ASAP7_75t_SL g826 ( .A1(n_791), .A2(n_754), .B1(n_767), .B2(n_800), .C(n_778), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_794), .Y(n_827) );
INVx2_ASAP7_75t_SL g828 ( .A(n_765), .Y(n_828) );
INVx4_ASAP7_75t_L g829 ( .A(n_781), .Y(n_829) );
INVx4_ASAP7_75t_L g830 ( .A(n_765), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_790), .B(n_774), .Y(n_831) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_765), .Y(n_832) );
INVx3_ASAP7_75t_L g833 ( .A(n_765), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_795), .Y(n_834) );
CKINVDCx16_ASAP7_75t_R g835 ( .A(n_784), .Y(n_835) );
NOR2xp33_ASAP7_75t_R g836 ( .A(n_763), .B(n_771), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_764), .B(n_779), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_768), .Y(n_838) );
INVx2_ASAP7_75t_SL g839 ( .A(n_765), .Y(n_839) );
AND2x2_ASAP7_75t_SL g840 ( .A(n_797), .B(n_772), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_795), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_792), .B(n_818), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_769), .B(n_810), .Y(n_843) );
NOR2x1_ASAP7_75t_SL g844 ( .A(n_803), .B(n_793), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_818), .B(n_819), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_806), .B(n_782), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_768), .B(n_780), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_793), .Y(n_848) );
AOI211xp5_ASAP7_75t_L g849 ( .A1(n_802), .A2(n_821), .B(n_812), .C(n_788), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_775), .A2(n_783), .B1(n_789), .B2(n_787), .C(n_786), .Y(n_850) );
OAI221xp5_ASAP7_75t_SL g851 ( .A1(n_803), .A2(n_821), .B1(n_816), .B2(n_775), .C(n_789), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_803), .A2(n_817), .B1(n_796), .B2(n_766), .Y(n_852) );
NAND2xp5_ASAP7_75t_SL g853 ( .A(n_798), .B(n_817), .Y(n_853) );
NOR2xp33_ASAP7_75t_R g854 ( .A(n_835), .B(n_796), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_840), .A2(n_815), .B1(n_820), .B2(n_817), .Y(n_855) );
BUFx2_ASAP7_75t_L g856 ( .A(n_825), .Y(n_856) );
INVx3_ASAP7_75t_L g857 ( .A(n_832), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_831), .B(n_804), .Y(n_858) );
NAND2x1p5_ASAP7_75t_L g859 ( .A(n_825), .B(n_817), .Y(n_859) );
NOR2xp33_ASAP7_75t_R g860 ( .A(n_829), .B(n_808), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_824), .B(n_801), .Y(n_861) );
CKINVDCx16_ASAP7_75t_R g862 ( .A(n_836), .Y(n_862) );
OR2x2_ASAP7_75t_L g863 ( .A(n_843), .B(n_805), .Y(n_863) );
BUFx2_ASAP7_75t_L g864 ( .A(n_829), .Y(n_864) );
NOR2x1p5_ASAP7_75t_L g865 ( .A(n_829), .B(n_773), .Y(n_865) );
INVx3_ASAP7_75t_L g866 ( .A(n_832), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_842), .B(n_762), .Y(n_867) );
INVx1_ASAP7_75t_SL g868 ( .A(n_836), .Y(n_868) );
AND3x2_ASAP7_75t_L g869 ( .A(n_849), .B(n_766), .C(n_814), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_837), .B(n_762), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g871 ( .A(n_826), .B(n_773), .C(n_777), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_823), .B(n_814), .Y(n_872) );
OAI33xp33_ASAP7_75t_L g873 ( .A1(n_846), .A2(n_811), .A3(n_813), .B1(n_809), .B2(n_799), .B3(n_807), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_827), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_830), .Y(n_875) );
OR2x2_ASAP7_75t_L g876 ( .A(n_845), .B(n_809), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_827), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_877), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_874), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_877), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_870), .B(n_834), .Y(n_881) );
BUFx2_ASAP7_75t_L g882 ( .A(n_860), .Y(n_882) );
INVx2_ASAP7_75t_SL g883 ( .A(n_865), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_862), .A2(n_851), .B1(n_852), .B2(n_848), .Y(n_884) );
NAND2x1_ASAP7_75t_L g885 ( .A(n_856), .B(n_830), .Y(n_885) );
AND2x4_ASAP7_75t_L g886 ( .A(n_872), .B(n_844), .Y(n_886) );
INVx4_ASAP7_75t_L g887 ( .A(n_862), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_867), .B(n_841), .Y(n_888) );
OAI21xp5_ASAP7_75t_SL g889 ( .A1(n_882), .A2(n_869), .B(n_868), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_887), .A2(n_868), .B1(n_864), .B2(n_855), .Y(n_890) );
XOR2x2_ASAP7_75t_SL g891 ( .A(n_884), .B(n_859), .Y(n_891) );
NAND2xp33_ASAP7_75t_SL g892 ( .A(n_887), .B(n_854), .Y(n_892) );
NAND3xp33_ASAP7_75t_SL g893 ( .A(n_885), .B(n_875), .C(n_859), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_878), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_883), .A2(n_858), .B1(n_863), .B2(n_861), .Y(n_895) );
INVxp67_ASAP7_75t_SL g896 ( .A(n_891), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_892), .A2(n_886), .B(n_853), .Y(n_897) );
XNOR2x1_ASAP7_75t_SL g898 ( .A(n_889), .B(n_828), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_896), .A2(n_895), .B1(n_890), .B2(n_893), .Y(n_899) );
OAI21xp5_ASAP7_75t_L g900 ( .A1(n_897), .A2(n_822), .B(n_871), .Y(n_900) );
OAI221xp5_ASAP7_75t_R g901 ( .A1(n_899), .A2(n_898), .B1(n_872), .B2(n_888), .C(n_881), .Y(n_901) );
AOI21xp5_ASAP7_75t_L g902 ( .A1(n_900), .A2(n_873), .B(n_894), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_902), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_903), .B(n_901), .Y(n_904) );
AND2x4_ASAP7_75t_L g905 ( .A(n_903), .B(n_879), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_905), .Y(n_906) );
XNOR2x1_ASAP7_75t_L g907 ( .A(n_904), .B(n_823), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_906), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_907), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_908), .B(n_905), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_909), .Y(n_911) );
OA21x2_ASAP7_75t_L g912 ( .A1(n_911), .A2(n_838), .B(n_828), .Y(n_912) );
AOI31xp33_ASAP7_75t_L g913 ( .A1(n_910), .A2(n_839), .A3(n_847), .B(n_876), .Y(n_913) );
NAND3xp33_ASAP7_75t_L g914 ( .A(n_912), .B(n_832), .C(n_850), .Y(n_914) );
AOI222xp33_ASAP7_75t_L g915 ( .A1(n_914), .A2(n_913), .B1(n_880), .B2(n_857), .C1(n_866), .C2(n_833), .Y(n_915) );
endmodule