module fake_jpeg_908_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_20),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_4),
.B(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_13),
.A2(n_11),
.B1(n_9),
.B2(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_7),
.B1(n_9),
.B2(n_14),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_18),
.A3(n_22),
.B1(n_14),
.B2(n_25),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_30),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_30),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

OAI322xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_28),
.A3(n_26),
.B1(n_21),
.B2(n_24),
.C1(n_16),
.C2(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_37),
.B1(n_41),
.B2(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_37),
.C(n_16),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_46),
.CI(n_24),
.CON(n_48),
.SN(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_46),
.C(n_39),
.Y(n_49)
);


endmodule