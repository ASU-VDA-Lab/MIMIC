module fake_jpeg_19811_n_214 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_47),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_2),
.B(n_3),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_22),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_29),
.B1(n_18),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_67),
.B1(n_71),
.B2(n_79),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_29),
.B1(n_31),
.B2(n_25),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_16),
.B(n_27),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_21),
.B1(n_18),
.B2(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_23),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_77),
.Y(n_102)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_38),
.A2(n_34),
.B1(n_24),
.B2(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_35),
.A2(n_30),
.B1(n_31),
.B2(n_15),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_22),
.B1(n_28),
.B2(n_6),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_94),
.B1(n_97),
.B2(n_103),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_26),
.B1(n_20),
.B2(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_23),
.B(n_15),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_65),
.B(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_4),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_106),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_58),
.B1(n_78),
.B2(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_66),
.Y(n_116)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_61),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_111),
.B(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_9),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_84),
.B1(n_90),
.B2(n_60),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_78),
.B(n_65),
.C(n_81),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_132),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_74),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_13),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_8),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_85),
.B1(n_83),
.B2(n_107),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_143),
.B1(n_149),
.B2(n_150),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_83),
.B1(n_85),
.B2(n_101),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_88),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_8),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_84),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_90),
.B1(n_60),
.B2(n_59),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_125),
.B1(n_133),
.B2(n_118),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_4),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_123),
.C(n_114),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_159),
.C(n_145),
.Y(n_171)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_112),
.C(n_117),
.D(n_120),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_152),
.B(n_137),
.C(n_142),
.D(n_144),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_129),
.B(n_127),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_169),
.B(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_153),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_175),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_169),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_144),
.C(n_138),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_182),
.C(n_164),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_180),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_135),
.C(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_191),
.C(n_182),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_150),
.B1(n_149),
.B2(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_158),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_190),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_161),
.B(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_157),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_176),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_198),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_179),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_188),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_175),
.C(n_139),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_161),
.B(n_146),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_199),
.B(n_202),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_184),
.B1(n_173),
.B2(n_183),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_194),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_118),
.C(n_109),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_109),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_211),
.Y(n_214)
);


endmodule