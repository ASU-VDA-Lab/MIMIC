module real_jpeg_22270_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_0),
.A2(n_21),
.B1(n_22),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_0),
.A2(n_36),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_0),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_2),
.A2(n_21),
.B(n_25),
.C(n_60),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_77),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_77),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_2),
.A2(n_10),
.B(n_49),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_2),
.B(n_93),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_50),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_23),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_4),
.Y(n_77)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_122),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_9),
.B(n_77),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_10),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_27),
.B(n_65),
.C(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_10),
.B(n_27),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_115),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_113),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_72),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_15),
.B(n_72),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_57),
.C(n_63),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_16),
.A2(n_17),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_18),
.B(n_39),
.C(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_24),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_20),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_24),
.B(n_25),
.C(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_42),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_22),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_26),
.A2(n_27),
.B(n_50),
.Y(n_60)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_28),
.A2(n_50),
.B(n_66),
.C(n_126),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_35),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_76),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_77),
.B(n_81),
.C(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_45),
.B(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_46),
.B(n_56),
.Y(n_153)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_52),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_48),
.B(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_50),
.B(n_89),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_50),
.B(n_62),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_51),
.B(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_59),
.A2(n_61),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_63),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_65),
.B(n_71),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_65),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_151),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_98),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_97),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_95),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_111),
.B2(n_112),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_110),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_101),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_172),
.B(n_178),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_155),
.B(n_171),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_142),
.B(n_154),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_131),
.B(n_141),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_123),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_136),
.B(n_140),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_157),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B1(n_162),
.B2(n_170),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_173),
.B(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);


endmodule