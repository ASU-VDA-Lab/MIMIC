module fake_jpeg_12840_n_196 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_33),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_0),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_68),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_107),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_79),
.B1(n_55),
.B2(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_78),
.B1(n_64),
.B2(n_65),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_59),
.C(n_66),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_83),
.B(n_81),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_67),
.B1(n_79),
.B2(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_101),
.B1(n_74),
.B2(n_72),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_72),
.B1(n_56),
.B2(n_80),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_116),
.B1(n_122),
.B2(n_125),
.Y(n_131)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_78),
.B1(n_64),
.B2(n_65),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_77),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_126),
.Y(n_140)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_71),
.B1(n_70),
.B2(n_69),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_83),
.B(n_62),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_127),
.Y(n_144)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_129),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_60),
.B1(n_57),
.B2(n_2),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_3),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_2),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_35),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_22),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_4),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_5),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_147),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_109),
.B(n_111),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_149),
.B(n_150),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_32),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_15),
.C(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_9),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_10),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_R g150 ( 
.A(n_118),
.B(n_13),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_14),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_15),
.B(n_16),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_168),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_23),
.Y(n_162)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_152),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_166),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_29),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_143),
.B1(n_149),
.B2(n_131),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_173),
.B1(n_159),
.B2(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_142),
.B1(n_42),
.B2(n_44),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_142),
.C(n_45),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_156),
.C(n_170),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_159),
.B1(n_155),
.B2(n_162),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_184),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_169),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_179),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_180),
.C(n_153),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_182),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_171),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_174),
.B(n_183),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_175),
.B(n_178),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_188),
.A3(n_164),
.B1(n_154),
.B2(n_49),
.C1(n_51),
.C2(n_40),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_176),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_46),
.Y(n_196)
);


endmodule