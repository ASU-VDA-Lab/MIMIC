module fake_jpeg_12516_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_48),
.Y(n_75)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_51),
.C(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_72),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_41),
.B1(n_49),
.B2(n_57),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_94),
.B1(n_40),
.B2(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_54),
.B(n_2),
.C(n_3),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_56),
.B(n_52),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_1),
.B(n_3),
.Y(n_103)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_95),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_44),
.B1(n_26),
.B2(n_28),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_1),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_103),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_23),
.C(n_39),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_105),
.C(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_104),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_4),
.B(n_5),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_29),
.C(n_37),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_24),
.C(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_31),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_14),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_6),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_114),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_119),
.B(n_108),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_104),
.B1(n_102),
.B2(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_122),
.B(n_124),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_118),
.B1(n_112),
.B2(n_109),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_126),
.C(n_125),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_32),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_34),
.C(n_38),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_115),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_117),
.Y(n_132)
);


endmodule