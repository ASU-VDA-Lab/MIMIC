module real_jpeg_32925_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_0),
.Y(n_115)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_0),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_45),
.B2(n_50),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_50),
.B1(n_104),
.B2(n_108),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_1),
.A2(n_50),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_45),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_2),
.A2(n_67),
.B1(n_258),
.B2(n_263),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_2),
.A2(n_67),
.B1(n_369),
.B2(n_372),
.Y(n_368)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_72),
.A3(n_78),
.B1(n_82),
.B2(n_90),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_3),
.A2(n_91),
.B1(n_202),
.B2(n_207),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_3),
.B(n_142),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_3),
.A2(n_100),
.B1(n_291),
.B2(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_3),
.B(n_347),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_3),
.A2(n_346),
.B(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_4),
.A2(n_282),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_4),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_5),
.Y(n_337)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_8),
.A2(n_121),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_9),
.A2(n_137),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_9),
.A2(n_137),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_9),
.A2(n_137),
.B1(n_391),
.B2(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_11),
.A2(n_152),
.B1(n_155),
.B2(n_158),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_11),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_11),
.A2(n_158),
.B1(n_242),
.B2(n_247),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_11),
.A2(n_158),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_11),
.A2(n_158),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_12),
.Y(n_331)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_14),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_14),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_176),
.B1(n_177),
.B2(n_181),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_15),
.A2(n_176),
.B1(n_217),
.B2(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_16),
.A2(n_263),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_16),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_409),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_321),
.B(n_408),
.Y(n_19)
);

OAI21x1_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_220),
.B(n_320),
.Y(n_20)
);

AOI211xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_128),
.B(n_195),
.C(n_196),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_22),
.A2(n_128),
.B(n_195),
.C(n_196),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_23),
.B(n_130),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_70),
.B1(n_126),
.B2(n_127),
.Y(n_23)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_24),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_24),
.B(n_126),
.C(n_129),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_40),
.B1(n_51),
.B2(n_65),
.Y(n_24)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_25),
.A2(n_240),
.B1(n_249),
.B2(n_250),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_25),
.B(n_91),
.Y(n_302)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_26),
.A2(n_66),
.B1(n_211),
.B2(n_219),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_27),
.A2(n_51),
.B1(n_212),
.B2(n_240),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_27),
.A2(n_40),
.B1(n_51),
.B2(n_399),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_27),
.A2(n_51),
.B1(n_399),
.B2(n_417),
.Y(n_416)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AO21x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_52),
.B(n_58),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_32),
.Y(n_180)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_37),
.Y(n_423)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_48),
.Y(n_218)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_49),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_49),
.Y(n_248)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_51),
.Y(n_219)
);

NAND2xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_58),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_61),
.Y(n_418)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_69),
.Y(n_401)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_97),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_71),
.A2(n_97),
.B1(n_98),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g159 ( 
.A1(n_82),
.A2(n_143),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_83),
.Y(n_440)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_84),
.Y(n_327)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_85),
.Y(n_344)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_91),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_91),
.B(n_235),
.Y(n_234)
);

OA21x2_ASAP7_75t_SL g250 ( 
.A1(n_91),
.A2(n_234),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_91),
.B(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_95),
.Y(n_238)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_112),
.B2(n_116),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_99),
.A2(n_116),
.B1(n_171),
.B2(n_175),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_99),
.A2(n_276),
.B1(n_283),
.B2(n_284),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_99),
.A2(n_175),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_100),
.A2(n_257),
.B1(n_264),
.B2(n_267),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_100),
.A2(n_277),
.B1(n_291),
.B2(n_298),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_100),
.A2(n_355),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_103),
.Y(n_267)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_107),
.Y(n_280)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_107),
.Y(n_359)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_110),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_115),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_115),
.Y(n_286)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_124),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_125),
.Y(n_297)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_168),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_131),
.B(n_169),
.C(n_185),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_141),
.B1(n_151),
.B2(n_159),
.Y(n_131)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_132),
.Y(n_365)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_141),
.A2(n_151),
.B1(n_159),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_141),
.A2(n_159),
.B1(n_368),
.B2(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_142),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g366 ( 
.A(n_159),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_184),
.B2(n_185),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_173),
.Y(n_309)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_174),
.Y(n_301)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_186),
.A2(n_377),
.B1(n_382),
.B2(n_390),
.Y(n_376)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_186),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_187),
.B(n_384),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_210),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_197),
.B(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_199),
.A2(n_200),
.B1(n_210),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_209),
.Y(n_371)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_209),
.Y(n_374)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_219),
.Y(n_249)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_314),
.B(n_319),
.Y(n_220)
);

OAI21x1_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_273),
.B(n_313),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_255),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_223),
.B(n_255),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_239),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_224),
.B(n_239),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_227),
.B(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B(n_234),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx4f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_248),
.Y(n_404)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_268),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_270),
.C(n_271),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_288),
.B(n_312),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_287),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_287),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_303),
.B(n_311),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_302),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_302),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_407),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_322),
.B(n_407),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_363),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_362),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_324),
.B(n_363),
.C(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_350),
.B1(n_360),
.B2(n_361),
.Y(n_324)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

OAI32xp33_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_328),
.A3(n_332),
.B1(n_338),
.B2(n_345),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g447 ( 
.A1(n_326),
.A2(n_328),
.A3(n_332),
.B1(n_338),
.B2(n_345),
.Y(n_447)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_351),
.Y(n_420)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_361),
.B(n_447),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_375),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_364),
.B(n_405),
.C(n_406),
.Y(n_424)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_398),
.B1(n_405),
.B2(n_406),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_385),
.B1(n_387),
.B2(n_389),
.Y(n_384)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_383),
.A2(n_429),
.B1(n_430),
.B2(n_436),
.Y(n_428)
);

INVx3_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_390),
.Y(n_436)
);

INVx8_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_398),
.Y(n_406)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_448),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_411),
.B(n_413),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_425),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_424),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_446),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_437),
.B2(n_438),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);


endmodule