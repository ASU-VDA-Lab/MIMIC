module real_jpeg_8709_n_17 (n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_1),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_69),
.B1(n_72),
.B2(n_84),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_84),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_84),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_3),
.B(n_35),
.Y(n_201)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_47),
.B(n_64),
.C(n_102),
.D(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_45),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_3),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_123),
.B(n_125),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_3),
.A2(n_34),
.B(n_41),
.C(n_159),
.D(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_34),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_38),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_140),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_143),
.B(n_169),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_9),
.A2(n_37),
.B1(n_69),
.B2(n_72),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_9),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_28),
.B1(n_69),
.B2(n_72),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_10),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_11),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_11),
.A2(n_69),
.B1(n_72),
.B2(n_117),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_117),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_117),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_12),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_69),
.B1(n_72),
.B2(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_105),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_105),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_14),
.A2(n_61),
.B1(n_69),
.B2(n_72),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_15),
.A2(n_69),
.B1(n_72),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_15),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_122),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_122),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_16),
.A2(n_50),
.B1(n_69),
.B2(n_72),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_51),
.B1(n_52),
.B2(n_75),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_31),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_27),
.A2(n_31),
.B(n_140),
.C(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_29),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_29),
.B(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_30),
.A2(n_33),
.B1(n_60),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_30),
.A2(n_33),
.B1(n_234),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_30),
.A2(n_219),
.B(n_257),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_33),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_33),
.A2(n_83),
.B(n_235),
.Y(n_298)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_38),
.B(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_48),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_41),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_41),
.A2(n_45),
.B1(n_254),
.B2(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_41),
.A2(n_45),
.B1(n_89),
.B2(n_272),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_43),
.B(n_46),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_65),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_47),
.A2(n_159),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.C(n_62),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_55),
.A2(n_57),
.B1(n_179),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_55),
.A2(n_214),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_57),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_57),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_57),
.A2(n_180),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_59),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_62),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_73),
.B(n_74),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_73),
.B1(n_116),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_63),
.A2(n_157),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_63),
.A2(n_73),
.B1(n_211),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_63),
.A2(n_73),
.B1(n_229),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_63),
.A2(n_73),
.B1(n_248),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_64),
.A2(n_68),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_72),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_69),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_72),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_73),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_73),
.A2(n_118),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_74),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.C(n_85),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_317),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_82),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_82),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_85),
.B(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_314),
.A3(n_324),
.B1(n_329),
.B2(n_330),
.C(n_332),
.Y(n_92)
);

AOI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_264),
.A3(n_302),
.B1(n_308),
.B2(n_313),
.C(n_333),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_222),
.C(n_261),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_194),
.B(n_221),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_173),
.B(n_193),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_151),
.B(n_172),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_128),
.B(n_150),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_100),
.B(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B(n_125),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_127),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_123),
.A2(n_124),
.B1(n_170),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_123),
.A2(n_124),
.B1(n_184),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_123),
.A2(n_124),
.B1(n_204),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_123),
.A2(n_124),
.B1(n_227),
.B2(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_123),
.A2(n_124),
.B(n_246),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_132),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_137),
.B(n_149),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_144),
.B(n_148),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_141),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_164),
.B2(n_171),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_163),
.C(n_171),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_175),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_189),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_190),
.C(n_191),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_182),
.B2(n_188),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_185),
.C(n_186),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_196),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_198),
.B(n_207),
.C(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_203),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_223),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_241),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_224),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_224),
.B(n_241),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_230),
.CI(n_231),
.CON(n_224),
.SN(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_240),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_259),
.B2(n_260),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_249),
.C(n_260),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_255),
.C(n_258),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_282),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_265),
.B(n_282),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.C(n_281),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_271),
.C(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_277),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_294),
.B(n_298),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_278),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_300),
.B2(n_301),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_292),
.B2(n_293),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_293),
.C(n_301),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_290),
.B(n_291),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_290),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_291),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_291),
.A2(n_316),
.B1(n_320),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_299),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_296),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_309),
.B(n_312),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_322),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_322),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.C(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);


endmodule