module fake_aes_12431_n_726 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_726);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_726;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_86), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_42), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_19), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_21), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_60), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_87), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_66), .B(n_82), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_51), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_65), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_28), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_56), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_18), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_26), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_14), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_62), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_72), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_13), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_76), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
BUFx2_ASAP7_75t_SL g119 ( .A(n_68), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_77), .B(n_55), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_9), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_38), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_0), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_5), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_70), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_1), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_69), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_96), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_109), .B(n_0), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_95), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_107), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_110), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_98), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_98), .Y(n_139) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_91), .A2(n_50), .B(n_89), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_130), .Y(n_141) );
INVx5_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_130), .B(n_6), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_94), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_101), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_110), .B(n_7), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_146), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVxp67_ASAP7_75t_SL g153 ( .A(n_131), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_142), .B(n_108), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_142), .B(n_118), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
AND3x2_ASAP7_75t_L g161 ( .A(n_133), .B(n_113), .C(n_128), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_131), .A2(n_93), .B1(n_123), .B2(n_100), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_142), .B(n_105), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_142), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_137), .A2(n_129), .B1(n_116), .B2(n_92), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_141), .A2(n_125), .B1(n_115), .B2(n_119), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_144), .B(n_148), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_142), .B(n_105), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVxp67_ASAP7_75t_SL g175 ( .A(n_141), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVxp33_ASAP7_75t_SL g179 ( .A(n_150), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_153), .B(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_153), .B(n_149), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_175), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_175), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_179), .B(n_133), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_163), .B(n_133), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_157), .B(n_149), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_163), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_163), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_169), .A2(n_137), .B1(n_148), .B2(n_144), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
BUFx5_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
NOR2x1p5_ASAP7_75t_L g194 ( .A(n_170), .B(n_116), .Y(n_194) );
NAND2xp33_ASAP7_75t_L g195 ( .A(n_169), .B(n_111), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_169), .A2(n_104), .B1(n_129), .B2(n_147), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_157), .B(n_145), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_156), .Y(n_199) );
NOR3xp33_ASAP7_75t_L g200 ( .A(n_170), .B(n_136), .C(n_135), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_169), .A2(n_147), .B1(n_145), .B2(n_139), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_139), .B(n_138), .C(n_121), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_163), .B(n_111), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_163), .B(n_114), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_168), .B(n_114), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_167), .B(n_117), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_168), .B(n_117), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_168), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_167), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_168), .B(n_120), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_168), .B(n_103), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_172), .B(n_120), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_161), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_172), .B(n_124), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_161), .B(n_124), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_186), .A2(n_159), .B(n_162), .Y(n_221) );
OA22x2_ASAP7_75t_L g222 ( .A1(n_191), .A2(n_135), .B1(n_162), .B2(n_174), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_187), .A2(n_160), .B(n_159), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_183), .A2(n_171), .B1(n_164), .B2(n_158), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_219), .B(n_164), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_193), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_183), .A2(n_171), .B1(n_158), .B2(n_160), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_184), .A2(n_159), .B1(n_160), .B2(n_162), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_184), .B(n_176), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_202), .A2(n_174), .B(n_166), .C(n_173), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
CKINVDCx8_ASAP7_75t_R g234 ( .A(n_213), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_219), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_182), .B(n_176), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_215), .B(n_176), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_219), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_193), .Y(n_239) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_198), .A2(n_174), .B(n_155), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_181), .A2(n_178), .B(n_177), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_193), .B(n_176), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_191), .A2(n_180), .B1(n_178), .B2(n_177), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_189), .A2(n_180), .B(n_178), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_193), .B(n_185), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
OAI21xp33_ASAP7_75t_L g247 ( .A1(n_214), .A2(n_126), .B(n_177), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_201), .A2(n_180), .B1(n_176), .B2(n_127), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_204), .A2(n_119), .B1(n_122), .B2(n_152), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_215), .B(n_8), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_194), .B(n_8), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_194), .B(n_9), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_200), .A2(n_154), .B1(n_152), .B2(n_102), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_251), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_234), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_247), .A2(n_195), .B(n_205), .C(n_212), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_251), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_244), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_226), .B(n_193), .Y(n_259) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_217), .A3(n_199), .B(n_209), .Y(n_260) );
BUFx2_ASAP7_75t_SL g261 ( .A(n_246), .Y(n_261) );
AO31x2_ASAP7_75t_L g262 ( .A1(n_228), .A2(n_217), .A3(n_199), .B(n_209), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_221), .A2(n_188), .B(n_190), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_240), .A2(n_192), .B(n_208), .Y(n_264) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_223), .A2(n_217), .B(n_199), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_203), .B(n_207), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_190), .B(n_188), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_233), .A2(n_220), .B(n_216), .C(n_206), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_230), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_226), .A2(n_218), .B1(n_211), .B2(n_210), .Y(n_272) );
AOI221x1_ASAP7_75t_L g273 ( .A1(n_249), .A2(n_152), .B1(n_154), .B2(n_209), .C(n_208), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_238), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_246), .B(n_210), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_224), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_258), .A2(n_235), .B(n_227), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_259), .A2(n_240), .B(n_243), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_258), .A2(n_235), .B(n_227), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_268), .A2(n_234), .B1(n_222), .B2(n_252), .C(n_253), .Y(n_280) );
BUFx12f_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_264), .A2(n_244), .B(n_248), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_269), .B(n_222), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_256), .A2(n_250), .B(n_252), .C(n_245), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_266), .A2(n_224), .B(n_239), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_273), .A2(n_243), .B(n_242), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_267), .A2(n_239), .B(n_232), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_264), .A2(n_232), .B(n_236), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_271), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_274), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_269), .B(n_222), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_225), .B(n_218), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
BUFx8_ASAP7_75t_SL g296 ( .A(n_255), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_273), .A2(n_192), .B(n_208), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_265), .A2(n_189), .B(n_192), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_257), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_282), .B(n_260), .Y(n_300) );
INVx8_ASAP7_75t_L g301 ( .A(n_281), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_282), .B(n_260), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_290), .B(n_291), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_278), .B(n_260), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_290), .B(n_260), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_297), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_285), .A2(n_263), .B(n_265), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_297), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_294), .A2(n_265), .B(n_275), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_283), .A2(n_262), .B(n_260), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_278), .A2(n_262), .B(n_275), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_295), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_280), .B(n_254), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_297), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_283), .B(n_261), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_298), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_297), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_262), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_292), .B(n_262), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_289), .A2(n_262), .B(n_275), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_292), .A2(n_257), .B1(n_261), .B2(n_237), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_287), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_284), .B(n_265), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_287), .Y(n_329) );
OA21x2_ASAP7_75t_L g330 ( .A1(n_277), .A2(n_237), .B(n_189), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_287), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_324), .B(n_299), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_301), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_306), .Y(n_334) );
INVxp67_ASAP7_75t_SL g335 ( .A(n_323), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_324), .Y(n_336) );
BUFx12f_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_328), .B(n_279), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_319), .B(n_276), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_319), .B(n_276), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_328), .B(n_286), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_319), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_320), .B(n_288), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_306), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_320), .B(n_300), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_306), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_320), .B(n_276), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_306), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_313), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_300), .B(n_10), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_302), .B(n_276), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_303), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_330), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_322), .B(n_281), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_301), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_305), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_308), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_305), .B(n_276), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_305), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_303), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_301), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_326), .B(n_10), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_310), .Y(n_374) );
INVx5_ASAP7_75t_L g375 ( .A(n_316), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_308), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_316), .B(n_270), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_301), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_326), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_321), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_321), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_310), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_329), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_355), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_342), .B(n_329), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_354), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_373), .B(n_304), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_332), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_336), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_373), .B(n_304), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_333), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_346), .B(n_304), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_337), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_342), .B(n_331), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_346), .B(n_304), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_332), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_352), .B(n_312), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_337), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_352), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_351), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_362), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_334), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_362), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_371), .B(n_312), .Y(n_408) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_359), .B(n_310), .Y(n_409) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_372), .B(n_322), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_358), .B(n_331), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_343), .Y(n_412) );
NOR2xp33_ASAP7_75t_SL g413 ( .A(n_372), .B(n_301), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_358), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_375), .B(n_316), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_360), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_360), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_363), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_363), .B(n_304), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_368), .B(n_304), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_334), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_380), .B(n_339), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_375), .B(n_316), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_380), .B(n_327), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_386), .B(n_327), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_350), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_337), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_381), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_339), .B(n_312), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_340), .B(n_312), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_344), .B(n_325), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_379), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_340), .B(n_325), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_348), .B(n_314), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_338), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_348), .B(n_325), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_338), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_366), .B(n_314), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_366), .B(n_325), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_375), .B(n_310), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_353), .B(n_311), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_353), .B(n_309), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_341), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_341), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_345), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_379), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_345), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_375), .B(n_316), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_353), .B(n_309), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_353), .B(n_311), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_344), .B(n_311), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_345), .B(n_311), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_347), .B(n_311), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_382), .B(n_317), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_382), .B(n_317), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_347), .B(n_311), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_347), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_383), .B(n_315), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_383), .B(n_317), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_349), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_377), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_349), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_463), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_392), .B(n_385), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_432), .B(n_385), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_396), .B(n_369), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_402), .B(n_375), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_399), .B(n_364), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_463), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_393), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_437), .B(n_364), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_400), .B(n_369), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_415), .B(n_375), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_389), .B(n_349), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_402), .B(n_361), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_435), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_419), .B(n_361), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_465), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_441), .B(n_377), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_390), .B(n_356), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_393), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_442), .B(n_361), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_391), .B(n_361), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_394), .B(n_356), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_403), .B(n_356), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_423), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_465), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_404), .B(n_357), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_420), .B(n_357), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_406), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_424), .B(n_357), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_414), .B(n_365), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_416), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_413), .A2(n_301), .B1(n_377), .B2(n_375), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_417), .B(n_365), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_418), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_422), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_438), .B(n_365), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_387), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_445), .B(n_377), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_426), .B(n_367), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_412), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_452), .B(n_377), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_412), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_440), .B(n_376), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_420), .B(n_376), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_446), .B(n_376), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_429), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_378), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_429), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_388), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_388), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_406), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_398), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_458), .B(n_378), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_436), .B(n_378), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_398), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_411), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_435), .B(n_367), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_421), .Y(n_524) );
AND2x2_ASAP7_75t_SL g525 ( .A(n_426), .B(n_367), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_411), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_397), .B(n_367), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_421), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_405), .B(n_407), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_449), .B(n_384), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_451), .Y(n_531) );
NAND2x1_ASAP7_75t_L g532 ( .A(n_409), .B(n_384), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_410), .A2(n_301), .B1(n_374), .B2(n_384), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_428), .Y(n_534) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_387), .A2(n_374), .B(n_384), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_439), .B(n_317), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_451), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_428), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_430), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_433), .B(n_335), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_447), .B(n_317), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_462), .B(n_335), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_443), .B(n_323), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_427), .B(n_315), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_444), .B(n_315), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_401), .B(n_323), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_425), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_425), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_434), .B(n_323), .Y(n_549) );
OAI21xp33_ASAP7_75t_L g550 ( .A1(n_454), .A2(n_307), .B(n_318), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_410), .A2(n_330), .B1(n_318), .B2(n_307), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_453), .B(n_318), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_434), .B(n_318), .Y(n_553) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_455), .B(n_330), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_464), .B(n_408), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g557 ( .A1(n_503), .A2(n_431), .B1(n_454), .B2(n_461), .C1(n_395), .C2(n_448), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_469), .B(n_431), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_480), .A2(n_461), .B1(n_460), .B2(n_450), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_495), .B(n_456), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_480), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_534), .B(n_459), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_494), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_469), .A2(n_551), .B1(n_512), .B2(n_514), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_468), .B(n_450), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_506), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_517), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_539), .B(n_11), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_529), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_508), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_497), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_539), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_468), .B(n_330), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_500), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_503), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_538), .B(n_330), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_520), .B(n_330), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_515), .B(n_12), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_498), .A2(n_237), .B1(n_296), .B2(n_15), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_475), .B(n_12), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_517), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_488), .B(n_13), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_516), .B(n_15), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_518), .B(n_521), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_522), .B(n_16), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_501), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_488), .B(n_16), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_524), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_490), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_526), .B(n_17), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_528), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_466), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_493), .B(n_17), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_487), .B(n_483), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_476), .B(n_18), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_493), .B(n_154), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_533), .A2(n_154), .B1(n_152), .B2(n_193), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_154), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_554), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_510), .B(n_152), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_471), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_478), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_467), .B(n_20), .Y(n_606) );
CKINVDCx14_ASAP7_75t_R g607 ( .A(n_486), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_528), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_487), .B(n_22), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_486), .B(n_23), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_484), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_471), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_472), .B(n_24), .Y(n_613) );
INVxp67_ASAP7_75t_SL g614 ( .A(n_466), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_481), .B(n_25), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_545), .B(n_552), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_477), .B(n_27), .Y(n_617) );
NOR2xp67_ASAP7_75t_L g618 ( .A(n_470), .B(n_30), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_545), .B(n_31), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_481), .B(n_32), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_489), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_502), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_552), .B(n_513), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_555), .A2(n_196), .B1(n_218), .B2(n_211), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_477), .B(n_33), .Y(n_625) );
AND2x2_ASAP7_75t_SL g626 ( .A(n_525), .B(n_34), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_504), .B(n_35), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_560), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_565), .A2(n_507), .B(n_525), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_607), .B(n_470), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_622), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_605), .Y(n_632) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_598), .A2(n_532), .B(n_523), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_557), .B(n_513), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_565), .A2(n_550), .B1(n_531), .B2(n_470), .C(n_537), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_607), .A2(n_531), .B1(n_537), .B2(n_479), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_611), .B(n_519), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_621), .B(n_519), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_558), .B(n_541), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_604), .A2(n_612), .B1(n_561), .B2(n_602), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_616), .B(n_546), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_574), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_581), .A2(n_537), .B1(n_531), .B2(n_477), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_593), .A2(n_542), .B1(n_536), .B2(n_553), .C1(n_544), .C2(n_511), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_573), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_602), .B(n_505), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_576), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_589), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_556), .B(n_473), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_571), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_623), .B(n_549), .Y(n_651) );
OAI322xp33_ASAP7_75t_L g652 ( .A1(n_598), .A2(n_509), .A3(n_492), .B1(n_496), .B2(n_499), .C1(n_523), .C2(n_482), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_626), .A2(n_527), .B1(n_505), .B2(n_535), .Y(n_653) );
AO221x1_ASAP7_75t_L g654 ( .A1(n_626), .A2(n_473), .B1(n_482), .B2(n_491), .C(n_548), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_590), .A2(n_505), .B1(n_491), .B2(n_543), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_564), .B(n_548), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_592), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_577), .A2(n_543), .B1(n_530), .B2(n_547), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_568), .B(n_547), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_572), .B(n_37), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_562), .B(n_39), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_587), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_577), .A2(n_211), .B1(n_43), .B2(n_45), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_597), .B(n_40), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_575), .B(n_48), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_559), .A2(n_49), .B1(n_52), .B2(n_53), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_593), .A2(n_54), .B(n_57), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_570), .A2(n_196), .B1(n_61), .B2(n_63), .C1(n_64), .C2(n_67), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_567), .B(n_90), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_595), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_640), .A2(n_570), .B(n_584), .C(n_596), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_631), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_641), .B(n_579), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_629), .A2(n_618), .B(n_582), .C(n_617), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_654), .A2(n_627), .B1(n_609), .B2(n_620), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_642), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g677 ( .A1(n_643), .A2(n_580), .B1(n_586), .B2(n_588), .C(n_619), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_668), .A2(n_601), .B(n_603), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_636), .A2(n_625), .B(n_617), .C(n_610), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_630), .B(n_595), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_634), .A2(n_615), .B1(n_613), .B2(n_599), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_632), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_628), .B(n_614), .Y(n_683) );
AOI221xp5_ASAP7_75t_SL g684 ( .A1(n_652), .A2(n_614), .B1(n_578), .B2(n_606), .C(n_563), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_670), .Y(n_685) );
OAI322xp33_ASAP7_75t_L g686 ( .A1(n_662), .A2(n_591), .A3(n_566), .B1(n_569), .B2(n_608), .C1(n_583), .C2(n_594), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_653), .B(n_625), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_637), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_652), .A2(n_591), .B1(n_566), .B2(n_569), .C(n_608), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_658), .A2(n_594), .B1(n_583), .B2(n_585), .C(n_563), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_633), .A2(n_635), .B(n_655), .C(n_642), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_644), .A2(n_625), .B1(n_617), .B2(n_585), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_650), .A2(n_600), .B1(n_624), .B2(n_73), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_661), .A2(n_58), .B(n_71), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_646), .A2(n_74), .B1(n_75), .B2(n_78), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_638), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_665), .A2(n_79), .B(n_80), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_646), .A2(n_667), .B(n_664), .C(n_666), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_663), .B(n_83), .C(n_84), .Y(n_699) );
O2A1O1Ixp5_ASAP7_75t_L g700 ( .A1(n_645), .A2(n_88), .B(n_647), .C(n_648), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_657), .B(n_639), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_649), .A2(n_669), .B(n_656), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_659), .Y(n_703) );
AOI21xp33_ASAP7_75t_SL g704 ( .A1(n_651), .A2(n_640), .B(n_636), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_704), .B(n_700), .C(n_687), .Y(n_705) );
OAI221xp5_ASAP7_75t_SL g706 ( .A1(n_691), .A2(n_674), .B1(n_675), .B2(n_692), .C(n_679), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_693), .B(n_678), .C(n_684), .Y(n_707) );
NOR2xp67_ASAP7_75t_L g708 ( .A(n_676), .B(n_685), .Y(n_708) );
NAND4xp75_ASAP7_75t_L g709 ( .A(n_678), .B(n_694), .C(n_690), .D(n_681), .Y(n_709) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_671), .B(n_698), .C(n_699), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_709), .B(n_672), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
NOR3xp33_ASAP7_75t_SL g713 ( .A(n_706), .B(n_677), .C(n_695), .Y(n_713) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_708), .B(n_686), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_712), .A2(n_707), .B1(n_705), .B2(n_682), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_711), .B(n_694), .C(n_697), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_714), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_716), .B(n_713), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_717), .Y(n_719) );
AOI22x1_ASAP7_75t_L g720 ( .A1(n_718), .A2(n_715), .B1(n_703), .B2(n_696), .Y(n_720) );
AOI22x1_ASAP7_75t_L g721 ( .A1(n_718), .A2(n_688), .B1(n_680), .B2(n_683), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_721), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_722), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_719), .B(n_720), .Y(n_724) );
AO21x1_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_701), .B(n_660), .Y(n_725) );
AOI211xp5_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_702), .B(n_689), .C(n_673), .Y(n_726) );
endmodule