module fake_jpeg_19523_n_70 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_56;
wire n_31;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_13),
.B1(n_25),
.B2(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_30),
.B1(n_35),
.B2(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_2),
.B1(n_5),
.B2(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_1),
.Y(n_54)
);

AO21x1_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_57),
.B(n_58),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_34),
.B(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_47),
.B1(n_46),
.B2(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_2),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_9),
.B(n_10),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_11),
.C(n_12),
.Y(n_64)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_55),
.C(n_17),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_16),
.B(n_22),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_63),
.C(n_27),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_62),
.B(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_23),
.Y(n_70)
);


endmodule