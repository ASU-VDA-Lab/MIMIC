module fake_jpeg_4935_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_25),
.B1(n_27),
.B2(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_30),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_20),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_31),
.B1(n_28),
.B2(n_26),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_51),
.B1(n_54),
.B2(n_64),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_53),
.B1(n_29),
.B2(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_35),
.A2(n_21),
.B1(n_19),
.B2(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_58),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_36),
.B1(n_39),
.B2(n_33),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_76),
.B1(n_79),
.B2(n_65),
.Y(n_89)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_75),
.B1(n_72),
.B2(n_68),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_38),
.B(n_37),
.C(n_40),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_45),
.B1(n_46),
.B2(n_62),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_40),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_59),
.B1(n_53),
.B2(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_101),
.B1(n_74),
.B2(n_75),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_72),
.B1(n_81),
.B2(n_78),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_99),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_51),
.B1(n_64),
.B2(n_43),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_103),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_62),
.B1(n_54),
.B2(n_63),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_80),
.B(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_50),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_52),
.B1(n_50),
.B2(n_60),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_79),
.B1(n_83),
.B2(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_40),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_114),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_124),
.B1(n_128),
.B2(n_57),
.Y(n_159)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_75),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_126),
.B(n_134),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_97),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_96),
.B1(n_94),
.B2(n_101),
.Y(n_139)
);

HAxp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_62),
.CON(n_126),
.SN(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_77),
.B1(n_81),
.B2(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_73),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_94),
.B(n_110),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_129),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_150),
.C(n_151),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_142),
.B(n_148),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_141),
.B1(n_145),
.B2(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_143),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_99),
.B1(n_77),
.B2(n_69),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_68),
.B1(n_37),
.B2(n_38),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_20),
.B(n_23),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_40),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_58),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_98),
.C(n_104),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_13),
.C(n_14),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_159),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_37),
.B1(n_38),
.B2(n_98),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_131),
.B(n_133),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_116),
.C(n_111),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_114),
.B1(n_113),
.B2(n_117),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_166),
.B(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_168),
.Y(n_195)
);

OR2x6_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_118),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_177),
.C(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_174),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_183),
.B1(n_142),
.B2(n_138),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_136),
.B1(n_143),
.B2(n_145),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_188),
.B1(n_196),
.B2(n_162),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_193),
.B(n_198),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_163),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_135),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_204),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_123),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_122),
.B1(n_93),
.B2(n_88),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_182),
.B(n_183),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_122),
.C(n_93),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.C(n_194),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_93),
.B1(n_88),
.B2(n_97),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_88),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_165),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_216),
.C(n_217),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_213),
.B1(n_219),
.B2(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_164),
.B1(n_178),
.B2(n_171),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_177),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_191),
.C(n_203),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_169),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_171),
.B1(n_11),
.B2(n_12),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_97),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_19),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_219),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_193),
.B1(n_196),
.B2(n_187),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_195),
.C(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_229),
.C(n_1),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_192),
.C(n_61),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_30),
.B1(n_22),
.B2(n_57),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_10),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_0),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_57),
.B1(n_61),
.B2(n_2),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_210),
.B1(n_61),
.B2(n_213),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_0),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_9),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_237),
.B(n_234),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_7),
.B(n_14),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_211),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_243),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_241),
.B(n_246),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_10),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_247),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_61),
.C(n_2),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_6),
.B(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_249),
.B(n_12),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_231),
.B(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_258),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_235),
.B1(n_232),
.B2(n_226),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_1),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_247),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_226),
.B1(n_225),
.B2(n_11),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_241),
.C(n_6),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_225),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_257),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_265),
.B(n_5),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_5),
.C(n_11),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_263),
.C(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_5),
.C(n_12),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_268),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_266),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_270),
.B(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_256),
.C(n_250),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_265),
.C(n_14),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_3),
.B(n_4),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_3),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_274),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_3),
.Y(n_279)
);


endmodule