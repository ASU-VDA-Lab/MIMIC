module fake_jpeg_24673_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_288;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_7),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_40),
.C(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_34),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_48),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_34),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_19),
.B(n_22),
.C(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_36),
.B1(n_28),
.B2(n_17),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_37),
.B1(n_28),
.B2(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_72),
.A2(n_86),
.B1(n_87),
.B2(n_27),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_36),
.B1(n_17),
.B2(n_34),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_82),
.B1(n_98),
.B2(n_23),
.Y(n_108)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_96),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_30),
.B1(n_37),
.B2(n_32),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_80),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_22),
.B(n_20),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_39),
.B1(n_45),
.B2(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_35),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_41),
.B1(n_32),
.B2(n_21),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_26),
.B1(n_31),
.B2(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_41),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_107),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_47),
.B(n_44),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_63),
.B(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_54),
.B1(n_44),
.B2(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_55),
.B(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_56),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_0),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_108),
.A2(n_101),
.B1(n_77),
.B2(n_104),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_23),
.B1(n_33),
.B2(n_58),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_121),
.B1(n_127),
.B2(n_78),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_0),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_133),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_136),
.B(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_63),
.B1(n_61),
.B2(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_73),
.B1(n_96),
.B2(n_92),
.Y(n_148)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_33),
.B1(n_35),
.B2(n_27),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_35),
.B1(n_27),
.B2(n_22),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_35),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_22),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_133),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_1),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_97),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_149),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_73),
.B1(n_95),
.B2(n_106),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_157),
.B1(n_135),
.B2(n_125),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_148),
.B1(n_155),
.B2(n_163),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_95),
.B(n_107),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_70),
.B(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_107),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_126),
.C(n_109),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_133),
.B(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_128),
.B1(n_116),
.B2(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_84),
.B1(n_93),
.B2(n_74),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_97),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_88),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_162),
.Y(n_186)
);

OAI22x1_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_19),
.B1(n_20),
.B2(n_85),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_125),
.B1(n_91),
.B2(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_117),
.B(n_88),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_103),
.B1(n_105),
.B2(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_79),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_133),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_132),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_189),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_132),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_194),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_190),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_176),
.B(n_178),
.Y(n_202)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_129),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_115),
.B1(n_110),
.B2(n_123),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_166),
.B1(n_153),
.B2(n_144),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_121),
.B1(n_110),
.B2(n_135),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_183),
.B1(n_195),
.B2(n_142),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_158),
.C(n_156),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_165),
.B1(n_154),
.B2(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_20),
.B1(n_19),
.B2(n_85),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_218),
.B1(n_220),
.B2(n_195),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_141),
.B1(n_167),
.B2(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_184),
.C(n_176),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_208),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_155),
.B1(n_163),
.B2(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_168),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_216),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_164),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_164),
.B1(n_68),
.B2(n_19),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_68),
.B1(n_2),
.B2(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_2),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_219),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_225),
.Y(n_246)
);

OAI21x1_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_178),
.B(n_181),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_230),
.B1(n_232),
.B2(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_236),
.C(n_237),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_171),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_183),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_239),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_211),
.B(n_205),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_188),
.C(n_193),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_188),
.C(n_191),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_190),
.B(n_173),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_201),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_186),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_243),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_252),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_224),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_215),
.B1(n_214),
.B2(n_204),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_235),
.B1(n_223),
.B2(n_195),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_182),
.B1(n_210),
.B2(n_208),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_253),
.B1(n_228),
.B2(n_219),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_196),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_218),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_213),
.C(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_237),
.C(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_230),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_255),
.C(n_247),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_3),
.B(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_221),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

AO221x1_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_174),
.B1(n_200),
.B2(n_216),
.C(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_274),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_5),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_275),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_283),
.A3(n_174),
.B1(n_257),
.B2(n_273),
.C1(n_263),
.C2(n_276),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_261),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_284),
.B(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_286),
.C(n_288),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_262),
.A3(n_259),
.B1(n_260),
.B2(n_265),
.C1(n_13),
.C2(n_6),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_289),
.B(n_6),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_15),
.B1(n_9),
.B2(n_11),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_15),
.B(n_9),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_282),
.B(n_12),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_11),
.C(n_13),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_11),
.B(n_13),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_293),
.B(n_14),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_14),
.Y(n_298)
);


endmodule