module fake_jpeg_650_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_10),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_51),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_67),
.B1(n_64),
.B2(n_53),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_54),
.B1(n_50),
.B2(n_53),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_64),
.B1(n_70),
.B2(n_66),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_57),
.B1(n_55),
.B2(n_54),
.Y(n_97)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_65),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_58),
.Y(n_96)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_97),
.B1(n_82),
.B2(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_75),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_52),
.B1(n_56),
.B2(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_59),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_76),
.Y(n_106)
);

NOR2x1_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_112),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_55),
.B(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_111),
.B(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_119),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_116),
.B1(n_16),
.B2(n_43),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_84),
.B1(n_58),
.B2(n_17),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_132),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_87),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_127),
.B(n_7),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_84),
.B1(n_58),
.B2(n_4),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_8),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_2),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_44),
.B(n_41),
.C(n_34),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_29),
.B(n_25),
.C(n_23),
.D(n_22),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_33),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_136),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_3),
.B(n_4),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_116),
.B(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_5),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_146),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_145),
.B(n_147),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_5),
.B(n_6),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_7),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_131),
.C(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_161),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_137),
.C(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_147),
.Y(n_171)
);

AOI321xp33_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_144),
.A3(n_150),
.B1(n_149),
.B2(n_145),
.C(n_134),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_153),
.C(n_148),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_128),
.B1(n_156),
.B2(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_154),
.B1(n_165),
.B2(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_161),
.C(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_171),
.B(n_166),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_130),
.B1(n_21),
.B2(n_20),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_177),
.B1(n_173),
.B2(n_175),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_9),
.B(n_11),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_12),
.B(n_13),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_15),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_12),
.B(n_13),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_15),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_14),
.Y(n_184)
);


endmodule