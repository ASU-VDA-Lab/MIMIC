module fake_jpeg_30484_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_21),
.Y(n_61)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_49),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_18),
.B(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_27),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_19),
.Y(n_73)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_58),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_63),
.B(n_81),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_83),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_91),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_54),
.B1(n_53),
.B2(n_48),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_88),
.B1(n_77),
.B2(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_31),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_41),
.B(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_29),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_29),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_28),
.B(n_14),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_101),
.B1(n_109),
.B2(n_112),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_66),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_83),
.B1(n_74),
.B2(n_72),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_68),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_86),
.B(n_76),
.C(n_85),
.D(n_10),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_91),
.B1(n_74),
.B2(n_73),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_59),
.B1(n_67),
.B2(n_78),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_114),
.B1(n_98),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_146),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_85),
.B1(n_67),
.B2(n_59),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_143),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_111),
.C(n_110),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_73),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_105),
.C(n_117),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_86),
.Y(n_141)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_71),
.B1(n_85),
.B2(n_89),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_65),
.B1(n_80),
.B2(n_76),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_120),
.B(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_156),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_103),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_165),
.Y(n_170)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_94),
.B1(n_109),
.B2(n_116),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_168),
.B1(n_135),
.B2(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_108),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_102),
.B1(n_107),
.B2(n_65),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_153),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_180),
.B1(n_148),
.B2(n_151),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_144),
.C(n_142),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_175),
.C(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_133),
.C(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_138),
.C(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_128),
.B1(n_127),
.B2(n_140),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_158),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_190),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_151),
.B(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_192),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_188),
.B(n_193),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_153),
.B1(n_152),
.B2(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_155),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_176),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_159),
.C(n_157),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_175),
.C(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_150),
.Y(n_198)
);

OAI211xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_147),
.B(n_167),
.C(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_208),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_204),
.C(n_206),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_179),
.B1(n_176),
.B2(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_181),
.C(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_169),
.B1(n_173),
.B2(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_197),
.Y(n_212)
);

OAI322xp33_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_187),
.A3(n_182),
.B1(n_13),
.B2(n_12),
.C1(n_14),
.C2(n_161),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_206),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_202),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_220),
.B(n_221),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_204),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_222),
.A2(n_211),
.B(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_216),
.B(n_13),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_5),
.B(n_6),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_228),
.B(n_5),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_216),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_227),
.C(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_230),
.Y(n_233)
);


endmodule