module real_jpeg_1693_n_21 (n_17, n_8, n_0, n_95, n_2, n_10, n_9, n_12, n_97, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_96, n_16, n_15, n_13, n_21);

input n_17;
input n_8;
input n_0;
input n_95;
input n_2;
input n_10;
input n_9;
input n_12;
input n_97;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_96;
input n_16;
input n_15;
input n_13;

output n_21;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_0),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_10),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_5),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_5),
.B(n_18),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_10),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_7),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_10),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_9),
.B(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

AOI221xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.C(n_30),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_34),
.B(n_40),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_26),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_10),
.B(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_11),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_52),
.B2(n_53),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_12),
.A2(n_52),
.B1(n_77),
.B2(n_85),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_95),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_96),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_97),
.Y(n_65)
);

AOI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_54),
.B1(n_76),
.B2(n_86),
.C(n_92),
.Y(n_21)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

NOR5xp2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.C(n_41),
.D(n_45),
.E(n_48),
.Y(n_24)
);

NOR5xp2_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_40),
.C(n_48),
.D(n_79),
.E(n_84),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_35),
.C(n_81),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_47),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_72),
.B(n_74),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_70),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_73),
.B(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_66),
.B(n_69),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);


endmodule