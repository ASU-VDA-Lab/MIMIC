module fake_jpeg_25474_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_7),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_29),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_32),
.B1(n_23),
.B2(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_32),
.B1(n_23),
.B2(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_38),
.B1(n_18),
.B2(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_68),
.Y(n_85)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_44),
.B1(n_36),
.B2(n_39),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_80),
.B1(n_91),
.B2(n_16),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_79),
.B1(n_43),
.B2(n_96),
.Y(n_106)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_32),
.B1(n_22),
.B2(n_23),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_22),
.B1(n_31),
.B2(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_39),
.B1(n_38),
.B2(n_30),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_38),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_96),
.B1(n_56),
.B2(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_38),
.B1(n_29),
.B2(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_21),
.A3(n_33),
.B1(n_42),
.B2(n_16),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_R g112 ( 
.A(n_95),
.B(n_31),
.Y(n_112)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_40),
.B1(n_43),
.B2(n_29),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_103),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_63),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_56),
.B1(n_51),
.B2(n_61),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_115),
.B1(n_81),
.B2(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_106),
.A2(n_116),
.B1(n_124),
.B2(n_18),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_121),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_40),
.C(n_62),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_81),
.C(n_76),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_113),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_33),
.B1(n_21),
.B2(n_60),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_48),
.B1(n_42),
.B2(n_55),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_90),
.B(n_85),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_9),
.B(n_10),
.Y(n_154)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_26),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_96),
.B(n_76),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_82),
.B(n_94),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_81),
.B1(n_74),
.B2(n_77),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_131),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_71),
.B1(n_73),
.B2(n_82),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_60),
.C(n_55),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_140),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_26),
.C(n_27),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_112),
.B(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_149),
.B(n_102),
.Y(n_174)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_150),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_73),
.B1(n_21),
.B2(n_28),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_25),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_107),
.B1(n_120),
.B2(n_108),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_73),
.B1(n_16),
.B2(n_28),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_26),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_120),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_100),
.B1(n_109),
.B2(n_99),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_99),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_139),
.C(n_134),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_159),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_120),
.B(n_102),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_171),
.B(n_177),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_178),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_175),
.B1(n_142),
.B2(n_151),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_0),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_100),
.B(n_98),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_180),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_119),
.B1(n_105),
.B2(n_117),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_186),
.B1(n_1),
.B2(n_2),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_28),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_187),
.B1(n_8),
.B2(n_10),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_25),
.B1(n_27),
.B2(n_8),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_126),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_209),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_135),
.C(n_128),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_193),
.B(n_167),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_149),
.B(n_154),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_199),
.B(n_203),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_198),
.C(n_207),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_157),
.B1(n_156),
.B2(n_187),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_25),
.C(n_7),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_1),
.B(n_3),
.Y(n_203)
);

AOI22x1_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_216),
.B1(n_186),
.B2(n_183),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_163),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_9),
.C(n_13),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_166),
.C(n_181),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_214),
.C(n_170),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_4),
.B(n_5),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_4),
.B(n_5),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_9),
.C(n_13),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_175),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_233),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_240),
.B(n_241),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_179),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_242),
.B1(n_216),
.B2(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_212),
.C(n_192),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_236),
.C(n_194),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_182),
.C(n_178),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_167),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_237),
.B(n_239),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_169),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_188),
.B1(n_202),
.B2(n_199),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_232),
.B1(n_237),
.B2(n_233),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_263),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_210),
.C(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_220),
.C(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_199),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_214),
.CI(n_213),
.CON(n_261),
.SN(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_275),
.C(n_277),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_234),
.B(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_278),
.Y(n_286)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_274),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_259),
.B1(n_248),
.B2(n_241),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_229),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_220),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_239),
.C(n_231),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_200),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_235),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_264),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_201),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_260),
.B(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_280),
.A2(n_256),
.B1(n_247),
.B2(n_245),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_287),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_284),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_246),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_165),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_248),
.B(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_269),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_232),
.B1(n_261),
.B2(n_254),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_244),
.B1(n_267),
.B2(n_270),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_244),
.B1(n_200),
.B2(n_240),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_292),
.B1(n_289),
.B2(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_269),
.C(n_275),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_303),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_265),
.C(n_274),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_165),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_306),
.C(n_299),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_306),
.Y(n_311)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_301),
.B1(n_297),
.B2(n_169),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_285),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_314),
.A2(n_8),
.B(n_11),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_309),
.C(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_318),
.B(n_321),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_6),
.B(n_11),
.C(n_14),
.D(n_320),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_319),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_322),
.B(n_323),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_11),
.B(n_14),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_327),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_14),
.Y(n_329)
);

AOI31xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_6),
.A3(n_328),
.B(n_324),
.Y(n_330)
);


endmodule