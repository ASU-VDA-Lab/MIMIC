module fake_jpeg_3764_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_41),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_24),
.B1(n_22),
.B2(n_15),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_18),
.B(n_13),
.Y(n_40)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_22),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_52),
.B1(n_36),
.B2(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_56),
.B1(n_50),
.B2(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_54),
.B(n_65),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_62),
.B(n_19),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_54),
.B1(n_56),
.B2(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_17),
.B1(n_26),
.B2(n_44),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_47),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_26),
.Y(n_91)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_17),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_44),
.C(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_90),
.B1(n_92),
.B2(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AO221x1_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_95),
.B1(n_62),
.B2(n_79),
.C(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_77),
.B1(n_82),
.B2(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_0),
.Y(n_111)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_78),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_1),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_78),
.B(n_26),
.C(n_74),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_94),
.C(n_14),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_108),
.B(n_111),
.Y(n_115)
);

NOR2xp67_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_14),
.C(n_5),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_5),
.C(n_8),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_1),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_8),
.Y(n_118)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_120),
.Y(n_122)
);

AOI31xp67_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_102),
.A3(n_99),
.B(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.C(n_11),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_112),
.B1(n_4),
.B2(n_2),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_11),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_119),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_130),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_2),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_4),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_127),
.CI(n_128),
.CON(n_134),
.SN(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);


endmodule