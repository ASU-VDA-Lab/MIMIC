module fake_jpeg_22008_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_43),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_19),
.B1(n_26),
.B2(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_55),
.B1(n_23),
.B2(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_57),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_42),
.Y(n_67)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_75),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_56),
.B1(n_41),
.B2(n_48),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_50),
.A3(n_59),
.B1(n_22),
.B2(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_19),
.B1(n_17),
.B2(n_16),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_34),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_41),
.B1(n_42),
.B2(n_31),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_20),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_34),
.C(n_36),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_16),
.B(n_30),
.C(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_30),
.B1(n_29),
.B2(n_21),
.Y(n_100)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_107),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_82),
.B1(n_64),
.B2(n_61),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_50),
.B(n_53),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_96),
.B(n_67),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_81),
.B1(n_74),
.B2(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_67),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_53),
.B(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_105),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_77),
.B(n_59),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_11),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_15),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_130),
.B1(n_89),
.B2(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_120),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_122),
.B(n_90),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_97),
.B1(n_95),
.B2(n_88),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_92),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_103),
.C(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_106),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_1),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_99),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_68),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_136),
.B(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_147),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_135),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_98),
.B(n_95),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_145),
.C(n_146),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_2),
.Y(n_163)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_110),
.B1(n_106),
.B2(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_143),
.B1(n_112),
.B2(n_121),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_96),
.C(n_109),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_132),
.B1(n_147),
.B2(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_161),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_157),
.B(n_140),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_115),
.B(n_125),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_118),
.B(n_114),
.C(n_111),
.D(n_128),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_139),
.A3(n_136),
.B1(n_141),
.B2(n_143),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_162),
.B1(n_4),
.B2(n_5),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_127),
.C(n_15),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_14),
.C(n_13),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_138),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_140),
.B(n_139),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_173),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_144),
.B1(n_134),
.B2(n_5),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_158),
.C(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_153),
.B(n_154),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_2),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_160),
.C(n_163),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_184),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_5),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_175),
.B(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_192),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_6),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_184),
.C(n_182),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_6),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_183),
.B1(n_181),
.B2(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_188),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_179),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_7),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_196),
.C(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_9),
.B1(n_199),
.B2(n_202),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_9),
.Y(n_205)
);


endmodule