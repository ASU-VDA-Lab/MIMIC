module fake_jpeg_21170_n_296 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_26),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_23),
.B1(n_15),
.B2(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_27),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_57),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_27),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_66),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

OAI22x1_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_60),
.B1(n_55),
.B2(n_54),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_72),
.B1(n_74),
.B2(n_79),
.Y(n_91)
);

NOR2x1_ASAP7_75t_R g69 ( 
.A(n_50),
.B(n_33),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_33),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_29),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_80),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_28),
.B1(n_37),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_28),
.B1(n_37),
.B2(n_35),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_29),
.B1(n_23),
.B2(n_15),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_58),
.B1(n_41),
.B2(n_42),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_23),
.B1(n_15),
.B2(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_74),
.B1(n_78),
.B2(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_94),
.Y(n_110)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_97),
.B(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_99),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_56),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_92),
.B1(n_96),
.B2(n_48),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_67),
.B1(n_71),
.B2(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_118),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_82),
.C(n_71),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_33),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_83),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_83),
.B1(n_84),
.B2(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_128),
.B1(n_129),
.B2(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_84),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_125),
.B(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_129),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_75),
.B(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_76),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_18),
.B1(n_12),
.B2(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_30),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_133),
.B(n_135),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_137),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_103),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_148),
.B(n_149),
.Y(n_161)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_141),
.Y(n_159)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_92),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_32),
.B(n_13),
.C(n_25),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_20),
.B(n_33),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_20),
.B(n_33),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_155),
.B(n_156),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_17),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_117),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_115),
.B1(n_117),
.B2(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_164),
.C(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_115),
.C(n_107),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_128),
.B1(n_113),
.B2(n_25),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_113),
.B(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_146),
.B1(n_131),
.B2(n_144),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_179),
.B1(n_141),
.B2(n_157),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_17),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_132),
.A2(n_149),
.B1(n_153),
.B2(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_177),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_17),
.B(n_25),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_96),
.B1(n_48),
.B2(n_24),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_30),
.Y(n_178)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_63),
.B1(n_62),
.B2(n_53),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_24),
.B1(n_18),
.B2(n_13),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_16),
.B(n_18),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_159),
.B1(n_173),
.B2(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_203),
.B1(n_179),
.B2(n_162),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_155),
.A3(n_156),
.B1(n_137),
.B2(n_16),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_63),
.C(n_62),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_200),
.C(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_53),
.C(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_167),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_32),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_11),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_10),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_183),
.B(n_1),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_175),
.C(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_215),
.C(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_175),
.C(n_161),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_161),
.B1(n_168),
.B2(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_220),
.B1(n_222),
.B2(n_191),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_183),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_186),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_183),
.B1(n_176),
.B2(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_10),
.B1(n_8),
.B2(n_2),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_53),
.B(n_10),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_0),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_8),
.B(n_1),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_0),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_32),
.C(n_22),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_233),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_207),
.B1(n_185),
.B2(n_190),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_191),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_199),
.B1(n_201),
.B2(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_237),
.B1(n_241),
.B2(n_220),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_209),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_240),
.B(n_242),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_204),
.C(n_199),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_215),
.C(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_217),
.B(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_237),
.C(n_22),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_218),
.C(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_236),
.B(n_229),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_2),
.B(n_3),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_32),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_225),
.C(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_221),
.B1(n_223),
.B2(n_213),
.Y(n_253)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_232),
.B(n_239),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_267),
.C(n_32),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_22),
.C(n_19),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_22),
.B(n_32),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_246),
.C(n_248),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_265),
.A2(n_251),
.B1(n_253),
.B2(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_272),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_253),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_277),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_275),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_6),
.C(n_7),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_266),
.C(n_267),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_6),
.B(n_7),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

BUFx4f_ASAP7_75t_SL g283 ( 
.A(n_270),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_269),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_283),
.B(n_284),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_278),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_286),
.C(n_279),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_289),
.B(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_271),
.C(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_294),
.B(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_6),
.Y(n_296)
);


endmodule