module fake_jpeg_29802_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_76),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_61),
.B(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_1),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_63),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_77),
.B(n_22),
.C(n_25),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_61),
.B1(n_63),
.B2(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_50),
.B1(n_61),
.B2(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_54),
.B1(n_68),
.B2(n_65),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_80),
.B1(n_76),
.B2(n_79),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_48),
.B1(n_69),
.B2(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_62),
.B1(n_64),
.B2(n_53),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_55),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_16),
.B(n_35),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_111),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_75),
.B(n_2),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_20),
.B1(n_46),
.B2(n_44),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_19),
.B1(n_43),
.B2(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_18),
.B(n_39),
.C(n_36),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_105),
.B1(n_101),
.B2(n_113),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_15),
.B1(n_32),
.B2(n_31),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_10),
.Y(n_141)
);

NAND2x1p5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_8),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_128),
.B1(n_11),
.B2(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_9),
.Y(n_135)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_141),
.B(n_143),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_9),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_139),
.C(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_28),
.C(n_30),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_12),
.C(n_13),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_127),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_11),
.B(n_29),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_125),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_136),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_134),
.B1(n_142),
.B2(n_146),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_152),
.C(n_118),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_147),
.B1(n_151),
.B2(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_157),
.B1(n_134),
.B2(n_148),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_133),
.B(n_150),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_150),
.Y(n_162)
);


endmodule