module fake_jpeg_31206_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_74),
.B1(n_46),
.B2(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_72),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_17),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_24),
.C(n_29),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_50),
.C(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_39),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_23),
.B1(n_25),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_23),
.B1(n_25),
.B2(n_36),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_76),
.B(n_91),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_71),
.B1(n_74),
.B2(n_37),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_35),
.B1(n_20),
.B2(n_38),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_19),
.B(n_31),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_79),
.B(n_87),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_69),
.B1(n_49),
.B2(n_41),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_80),
.A2(n_104),
.A3(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_89),
.Y(n_143)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_50),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_97),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_17),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_65),
.Y(n_94)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_31),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_112),
.C(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_46),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_34),
.B1(n_38),
.B2(n_35),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_32),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_31),
.B(n_19),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_26),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_19),
.A3(n_31),
.B1(n_18),
.B2(n_20),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_17),
.B1(n_19),
.B2(n_31),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_34),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_19),
.B(n_33),
.C(n_26),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_64),
.B(n_32),
.C(n_15),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_32),
.C(n_37),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_93),
.B1(n_38),
.B2(n_35),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_32),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_106),
.B(n_105),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_131),
.B1(n_146),
.B2(n_40),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_82),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_109),
.B1(n_47),
.B2(n_40),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_80),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_91),
.A2(n_28),
.B(n_33),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_90),
.B(n_18),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_28),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_136),
.C(n_143),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_80),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_89),
.B1(n_110),
.B2(n_112),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_172),
.B1(n_120),
.B2(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_89),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_152),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_96),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_157),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_156),
.A2(n_158),
.B1(n_166),
.B2(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_93),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_175),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_102),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_90),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_170),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_104),
.C(n_94),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_146),
.B1(n_140),
.B2(n_125),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_105),
.B1(n_86),
.B2(n_116),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_106),
.B1(n_81),
.B2(n_107),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_107),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_141),
.B(n_18),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_173),
.A2(n_117),
.B(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_88),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_122),
.A2(n_36),
.B1(n_84),
.B2(n_116),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_84),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_118),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_196),
.B1(n_202),
.B2(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_193),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_185),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_154),
.C(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_18),
.C(n_13),
.Y(n_236)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_171),
.B(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_138),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_119),
.B1(n_138),
.B2(n_127),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_208),
.B1(n_172),
.B2(n_174),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_141),
.B(n_127),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_201),
.B(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_120),
.B1(n_119),
.B2(n_142),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_130),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_207),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_130),
.B(n_123),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_47),
.B1(n_44),
.B2(n_36),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_148),
.A2(n_44),
.B1(n_36),
.B2(n_45),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_148),
.A2(n_123),
.B(n_45),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_45),
.B1(n_18),
.B2(n_15),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_151),
.B(n_14),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_149),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_220),
.B(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_215),
.B(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_168),
.B(n_175),
.Y(n_220)
);

AO32x1_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_162),
.A3(n_173),
.B1(n_156),
.B2(n_157),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_240),
.B1(n_181),
.B2(n_207),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_173),
.B(n_174),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_232),
.B(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_228),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_153),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_234),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_203),
.A2(n_153),
.B1(n_160),
.B2(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_237),
.C(n_197),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_12),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_11),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_185),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_189),
.B(n_183),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_235),
.B(n_214),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_221),
.B(n_227),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_247),
.B1(n_258),
.B2(n_213),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_200),
.B1(n_190),
.B2(n_202),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_252),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_254),
.B(n_217),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_186),
.C(n_190),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_206),
.B1(n_197),
.B2(n_199),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_255),
.A2(n_265),
.B1(n_240),
.B2(n_220),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_197),
.B1(n_186),
.B2(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_188),
.C(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_263),
.C(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_188),
.C(n_179),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_210),
.B1(n_11),
.B2(n_2),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_274),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_279),
.B1(n_244),
.B2(n_258),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_211),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_273),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_215),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_212),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_285),
.B(n_0),
.C(n_3),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_225),
.C(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_287),
.C(n_257),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_283),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_218),
.B1(n_222),
.B2(n_223),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_280),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_216),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_284),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_SL g283 ( 
.A(n_249),
.B(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_0),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_233),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_293),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_272),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_255),
.B1(n_264),
.B2(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_247),
.B1(n_256),
.B2(n_242),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_256),
.B1(n_254),
.B2(n_250),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_297),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_304),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_250),
.B1(n_252),
.B2(n_263),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_298),
.B(n_305),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_0),
.C(n_1),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_284),
.C(n_281),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_274),
.B(n_286),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_308),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_278),
.CI(n_297),
.CON(n_308),
.SN(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_277),
.B(n_290),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_313),
.B(n_294),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_287),
.C(n_272),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_320),
.C(n_291),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g313 ( 
.A(n_289),
.B(n_283),
.Y(n_313)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_270),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_319),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_325),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_308),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_309),
.A2(n_316),
.B(n_311),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_323),
.A2(n_324),
.B(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_288),
.C(n_293),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_303),
.B1(n_305),
.B2(n_282),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_295),
.C(n_282),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_319),
.B(n_295),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_335),
.B(n_5),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_328),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_336),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_310),
.B(n_307),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_314),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_339),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_312),
.Y(n_340)
);

AOI31xp33_ASAP7_75t_L g344 ( 
.A1(n_340),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_317),
.A3(n_330),
.B1(n_296),
.B2(n_324),
.C1(n_308),
.C2(n_299),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g347 ( 
.A1(n_341),
.A2(n_343),
.A3(n_344),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_280),
.A3(n_298),
.B1(n_276),
.B2(n_322),
.C1(n_8),
.C2(n_4),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_345),
.B(n_6),
.Y(n_348)
);

AOI31xp33_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_349),
.A3(n_9),
.B(n_10),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_348),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_8),
.C(n_9),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_350),
.C(n_342),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_345),
.Y(n_353)
);


endmodule