module fake_jpeg_8063_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_46),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_57),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_53),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_19),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_30),
.B1(n_25),
.B2(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_21),
.B1(n_19),
.B2(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_26),
.B1(n_34),
.B2(n_23),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_42),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_83),
.B(n_88),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_42),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_80),
.C(n_20),
.Y(n_103)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_79),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_49),
.B(n_56),
.C(n_38),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_44),
.B(n_42),
.C(n_45),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_23),
.B1(n_29),
.B2(n_17),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_96),
.B1(n_97),
.B2(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_60),
.B1(n_57),
.B2(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_96),
.Y(n_127)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_29),
.B1(n_23),
.B2(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_26),
.B1(n_29),
.B2(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_101),
.B(n_105),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_64),
.B1(n_51),
.B2(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_112),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_79),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_27),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_113),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_64),
.B1(n_69),
.B2(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_58),
.B1(n_72),
.B2(n_18),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_80),
.C(n_74),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_88),
.C(n_74),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_72),
.B1(n_43),
.B2(n_40),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_27),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_120),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_93),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_127),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_79),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_83),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_100),
.B(n_101),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_136),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_133),
.A2(n_145),
.B(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_144),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_33),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_111),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_147),
.C(n_149),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_83),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_45),
.B(n_37),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_72),
.B(n_93),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_50),
.C(n_37),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_104),
.C(n_99),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_90),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_106),
.A2(n_45),
.B(n_37),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_45),
.B(n_84),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_102),
.B1(n_125),
.B2(n_124),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_157),
.A2(n_161),
.B1(n_164),
.B2(n_166),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_175),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_113),
.B(n_99),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_162),
.B(n_165),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_122),
.B1(n_110),
.B2(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_112),
.B1(n_110),
.B2(n_100),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_123),
.B(n_115),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_81),
.B1(n_121),
.B2(n_115),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_120),
.B1(n_119),
.B2(n_93),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_120),
.B1(n_114),
.B2(n_95),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_89),
.B1(n_84),
.B2(n_95),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_139),
.B1(n_133),
.B2(n_143),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_153),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_130),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_31),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_148),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_43),
.B1(n_40),
.B2(n_36),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_142),
.C(n_149),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_33),
.B(n_35),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_130),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_185),
.A2(n_201),
.B(n_204),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_194),
.C(n_138),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_150),
.B1(n_128),
.B2(n_135),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_207),
.B(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_167),
.C(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_135),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

XOR2x2_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_147),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_200),
.B(n_28),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_132),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_132),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_209),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_33),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_205),
.B(n_197),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_180),
.CI(n_178),
.CON(n_213),
.SN(n_213)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_213),
.B(n_24),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_200),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_237),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_209),
.A2(n_167),
.B1(n_157),
.B2(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_173),
.B1(n_161),
.B2(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_165),
.B(n_174),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_224),
.B(n_190),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_178),
.B1(n_134),
.B2(n_152),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_225),
.B1(n_232),
.B2(n_233),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_156),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_152),
.B1(n_179),
.B2(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_141),
.B1(n_181),
.B2(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_229),
.C(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_33),
.C(n_35),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_185),
.B1(n_202),
.B2(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_28),
.B1(n_24),
.B2(n_33),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_33),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_241),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_192),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_248),
.C(n_257),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_204),
.B1(n_190),
.B2(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_254),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_186),
.C(n_191),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_186),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_217),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_229),
.C(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_0),
.C(n_1),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_0),
.C(n_1),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_245),
.B(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

AO221x1_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_235),
.B1(n_232),
.B2(n_233),
.C(n_236),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_265),
.B1(n_269),
.B2(n_271),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_219),
.B1(n_234),
.B2(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_225),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_266),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_213),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_273),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_244),
.A2(n_221),
.B(n_213),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_237),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_240),
.B(n_9),
.CI(n_15),
.CON(n_277),
.SN(n_277)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_11),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_243),
.C(n_241),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_285),
.C(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_273),
.A2(n_260),
.B1(n_261),
.B2(n_249),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_289),
.B1(n_277),
.B2(n_10),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_249),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_288),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_11),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_248),
.C(n_257),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_254),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_292),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_16),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_8),
.C(n_14),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_276),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_304),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_262),
.Y(n_300)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_0),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_279),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_303),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_277),
.B1(n_279),
.B2(n_271),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_288),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_265),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_307),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_281),
.C(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_297),
.C(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_7),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_295),
.B(n_10),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_7),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_10),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_320),
.B(n_321),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_319),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_7),
.B(n_14),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_6),
.B(n_13),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_323),
.B1(n_12),
.B2(n_16),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_12),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_314),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_324),
.B(n_317),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_323),
.C(n_311),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.B(n_329),
.Y(n_332)
);

AOI321xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_326),
.A3(n_12),
.B1(n_2),
.B2(n_4),
.C(n_1),
.Y(n_333)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_0),
.B(n_2),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_4),
.Y(n_335)
);


endmodule