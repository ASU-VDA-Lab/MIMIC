module fake_jpeg_6185_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_27),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_47),
.B1(n_26),
.B2(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_59),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_56),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_17),
.B1(n_23),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_25),
.B1(n_16),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_55),
.B1(n_22),
.B2(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_25),
.B1(n_16),
.B2(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_30),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_20),
.B1(n_1),
.B2(n_3),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_21),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_41),
.B(n_26),
.C(n_31),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_38),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_56),
.B(n_61),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_46),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_73),
.B1(n_42),
.B2(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_59),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_24),
.C(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_72),
.Y(n_81)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_15),
.B1(n_20),
.B2(n_29),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_46),
.B1(n_54),
.B2(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_29),
.B1(n_20),
.B2(n_26),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_52),
.B1(n_58),
.B2(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_84),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_93),
.B1(n_96),
.B2(n_52),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_58),
.B1(n_51),
.B2(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_100),
.B(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_119),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_65),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_91),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_65),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_75),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_96),
.C(n_85),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_109),
.B1(n_119),
.B2(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_71),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_48),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_108),
.C(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_132),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_85),
.B1(n_79),
.B2(n_52),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_45),
.A3(n_53),
.B1(n_51),
.B2(n_14),
.C1(n_11),
.C2(n_50),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_78),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_117),
.B(n_103),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_151),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_108),
.B(n_114),
.C(n_113),
.D(n_107),
.Y(n_142)
);

OA21x2_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_149),
.B(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_146),
.C(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_102),
.C(n_118),
.Y(n_148)
);

AOI21x1_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_64),
.B(n_60),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_76),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_164),
.B(n_147),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_122),
.B1(n_140),
.B2(n_138),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_162),
.A2(n_175),
.B1(n_176),
.B2(n_0),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_128),
.B1(n_133),
.B2(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

OAI322xp33_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_125),
.A3(n_128),
.B1(n_129),
.B2(n_123),
.C1(n_130),
.C2(n_137),
.Y(n_165)
);

AOI321xp33_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_147),
.A3(n_148),
.B1(n_153),
.B2(n_141),
.C(n_14),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_125),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_64),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_78),
.B1(n_72),
.B2(n_60),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_78),
.B1(n_72),
.B2(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_185),
.C(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_11),
.C(n_1),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_182),
.C(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_172),
.C(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_3),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_5),
.C(n_6),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_200),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_185),
.B(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_174),
.C(n_170),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_8),
.C(n_9),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_7),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_187),
.C(n_8),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_209),
.C(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_183),
.B1(n_177),
.B2(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_207),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_7),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_199),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_202),
.C(n_208),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_217),
.B(n_195),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_201),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_215),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_214),
.B(n_9),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_10),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_10),
.C(n_225),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.Y(n_229)
);


endmodule