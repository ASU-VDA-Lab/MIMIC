module real_jpeg_7116_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_1),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_1),
.A2(n_205),
.B(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_1),
.B(n_182),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_1),
.B(n_364),
.C(n_367),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_1),
.A2(n_78),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_1),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_1),
.B(n_138),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_1),
.A2(n_27),
.B1(n_407),
.B2(n_415),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_37),
.B1(n_40),
.B2(n_45),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_2),
.A2(n_45),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_2),
.A2(n_45),
.B1(n_78),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_45),
.B1(n_141),
.B2(n_224),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_121),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_121),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_3),
.A2(n_121),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_5),
.A2(n_103),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_5),
.A2(n_187),
.B1(n_249),
.B2(n_286),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_5),
.A2(n_286),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_5),
.A2(n_286),
.B1(n_396),
.B2(n_397),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_77),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_28),
.B1(n_77),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_77),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_49),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_49),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_7),
.A2(n_49),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_8),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_8),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_8),
.Y(n_302)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_12),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_12),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_12),
.A2(n_143),
.B1(n_179),
.B2(n_276),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_12),
.A2(n_29),
.B1(n_179),
.B2(n_390),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_12),
.A2(n_54),
.B1(n_179),
.B2(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_13),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_13),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_14),
.A2(n_103),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_14),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_14),
.A2(n_123),
.B1(n_283),
.B2(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_14),
.A2(n_54),
.B1(n_283),
.B2(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_14),
.A2(n_283),
.B1(n_408),
.B2(n_410),
.Y(n_407)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_15),
.Y(n_492)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_16),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_17),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_490),
.B(n_493),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_478),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI31xp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_211),
.A3(n_234),
.B(n_475),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_190),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_23),
.B(n_190),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_113),
.C(n_153),
.Y(n_23)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_24),
.B(n_113),
.CI(n_153),
.CON(n_352),
.SN(n_352)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_79),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_26),
.B(n_81),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_26),
.A2(n_80),
.B1(n_81),
.B2(n_112),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_26),
.A2(n_46),
.B1(n_80),
.B2(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_27),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_27),
.A2(n_257),
.B1(n_263),
.B2(n_267),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_27),
.A2(n_267),
.B(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_27),
.A2(n_162),
.B(n_389),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_27),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_27),
.A2(n_301),
.B1(n_395),
.B2(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_27),
.A2(n_36),
.B(n_299),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_31),
.Y(n_272)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_33),
.Y(n_419)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_36),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_43),
.Y(n_409)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_44),
.Y(n_262)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_44),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_46),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_57),
.B(n_72),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_48),
.A2(n_58),
.B1(n_73),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_51),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_125)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_52),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_52),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_52),
.Y(n_383)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_57),
.B(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_57),
.A2(n_146),
.B(n_147),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_57),
.A2(n_72),
.B(n_147),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_57),
.A2(n_146),
.B1(n_151),
.B2(n_169),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_57),
.A2(n_459),
.B(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_58),
.A2(n_73),
.B1(n_369),
.B2(n_372),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_58),
.A2(n_73),
.B1(n_372),
.B2(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_58),
.A2(n_73),
.B1(n_381),
.B2(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_59)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_60),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_67),
.Y(n_367)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_100),
.B(n_105),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_82),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_82),
.A2(n_182),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_82),
.A2(n_182),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_83),
.A2(n_176),
.B(n_181),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_83),
.A2(n_111),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_83),
.A2(n_111),
.B1(n_176),
.B2(n_285),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_83),
.A2(n_485),
.B(n_486),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_95),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_95),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_95),
.Y(n_444)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_96),
.Y(n_279)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_96),
.Y(n_335)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_98),
.Y(n_436)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_100),
.B(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_102),
.Y(n_287)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_105),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_109),
.Y(n_233)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_111),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_111),
.A2(n_201),
.B(n_207),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_144),
.B(n_152),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_144),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_124),
.B1(n_138),
.B2(n_139),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_125),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_131)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_124),
.B(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_124),
.A2(n_139),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_124),
.A2(n_222),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_124),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_124),
.A2(n_138),
.B1(n_332),
.B2(n_443),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_124),
.A2(n_138),
.B(n_483),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_125),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_125),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_125),
.A2(n_294),
.B1(n_295),
.B2(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_126),
.Y(n_371)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_127),
.Y(n_438)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_129),
.Y(n_432)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_186),
.Y(n_197)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g427 ( 
.A1(n_143),
.A2(n_428),
.A3(n_430),
.B1(n_433),
.B2(n_437),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_145),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_146),
.B(n_370),
.Y(n_405)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_148),
.Y(n_439)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_191),
.CI(n_210),
.CON(n_190),
.SN(n_190)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_174),
.C(n_183),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_154),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_166),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_155),
.A2(n_166),
.B1(n_167),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_155),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_157),
.A2(n_258),
.B(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_158),
.Y(n_303)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_164),
.Y(n_415)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_170),
.Y(n_447)
);

INVx5_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_172),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_174),
.A2(n_175),
.B1(n_183),
.B2(n_184),
.Y(n_346)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_190),
.B(n_213),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_200),
.B2(n_209),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_199),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_194),
.B(n_219),
.C(n_227),
.Y(n_487)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_199),
.C(n_200),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_197),
.A2(n_223),
.B(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_209),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_200),
.B(n_214),
.C(n_217),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_212),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_227),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_223),
.Y(n_483)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_229),
.Y(n_485)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_353),
.B(n_469),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_338),
.C(n_350),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_317),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_237),
.A2(n_471),
.B(n_472),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_305),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_238),
.B(n_305),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_288),
.C(n_297),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_239),
.B(n_337),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_273),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_240),
.B(n_274),
.C(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_256),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_241),
.B(n_256),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_245),
.A3(n_246),
.B1(n_248),
.B2(n_253),
.Y(n_241)
);

INVx4_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_261),
.Y(n_390)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_270),
.Y(n_396)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_271),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_297),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.C(n_293),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_289),
.B(n_290),
.CI(n_293),
.CON(n_319),
.SN(n_319)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_304),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_302),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_315),
.C(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_336),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_318),
.B(n_336),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_319),
.B(n_467),
.Y(n_466)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_319),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_320),
.B(n_321),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_328),
.C(n_330),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_322),
.A2(n_323),
.B1(n_328),
.B2(n_329),
.Y(n_454)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_330),
.B(n_454),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

A2O1A1O1Ixp25_ASAP7_75t_L g469 ( 
.A1(n_338),
.A2(n_350),
.B(n_470),
.C(n_473),
.D(n_474),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_349),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_339),
.B(n_349),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_343),
.C(n_348),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_345),
.B1(n_347),
.B2(n_348),
.Y(n_342)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_345),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_351),
.B(n_352),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_352),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_464),
.B(n_468),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_449),
.B(n_463),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_423),
.B(n_448),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_391),
.B(n_422),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_376),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_358),
.B(n_376),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_368),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_368),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_434),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_SL g443 ( 
.A1(n_370),
.A2(n_433),
.B(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_388),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_387),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_387),
.C(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_380),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_403),
.B(n_421),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_402),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_402),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_396),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_413),
.B(n_420),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_405),
.B(n_406),
.Y(n_420)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx4_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_425),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_441),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_442),
.C(n_445),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_440),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_440),
.Y(n_457)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_450),
.B(n_451),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_456),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_458),
.C(n_461),
.Y(n_465)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_461),
.B2(n_462),
.Y(n_456)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_457),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_458),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_466),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_488),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_481),
.Y(n_489)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_481),
.Y(n_498)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_484),
.CI(n_487),
.CON(n_481),
.SN(n_481)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx13_ASAP7_75t_L g495 ( 
.A(n_492),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);


endmodule