module fake_netlist_5_1510_n_190 (n_16, n_0, n_12, n_9, n_25, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_190);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_190;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_146;
wire n_136;
wire n_86;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_101;
wire n_75;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_29;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_188;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_154;
wire n_148;
wire n_71;
wire n_138;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_27;
wire n_170;
wire n_64;
wire n_77;
wire n_102;
wire n_161;
wire n_106;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVxp67_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_18),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AND3x1_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_0),
.C(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_4),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2x1p5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_49),
.B1(n_65),
.B2(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_44),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_79),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_64),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_54),
.B1(n_63),
.B2(n_52),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_53),
.C(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_81),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_73),
.B(n_71),
.C(n_74),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_72),
.B(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_71),
.B1(n_77),
.B2(n_83),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_90),
.Y(n_105)
);

OAI21x1_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_95),
.B(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_85),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_102),
.B(n_99),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_93),
.B(n_96),
.C(n_94),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_94),
.B(n_96),
.C(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_92),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_108),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_83),
.B1(n_68),
.B2(n_77),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_46),
.B1(n_77),
.B2(n_85),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_92),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_73),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_122),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_128),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_117),
.Y(n_146)
);

NAND2x1_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_126),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_122),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_123),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_123),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_125),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_146),
.C(n_125),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_120),
.B1(n_144),
.B2(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_154),
.C(n_156),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_143),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_147),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_138),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_151),
.C(n_136),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_136),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_120),
.Y(n_169)
);

NOR2x1p5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_51),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_48),
.C(n_47),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_120),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_54),
.C(n_47),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_171),
.B(n_159),
.C(n_160),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

OR5x1_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_166),
.C(n_173),
.D(n_172),
.E(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_54),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_75),
.C(n_110),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_71),
.B(n_106),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_86),
.C(n_92),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_177),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_10),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_180),
.A3(n_176),
.B1(n_179),
.B2(n_181),
.C1(n_86),
.C2(n_102),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g187 ( 
.A(n_185),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_183),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_186),
.B1(n_188),
.B2(n_89),
.C(n_88),
.Y(n_190)
);


endmodule