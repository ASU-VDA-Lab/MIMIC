module fake_netlist_1_4811_n_588 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_588);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_588;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_39), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_70), .Y(n_84) );
BUFx10_ASAP7_75t_L g85 ( .A(n_30), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_34), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_28), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_56), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_5), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_77), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_36), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_26), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_69), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_59), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_54), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_65), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_52), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_32), .Y(n_102) );
BUFx2_ASAP7_75t_SL g103 ( .A(n_17), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_51), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_46), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_49), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_24), .Y(n_107) );
OR2x2_ASAP7_75t_L g108 ( .A(n_19), .B(n_72), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_42), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_81), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_48), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_50), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_15), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_7), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_31), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_64), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_6), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_120), .B(n_0), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_85), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_93), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_93), .Y(n_124) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_94), .A2(n_38), .B(n_79), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_85), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_119), .B(n_0), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_111), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_82), .B(n_1), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_91), .B(n_1), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_101), .A2(n_2), .B1(n_3), .B2(n_6), .Y(n_133) );
BUFx8_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_101), .A2(n_2), .B1(n_3), .B2(n_7), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_89), .B(n_8), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_83), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_84), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
OAI22xp5_ASAP7_75t_SL g143 ( .A1(n_116), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_98), .B(n_11), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_138), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_122), .B(n_86), .Y(n_149) );
INVxp67_ASAP7_75t_SL g150 ( .A(n_122), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_138), .A2(n_115), .B1(n_109), .B2(n_103), .Y(n_151) );
NAND2xp33_ASAP7_75t_L g152 ( .A(n_122), .B(n_87), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_122), .B(n_87), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_125), .A2(n_95), .B(n_117), .Y(n_155) );
OR2x2_ASAP7_75t_L g156 ( .A(n_136), .B(n_89), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_123), .A2(n_103), .B1(n_114), .B2(n_108), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_123), .A2(n_108), .B1(n_113), .B2(n_102), .Y(n_159) );
INVx4_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
NAND3xp33_ASAP7_75t_L g161 ( .A(n_124), .B(n_118), .C(n_90), .Y(n_161) );
INVx6_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_124), .A2(n_92), .B1(n_99), .B2(n_104), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_142), .A2(n_105), .B1(n_112), .B2(n_107), .Y(n_165) );
BUFx4f_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_136), .B(n_100), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_133), .A2(n_100), .B1(n_110), .B2(n_107), .Y(n_168) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_125), .A2(n_112), .B(n_110), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_136), .B(n_106), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_126), .B(n_145), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g172 ( .A1(n_121), .A2(n_106), .B1(n_97), .B2(n_88), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_145), .B(n_96), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_173), .A2(n_131), .B1(n_132), .B2(n_144), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_151), .A2(n_126), .B1(n_140), .B2(n_139), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_150), .B(n_88), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_153), .B(n_97), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_168), .A2(n_133), .B1(n_137), .B2(n_143), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_170), .B(n_144), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_160), .B(n_132), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_160), .B(n_121), .Y(n_185) );
NOR2xp33_ASAP7_75t_R g186 ( .A(n_152), .B(n_134), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g187 ( .A(n_160), .B(n_57), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_146), .A2(n_128), .B1(n_137), .B2(n_143), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
AND2x6_ASAP7_75t_SL g191 ( .A(n_149), .B(n_128), .Y(n_191) );
BUFx8_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_160), .B(n_134), .Y(n_193) );
O2A1O1Ixp5_ASAP7_75t_L g194 ( .A1(n_166), .A2(n_171), .B(n_167), .C(n_148), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_166), .B(n_134), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_166), .B(n_125), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_147), .B(n_47), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_166), .B(n_130), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_146), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_168), .A2(n_130), .B1(n_12), .B2(n_13), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_156), .B(n_130), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_156), .B(n_141), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_172), .B(n_141), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_148), .B(n_45), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_165), .B(n_141), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_159), .B(n_53), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_158), .B(n_11), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_173), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_196), .A2(n_169), .B(n_161), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_209), .B(n_163), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_209), .A2(n_173), .B1(n_161), .B2(n_162), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_169), .B(n_157), .Y(n_214) );
OAI21xp33_ASAP7_75t_L g215 ( .A1(n_182), .A2(n_173), .B(n_129), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_183), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_183), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_192), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_191), .B(n_173), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_205), .B(n_129), .Y(n_220) );
NOR2x1_ASAP7_75t_L g221 ( .A(n_176), .B(n_169), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_199), .A2(n_169), .B(n_141), .C(n_135), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_191), .B(n_162), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_185), .A2(n_202), .B(n_199), .Y(n_224) );
NOR3xp33_ASAP7_75t_L g225 ( .A(n_188), .B(n_173), .C(n_157), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_157), .B(n_162), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_209), .A2(n_162), .B1(n_173), .B2(n_141), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_174), .A2(n_162), .B(n_164), .Y(n_228) );
BUFx4f_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_175), .B(n_178), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_205), .B(n_141), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_179), .B(n_173), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_189), .A2(n_164), .B(n_55), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_189), .B(n_135), .Y(n_235) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_186), .B(n_135), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_177), .A2(n_164), .B(n_135), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_200), .B(n_12), .C(n_13), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_207), .B(n_14), .Y(n_239) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_187), .A2(n_164), .B(n_135), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_190), .B(n_135), .Y(n_241) );
NOR2xp33_ASAP7_75t_SL g242 ( .A(n_192), .B(n_129), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_190), .A2(n_129), .B(n_164), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_187), .A2(n_164), .B(n_44), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_181), .Y(n_245) );
CKINVDCx10_ASAP7_75t_R g246 ( .A(n_192), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_181), .A2(n_43), .B(n_78), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_212), .B(n_208), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_222), .A2(n_208), .B(n_203), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_214), .A2(n_206), .B(n_201), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_234), .A2(n_210), .B(n_194), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_233), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_245), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_235), .A2(n_193), .B(n_195), .Y(n_254) );
AOI21xp33_ASAP7_75t_L g255 ( .A1(n_221), .A2(n_204), .B(n_197), .Y(n_255) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_198), .A3(n_200), .B(n_210), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_217), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_180), .B1(n_210), .B2(n_16), .Y(n_258) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_180), .B(n_58), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_235), .A2(n_41), .B(n_76), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_218), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_211), .A2(n_40), .B(n_75), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_241), .A2(n_37), .B(n_74), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_212), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_219), .B(n_14), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_230), .B(n_15), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_223), .B(n_16), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_244), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_241), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_232), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_220), .Y(n_277) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_274), .A2(n_215), .B(n_220), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_268), .B(n_238), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_272), .A2(n_213), .B(n_227), .Y(n_280) );
CKINVDCx8_ASAP7_75t_R g281 ( .A(n_271), .Y(n_281) );
BUFx12f_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_268), .B(n_239), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_250), .A2(n_231), .B(n_236), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_258), .A2(n_239), .B1(n_225), .B2(n_223), .C(n_224), .Y(n_285) );
AOI21x1_ASAP7_75t_L g286 ( .A1(n_274), .A2(n_231), .B(n_237), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_261), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_261), .B(n_247), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_261), .B(n_226), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_261), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_250), .A2(n_228), .B(n_61), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_257), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_252), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_261), .B(n_18), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_261), .B(n_18), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_272), .A2(n_19), .B(n_20), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_249), .A2(n_21), .B(n_23), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_252), .B(n_80), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_257), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_249), .A2(n_25), .B(n_27), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_253), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_274), .A2(n_29), .B(n_33), .Y(n_302) );
INVx4_ASAP7_75t_SL g303 ( .A(n_282), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_299), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_299), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_293), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_301), .B(n_263), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_292), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_294), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_294), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_279), .B(n_248), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_295), .B(n_248), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_282), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_289), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_281), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_283), .B(n_253), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_316), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_316), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_321), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_324), .B(n_288), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_321), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_324), .B(n_256), .Y(n_334) );
INVxp33_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_306), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_326), .A2(n_285), .B1(n_273), .B2(n_263), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_309), .B(n_256), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_309), .B(n_256), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_310), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_314), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_303), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_326), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_318), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_317), .B(n_256), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_317), .B(n_256), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_313), .B(n_256), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_311), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_348), .B(n_313), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_349), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_352), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_336), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_350), .B(n_312), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_342), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_350), .B(n_323), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_353), .B(n_323), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_351), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_352), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_353), .B(n_259), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_335), .B(n_322), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_343), .B(n_355), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_343), .B(n_325), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_259), .Y(n_376) );
INVx4_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_355), .B(n_320), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_341), .B(n_303), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_337), .A2(n_289), .B1(n_296), .B2(n_288), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_334), .B(n_259), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_344), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_330), .B(n_303), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_331), .B(n_269), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_259), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_337), .A2(n_271), .B1(n_280), .B2(n_266), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_331), .B(n_303), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_347), .B(n_271), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_338), .B(n_288), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_339), .B(n_329), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_333), .B(n_329), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_339), .B(n_287), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_345), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_329), .B(n_287), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_354), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_333), .B(n_269), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_358), .B(n_271), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_357), .B(n_271), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_374), .B(n_357), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_363), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_366), .B(n_340), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_366), .B(n_340), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_359), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_391), .B(n_330), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_391), .B(n_330), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_392), .B(n_357), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_392), .B(n_340), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_367), .B(n_340), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_367), .B(n_351), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_368), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_403), .A2(n_290), .B(n_354), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_359), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_395), .B(n_332), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_394), .B(n_332), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g423 ( .A(n_377), .B(n_271), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_374), .B(n_356), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_360), .B(n_356), .Y(n_426) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_265), .B(n_300), .C(n_297), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_395), .B(n_332), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_364), .B(n_332), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_364), .B(n_332), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_359), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_378), .B(n_328), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_394), .B(n_332), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_360), .B(n_328), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_361), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_378), .B(n_328), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_393), .B(n_327), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_327), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_394), .B(n_327), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_394), .B(n_270), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_372), .B(n_290), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_371), .B(n_270), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_377), .B(n_265), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_371), .B(n_376), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_372), .B(n_284), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_382), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_377), .B(n_287), .Y(n_447) );
OAI21xp33_ASAP7_75t_SL g448 ( .A1(n_377), .A2(n_389), .B(n_379), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_383), .B(n_287), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_376), .B(n_270), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_375), .B(n_255), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_382), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_397), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_381), .B(n_251), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_375), .B(n_257), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_369), .B(n_277), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_373), .B(n_60), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_381), .B(n_251), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_384), .B(n_255), .Y(n_459) );
OAI21xp33_ASAP7_75t_SL g460 ( .A1(n_406), .A2(n_404), .B(n_380), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_437), .Y(n_461) );
AOI32xp33_ASAP7_75t_L g462 ( .A1(n_448), .A2(n_388), .A3(n_383), .B1(n_369), .B2(n_387), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_453), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_444), .B(n_402), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_425), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_412), .B(n_383), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_408), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_437), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_423), .B(n_383), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_451), .A2(n_390), .B(n_385), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_455), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_417), .B(n_361), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_447), .B(n_362), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_426), .B(n_402), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_409), .A2(n_384), .B1(n_386), .B2(n_398), .C(n_396), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_438), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_405), .B(n_370), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_405), .B(n_370), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_446), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_412), .B(n_396), .Y(n_486) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_455), .B(n_401), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_432), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_432), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_410), .B(n_386), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_444), .B(n_398), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_416), .B(n_401), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_413), .B(n_399), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_436), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_449), .B(n_385), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_436), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_414), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_411), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_457), .A2(n_390), .B1(n_387), .B2(n_362), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_456), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_414), .B(n_400), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_413), .B(n_390), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_429), .B(n_399), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_411), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_447), .B(n_400), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_480), .B(n_487), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_505), .B(n_430), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_470), .B(n_415), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_480), .B(n_415), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
NAND2xp33_ASAP7_75t_SL g514 ( .A(n_470), .B(n_475), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_490), .B(n_439), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_490), .B(n_439), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_464), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_491), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_492), .B(n_459), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_500), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_460), .A2(n_443), .B(n_419), .C(n_427), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_492), .A2(n_430), .B1(n_429), .B2(n_421), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_468), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_500), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
BUFx2_ASAP7_75t_SL g527 ( .A(n_488), .Y(n_527) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_472), .A2(n_458), .B1(n_454), .B2(n_442), .C1(n_450), .C2(n_441), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_496), .A2(n_456), .B(n_431), .C(n_420), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_496), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_504), .A2(n_428), .B1(n_421), .B2(n_433), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g532 ( .A1(n_462), .A2(n_443), .B(n_428), .Y(n_532) );
OAI22xp33_ASAP7_75t_SL g533 ( .A1(n_471), .A2(n_443), .B1(n_449), .B2(n_422), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_504), .A2(n_433), .B1(n_450), .B2(n_442), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_467), .B(n_422), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_469), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g537 ( .A1(n_479), .A2(n_443), .B(n_420), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_495), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_481), .B(n_435), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_535), .B(n_494), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_538), .Y(n_541) );
AOI211xp5_ASAP7_75t_L g542 ( .A1(n_522), .A2(n_502), .B(n_479), .C(n_477), .Y(n_542) );
OAI21xp33_ASAP7_75t_L g543 ( .A1(n_532), .A2(n_498), .B(n_465), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_530), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_527), .Y(n_545) );
NAND4xp75_ASAP7_75t_L g546 ( .A(n_508), .B(n_501), .C(n_477), .D(n_466), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_514), .A2(n_502), .B1(n_499), .B2(n_473), .C(n_485), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_528), .A2(n_495), .B1(n_486), .B2(n_489), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_520), .A2(n_474), .B1(n_497), .B2(n_478), .C(n_482), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_512), .A2(n_461), .B1(n_493), .B2(n_506), .C(n_484), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_539), .B(n_483), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_526), .A2(n_503), .B1(n_507), .B2(n_449), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_513), .A2(n_440), .B(n_361), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_535), .B(n_422), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_526), .A2(n_435), .B1(n_431), .B2(n_400), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_533), .B(n_440), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_528), .A2(n_458), .B1(n_454), .B2(n_370), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g558 ( .A1(n_537), .A2(n_362), .B1(n_267), .B2(n_302), .C(n_291), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_534), .A2(n_267), .B(n_262), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_537), .A2(n_264), .B1(n_260), .B2(n_276), .Y(n_560) );
AO21x1_ASAP7_75t_L g561 ( .A1(n_539), .A2(n_260), .B(n_277), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_518), .A2(n_276), .B1(n_264), .B2(n_254), .C(n_277), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g563 ( .A1(n_538), .A2(n_264), .B1(n_276), .B2(n_275), .C(n_67), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_519), .A2(n_276), .B1(n_275), .B2(n_66), .C(n_68), .Y(n_564) );
NOR3x1_ASAP7_75t_L g565 ( .A(n_511), .B(n_62), .C(n_63), .Y(n_565) );
NAND4xp25_ASAP7_75t_L g566 ( .A(n_531), .B(n_275), .C(n_71), .D(n_73), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_515), .B(n_516), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_529), .B(n_536), .C(n_524), .Y(n_568) );
NOR4xp75_ASAP7_75t_L g569 ( .A(n_517), .B(n_509), .C(n_523), .D(n_510), .Y(n_569) );
NOR3xp33_ASAP7_75t_L g570 ( .A(n_542), .B(n_543), .C(n_546), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_548), .A2(n_557), .B1(n_545), .B2(n_568), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_565), .B(n_566), .C(n_547), .D(n_563), .Y(n_572) );
NAND3xp33_ASAP7_75t_SL g573 ( .A(n_569), .B(n_561), .C(n_550), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_541), .B(n_544), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_567), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_573), .B(n_552), .C(n_564), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_575), .B(n_551), .Y(n_577) );
NAND3xp33_ASAP7_75t_SL g578 ( .A(n_570), .B(n_549), .C(n_556), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_578), .B(n_571), .C(n_572), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_577), .B(n_574), .Y(n_580) );
XNOR2xp5_ASAP7_75t_L g581 ( .A(n_579), .B(n_576), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_580), .B(n_553), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_582), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_581), .B1(n_525), .B2(n_521), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_584), .A2(n_540), .B(n_555), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_585), .A2(n_553), .B(n_554), .Y(n_586) );
NAND2x1_ASAP7_75t_L g587 ( .A(n_586), .B(n_560), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_587), .A2(n_559), .B1(n_562), .B2(n_558), .Y(n_588) );
endmodule