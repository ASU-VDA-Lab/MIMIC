module real_jpeg_28340_n_17 (n_8, n_0, n_2, n_338, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_338;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_0),
.A2(n_55),
.B1(n_57),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_0),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_77),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_77),
.Y(n_202)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_2),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_55),
.B1(n_57),
.B2(n_134),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_134),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_134),
.Y(n_271)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_4),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_4),
.A2(n_35),
.B1(n_55),
.B2(n_57),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_66),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_8),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_8),
.A2(n_31),
.B1(n_55),
.B2(n_57),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_9),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_55),
.B1(n_57),
.B2(n_169),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_169),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_169),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_10),
.B(n_57),
.Y(n_56)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_10),
.A2(n_56),
.B(n_57),
.C(n_61),
.D(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_10),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_10),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_81),
.B(n_85),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_25),
.B(n_119),
.C(n_120),
.D(n_124),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_10),
.B(n_25),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_23),
.B(n_24),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_103),
.Y(n_176)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_11),
.A2(n_57),
.B(n_62),
.C(n_63),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_12),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_12),
.A2(n_55),
.B1(n_57),
.B2(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_152),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_152),
.Y(n_298)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_55),
.B1(n_57),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_14),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_15),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_15),
.A2(n_55),
.B1(n_57),
.B2(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_84),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_84),
.Y(n_219)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_21),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_21),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_21),
.A2(n_26),
.B1(n_202),
.B2(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_21),
.A2(n_26),
.B1(n_34),
.B2(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_22),
.A2(n_28),
.B(n_103),
.C(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_24),
.A2(n_25),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_24),
.A2(n_57),
.A3(n_119),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_26),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_26),
.B(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_26),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_33),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_33),
.B(n_335),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_334),
.B(n_336),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_322),
.B(n_333),
.Y(n_39)
);

OAI321xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_286),
.A3(n_315),
.B1(n_320),
.B2(n_321),
.C(n_338),
.Y(n_40)
);

AOI321xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_236),
.A3(n_275),
.B1(n_280),
.B2(n_285),
.C(n_339),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_189),
.C(n_232),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_160),
.B(n_188),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_139),
.B(n_159),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_114),
.B(n_138),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_90),
.B(n_113),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_68),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_48),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_60),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_50),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_55),
.B(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_63),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_61),
.A2(n_63),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_61),
.A2(n_63),
.B1(n_252),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_67),
.A2(n_78),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_67),
.A2(n_156),
.B1(n_187),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_67),
.A2(n_156),
.B1(n_210),
.B2(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_67),
.A2(n_156),
.B(n_261),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_75),
.C(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_72),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_72),
.A2(n_120),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_72),
.A2(n_120),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_72),
.A2(n_120),
.B1(n_264),
.B2(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_72),
.A2(n_120),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_76),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_89),
.B1(n_133),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_81),
.A2(n_89),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_81),
.A2(n_208),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_81),
.A2(n_98),
.B(n_226),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_88),
.A2(n_95),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx5_ASAP7_75t_SL g225 ( 
.A(n_88),
.Y(n_225)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_103),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_112),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_99),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_98),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_106),
.B(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_107),
.B(n_111),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_104),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_116),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_130),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_127),
.C(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_126),
.A2(n_145),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_126),
.A2(n_197),
.B1(n_222),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_126),
.A2(n_197),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_153),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_154),
.C(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_148),
.C(n_150),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_201),
.B(n_203),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_149),
.A2(n_203),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_149),
.A2(n_243),
.B1(n_271),
.B2(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_149),
.A2(n_243),
.B1(n_298),
.B2(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_164),
.B(n_165),
.C(n_174),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_173),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_182),
.C(n_185),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_178),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_190),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_212),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_191),
.B(n_212),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_205),
.C(n_211),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_195),
.C(n_204),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_204),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B(n_199),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_211),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_209),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_223),
.C(n_231),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_218),
.C(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_219),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_227),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_233),
.B(n_234),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_256),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_248),
.C(n_255),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_248),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_247),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_239),
.Y(n_247)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_245),
.C(n_247),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_254),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_254),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_269),
.B(n_272),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_274),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_266),
.B1(n_267),
.B2(n_273),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_262),
.B(n_265),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_262),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_265),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_265),
.A2(n_288),
.B1(n_289),
.B2(n_300),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_273),
.C(n_274),
.Y(n_316)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_276),
.A2(n_281),
.B(n_284),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_303),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_303),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_300),
.C(n_301),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_299),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_296),
.C(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_293),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_294),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_296),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_307),
.C(n_311),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_297),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_299),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_306),
.C(n_314),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_302),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_308),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_313),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_326),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_328),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_331),
.C(n_332),
.Y(n_335)
);


endmodule