module fake_jpeg_26405_n_330 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_6),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_69),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_20),
.B1(n_18),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_36),
.B1(n_24),
.B2(n_28),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_26),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_29),
.B1(n_23),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_23),
.B1(n_18),
.B2(n_22),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_76),
.B1(n_79),
.B2(n_27),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_46),
.B1(n_17),
.B2(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_45),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_48),
.B(n_43),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_28),
.B1(n_24),
.B2(n_36),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_47),
.C(n_43),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_48),
.CI(n_36),
.CON(n_94),
.SN(n_94)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_36),
.B1(n_27),
.B2(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_89),
.B1(n_116),
.B2(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_47),
.B1(n_44),
.B2(n_36),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_117),
.B1(n_102),
.B2(n_109),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_97),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_96),
.B(n_104),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_28),
.B1(n_24),
.B2(n_43),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_80),
.B1(n_68),
.B2(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_0),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_0),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_111),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_54),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_78),
.A3(n_57),
.B1(n_50),
.B2(n_7),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_33),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_33),
.B1(n_32),
.B2(n_3),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_97),
.B1(n_98),
.B2(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_50),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_64),
.B1(n_80),
.B2(n_70),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_127),
.B1(n_138),
.B2(n_141),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_64),
.C(n_59),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_150),
.C(n_115),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_125),
.B1(n_137),
.B2(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_84),
.B1(n_83),
.B2(n_104),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_58),
.B(n_57),
.C(n_59),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_133),
.B(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_144),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_57),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_78),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_88),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_50),
.C(n_8),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_151),
.B(n_155),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_104),
.C(n_107),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_160),
.B(n_172),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_125),
.B1(n_127),
.B2(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_154),
.A2(n_165),
.B1(n_176),
.B2(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_133),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_175),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_128),
.B(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_92),
.B1(n_94),
.B2(n_99),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_181),
.B1(n_150),
.B2(n_126),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_163),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_88),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_166),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_94),
.B1(n_96),
.B2(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_91),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_94),
.B1(n_89),
.B2(n_117),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_183),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_97),
.B1(n_98),
.B2(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_100),
.B1(n_101),
.B2(n_108),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_101),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_174),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_103),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_105),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_108),
.B1(n_111),
.B2(n_110),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_108),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_119),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_180),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_142),
.B1(n_138),
.B2(n_122),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_119),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_122),
.A2(n_85),
.B1(n_81),
.B2(n_93),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_162),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_145),
.B(n_126),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_204),
.B(n_210),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_197),
.B1(n_200),
.B2(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_196),
.B(n_198),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_159),
.B1(n_161),
.B2(n_151),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_150),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_139),
.B1(n_137),
.B2(n_124),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_134),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_204),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_134),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_203),
.B(n_164),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_136),
.B(n_124),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_213),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_136),
.C(n_129),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.C(n_157),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_129),
.C(n_131),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_87),
.B(n_131),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_168),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_81),
.B1(n_143),
.B2(n_114),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_176),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_163),
.B1(n_169),
.B2(n_167),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_175),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_222),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_209),
.C(n_193),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_241),
.C(n_152),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_154),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_158),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_190),
.B(n_166),
.CI(n_158),
.CON(n_232),
.SN(n_232)
);

OAI322xp33_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_190),
.A3(n_195),
.B1(n_205),
.B2(n_213),
.C1(n_199),
.C2(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_199),
.B(n_164),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_206),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_170),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_194),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_240),
.B(n_242),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_182),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_265),
.B(n_241),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_188),
.B1(n_197),
.B2(n_200),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_257),
.B1(n_259),
.B2(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_253),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_95),
.Y(n_283)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_93),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_188),
.B1(n_215),
.B2(n_152),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_207),
.B1(n_216),
.B2(n_210),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_218),
.C(n_227),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_212),
.B1(n_202),
.B2(n_195),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_238),
.A2(n_193),
.B1(n_202),
.B2(n_155),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_231),
.B1(n_174),
.B2(n_221),
.Y(n_276)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_221),
.A2(n_155),
.B(n_180),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_271),
.C(n_273),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_260),
.A2(n_187),
.B1(n_230),
.B2(n_237),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_272),
.B1(n_278),
.B2(n_256),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_222),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_248),
.C(n_254),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_237),
.B1(n_226),
.B2(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_240),
.C(n_217),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_280),
.B(n_265),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_239),
.C(n_235),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_276),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_239),
.C(n_242),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_232),
.B1(n_184),
.B2(n_229),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_232),
.B(n_81),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_50),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_143),
.C(n_95),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_264),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_255),
.B1(n_244),
.B2(n_247),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_249),
.B1(n_257),
.B2(n_247),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_255),
.B1(n_251),
.B2(n_245),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_245),
.B(n_250),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_277),
.C(n_275),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_7),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_10),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_7),
.B(n_9),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_16),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_266),
.B(n_271),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_303),
.B(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_286),
.C(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_304),
.C(n_285),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_307),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_273),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_270),
.C(n_11),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_10),
.B(n_13),
.Y(n_306)
);

OAI221xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_316),
.Y(n_318)
);

OAI221xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_294),
.B1(n_295),
.B2(n_290),
.C(n_297),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_15),
.B(n_16),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_297),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_309),
.B(n_311),
.C(n_301),
.D(n_304),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_317),
.B(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_14),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_15),
.B(n_16),
.C(n_319),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_318),
.C(n_322),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_325),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_326),
.B(n_320),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_327),
.Y(n_330)
);


endmodule