module fake_jpeg_30002_n_399 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_399);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_399;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_332;
wire n_92;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_66),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_35),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_76),
.Y(n_105)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_32),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_25),
.B1(n_23),
.B2(n_39),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_86),
.A2(n_36),
.B1(n_26),
.B2(n_37),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_90),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_96),
.Y(n_135)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_41),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_110),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_41),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_61),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_119),
.Y(n_149)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_49),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_35),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_27),
.A3(n_24),
.B1(n_43),
.B2(n_33),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_76),
.C(n_39),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_138),
.B(n_147),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_34),
.B(n_50),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_145),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_71),
.B1(n_69),
.B2(n_83),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_154),
.B1(n_149),
.B2(n_109),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_48),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_48),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_98),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_94),
.A2(n_62),
.B1(n_58),
.B2(n_56),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_27),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_94),
.A2(n_53),
.B1(n_39),
.B2(n_50),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_86),
.B1(n_119),
.B2(n_108),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_43),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_105),
.B1(n_124),
.B2(n_106),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_172),
.B1(n_177),
.B2(n_181),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_107),
.B1(n_101),
.B2(n_115),
.Y(n_171)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_116),
.B(n_31),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_179),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_100),
.B1(n_118),
.B2(n_120),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_128),
.B1(n_125),
.B2(n_108),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_133),
.A2(n_100),
.B1(n_97),
.B2(n_120),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_146),
.Y(n_198)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_118),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_191),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_131),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_199),
.Y(n_208)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_139),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_200),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_134),
.Y(n_200)
);

INVx6_ASAP7_75t_SL g201 ( 
.A(n_170),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_169),
.B(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_204),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_150),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_168),
.Y(n_214)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_167),
.B1(n_164),
.B2(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_216),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_179),
.C(n_164),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_211),
.C(n_219),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_203),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_221),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_176),
.C(n_182),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_180),
.B(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_212),
.B(n_222),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_181),
.B(n_149),
.Y(n_215)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_177),
.B1(n_184),
.B2(n_168),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_222),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_160),
.B1(n_149),
.B2(n_174),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_194),
.B1(n_190),
.B2(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_150),
.C(n_166),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_136),
.B(n_130),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_194),
.B1(n_188),
.B2(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_247),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_206),
.C(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_236),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_198),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_229),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_215),
.B1(n_218),
.B2(n_220),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_189),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_242),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_230),
.B(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_197),
.C(n_191),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_187),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_197),
.C(n_191),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_220),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_187),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_210),
.B1(n_216),
.B2(n_201),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_225),
.B1(n_247),
.B2(n_230),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_241),
.B1(n_240),
.B2(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_243),
.B(n_202),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_262),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_193),
.B(n_212),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_188),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_213),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_226),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_211),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_219),
.B(n_188),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_155),
.Y(n_294)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_271),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_SL g276 ( 
.A(n_253),
.B(n_230),
.C(n_226),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_276),
.B(n_264),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_293),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_244),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_279),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_231),
.B1(n_244),
.B2(n_188),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_292),
.B1(n_255),
.B2(n_252),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_240),
.B1(n_196),
.B2(n_234),
.Y(n_284)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_259),
.B(n_201),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_287),
.B(n_294),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_170),
.C(n_173),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_295),
.C(n_278),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_141),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_260),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_256),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_262),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_209),
.B1(n_190),
.B2(n_136),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_141),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_173),
.C(n_166),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_298),
.A2(n_275),
.B1(n_285),
.B2(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_304),
.Y(n_328)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_279),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_306),
.Y(n_319)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_263),
.C(n_252),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_266),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_314),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_261),
.C(n_257),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_311),
.C(n_282),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_257),
.C(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_290),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_313),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_289),
.Y(n_314)
);

NOR4xp25_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_317),
.C(n_22),
.D(n_20),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_249),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_320),
.A2(n_325),
.B1(n_329),
.B2(n_296),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_276),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_324),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_283),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_286),
.B1(n_249),
.B2(n_277),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_142),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_303),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_327),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_297),
.A2(n_251),
.B1(n_292),
.B2(n_209),
.Y(n_329)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_310),
.C(n_311),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_336),
.C(n_318),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_309),
.A2(n_297),
.B(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_251),
.C(n_162),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_337),
.B(n_341),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_347),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_302),
.B1(n_300),
.B2(n_18),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_342),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_300),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_162),
.C(n_130),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_37),
.Y(n_344)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_20),
.B1(n_142),
.B2(n_153),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_349),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_129),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_129),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_350),
.B(n_336),
.C(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_353),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_348),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_322),
.C(n_324),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_354),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_328),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_358),
.B(n_340),
.Y(n_366)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_337),
.A2(n_327),
.B(n_334),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_155),
.Y(n_368)
);

OAI31xp33_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_340),
.A3(n_347),
.B(n_334),
.Y(n_365)
);

AOI322xp5_ASAP7_75t_L g379 ( 
.A1(n_365),
.A2(n_370),
.A3(n_371),
.B1(n_372),
.B2(n_42),
.C1(n_31),
.C2(n_26),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_366),
.B(n_369),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_105),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_128),
.C(n_92),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_374),
.Y(n_378)
);

AOI211xp5_ASAP7_75t_L g370 ( 
.A1(n_359),
.A2(n_49),
.B(n_44),
.C(n_40),
.Y(n_370)
);

OA21x2_ASAP7_75t_SL g371 ( 
.A1(n_362),
.A2(n_155),
.B(n_79),
.Y(n_371)
);

AOI31xp67_ASAP7_75t_L g372 ( 
.A1(n_355),
.A2(n_360),
.A3(n_351),
.B(n_44),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_155),
.B(n_40),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_3),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_88),
.C(n_91),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_382),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_377),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_32),
.C(n_42),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_379),
.A2(n_380),
.B(n_4),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_363),
.A2(n_1),
.B(n_2),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_2),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_378),
.B(n_5),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_3),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_383),
.B(n_3),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_365),
.C(n_123),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_386),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_4),
.C(n_5),
.Y(n_390)
);

AOI322xp5_ASAP7_75t_L g393 ( 
.A1(n_388),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_13),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_393),
.C(n_384),
.Y(n_395)
);

AOI322xp5_ASAP7_75t_L g392 ( 
.A1(n_389),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_392),
.Y(n_394)
);

AO221x1_ASAP7_75t_L g396 ( 
.A1(n_395),
.A2(n_391),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_394),
.B(n_15),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_6),
.C(n_15),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_17),
.Y(n_399)
);


endmodule