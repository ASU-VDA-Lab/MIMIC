module fake_jpeg_3603_n_226 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_11),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_96),
.Y(n_120)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_56),
.B1(n_54),
.B2(n_65),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_99),
.B1(n_71),
.B2(n_58),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_56),
.B1(n_74),
.B2(n_68),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_75),
.B1(n_67),
.B2(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_65),
.B1(n_60),
.B2(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_113),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_112),
.Y(n_133)
);

OR2x2_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_79),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_119),
.B(n_98),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_81),
.B1(n_73),
.B2(n_71),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_69),
.B1(n_63),
.B2(n_55),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_98),
.B1(n_70),
.B2(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_59),
.Y(n_113)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_117),
.Y(n_134)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_97),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_73),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_141),
.B1(n_7),
.B2(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_137),
.Y(n_151)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_5),
.Y(n_149)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_139),
.B1(n_127),
.B2(n_134),
.Y(n_153)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_68),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_1),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_30),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_55),
.B1(n_25),
.B2(n_26),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_23),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_33),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_141)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_147),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_115),
.B(n_111),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_150),
.B(n_16),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_115),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_36),
.C(n_44),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_51),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_2),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_153),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_5),
.B(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_6),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_160),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_29),
.B1(n_49),
.B2(n_48),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_162),
.B1(n_13),
.B2(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_7),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_12),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_32),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_16),
.B(n_17),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_170),
.Y(n_195)
);

NAND2xp67_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_136),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_149),
.B(n_150),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_131),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_176),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_35),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_147),
.C(n_159),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_183)
);

OAI22x1_ASAP7_75t_SL g194 ( 
.A1(n_183),
.A2(n_162),
.B1(n_18),
.B2(n_28),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_193),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_168),
.B1(n_173),
.B2(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_201),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_210)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_190),
.B(n_175),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_176),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_183),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_172),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_196),
.B1(n_169),
.B2(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_211),
.A2(n_213),
.B1(n_214),
.B2(n_180),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_196),
.B(n_144),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_198),
.B(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_191),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_219),
.B1(n_210),
.B2(n_202),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_188),
.C(n_212),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_183),
.A3(n_194),
.B1(n_157),
.B2(n_186),
.C1(n_182),
.C2(n_50),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_21),
.C(n_31),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_170),
.Y(n_226)
);


endmodule