module real_jpeg_4238_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_0),
.A2(n_151),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_0),
.A2(n_190),
.B1(n_197),
.B2(n_219),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_0),
.A2(n_219),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_0),
.A2(n_40),
.B1(n_59),
.B2(n_219),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_47),
.B1(n_70),
.B2(n_74),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_1),
.A2(n_74),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_1),
.A2(n_74),
.B1(n_177),
.B2(n_398),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_1),
.A2(n_74),
.B1(n_114),
.B2(n_412),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_54),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_54),
.B1(n_113),
.B2(n_117),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_2),
.A2(n_54),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_2),
.A2(n_54),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_46),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_60),
.B1(n_107),
.B2(n_110),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_3),
.A2(n_60),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_3),
.A2(n_60),
.B1(n_291),
.B2(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_176),
.B1(n_210),
.B2(n_214),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_4),
.A2(n_109),
.B1(n_118),
.B2(n_176),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_4),
.A2(n_51),
.B1(n_176),
.B2(n_348),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_5),
.Y(n_232)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_5),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_5),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_5),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_6),
.Y(n_342)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_6),
.Y(n_349)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_7),
.Y(n_345)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_8),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_9),
.Y(n_545)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_12),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_14),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_14),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_14),
.A2(n_80),
.B1(n_356),
.B2(n_360),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_14),
.A2(n_80),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_14),
.A2(n_80),
.B1(n_314),
.B2(n_451),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_15),
.A2(n_190),
.B1(n_196),
.B2(n_197),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_15),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_15),
.A2(n_148),
.B1(n_196),
.B2(n_259),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_15),
.A2(n_196),
.B1(n_346),
.B2(n_375),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_15),
.A2(n_196),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_17),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_17),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_17),
.B(n_185),
.C(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_17),
.B(n_97),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_17),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_17),
.B(n_146),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_17),
.B(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_18),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_18),
.A2(n_177),
.B1(n_283),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_18),
.A2(n_283),
.B1(n_289),
.B2(n_407),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_L g464 ( 
.A1(n_18),
.A2(n_283),
.B1(n_342),
.B2(n_465),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_540),
.B(n_542),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_55),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_24),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_24),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_25),
.B(n_171),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_25),
.A2(n_56),
.B1(n_414),
.B2(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_29),
.Y(n_290)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_30),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_30),
.Y(n_376)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_32),
.Y(n_340)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_34),
.A2(n_337),
.A3(n_341),
.B1(n_343),
.B2(n_347),
.Y(n_336)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_36),
.A2(n_368),
.B(n_369),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_36),
.B(n_371),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_37)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_40),
.Y(n_415)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_41),
.Y(n_465)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_53),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_55),
.B(n_65),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_61),
.B1(n_69),
.B2(n_75),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_75),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_56),
.A2(n_370),
.B(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_56),
.A2(n_61),
.B1(n_69),
.B2(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_61),
.A2(n_439),
.B(n_466),
.Y(n_476)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_157),
.B(n_539),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_153),
.C(n_154),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_66),
.A2(n_67),
.B1(n_535),
.B2(n_536),
.Y(n_534)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_81),
.C(n_119),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_68),
.B(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_81),
.A2(n_119),
.B1(n_120),
.B2(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_81),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_81)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_82),
.A2(n_111),
.B1(n_311),
.B2(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_82),
.A2(n_111),
.B1(n_406),
.B2(n_411),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_82),
.A2(n_106),
.B1(n_111),
.B2(n_516),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_97),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_91),
.B2(n_96),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_85),
.Y(n_296)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_86),
.Y(n_300)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_90),
.Y(n_274)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_90),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_90),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_97),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

AOI22x1_ASAP7_75t_L g440 ( 
.A1(n_97),
.A2(n_155),
.B1(n_317),
.B2(n_441),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_97),
.A2(n_155),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_105),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_101),
.Y(n_403)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_103),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_103),
.Y(n_398)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_104),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_104),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_111),
.B(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_111),
.A2(n_311),
.B(n_316),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_119),
.A2(n_120),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_119),
.B(n_511),
.C(n_514),
.Y(n_522)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_145),
.B(n_147),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_167),
.B(n_172),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_121),
.A2(n_145),
.B1(n_218),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_121),
.A2(n_172),
.B(n_258),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_121),
.A2(n_145),
.B1(n_378),
.B2(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_122),
.B(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_122),
.A2(n_146),
.B1(n_397),
.B2(n_399),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_122),
.A2(n_146),
.B1(n_399),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_122),
.A2(n_146),
.B1(n_421),
.B2(n_455),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_135),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_126),
.Y(n_424)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_135),
.A2(n_218),
.B(n_222),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_141),
.B2(n_143),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_140),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_140),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_141),
.Y(n_325)
);

BUFx8_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_142),
.Y(n_282)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_142),
.Y(n_359)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_145),
.A2(n_222),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_147),
.Y(n_455)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g297 ( 
.A(n_150),
.B(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_153),
.B(n_154),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_155),
.A2(n_266),
.B(n_275),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_155),
.B(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_155),
.A2(n_275),
.B(n_479),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_533),
.B(n_538),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_505),
.B(n_530),
.Y(n_158)
);

OAI311xp33_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_383),
.A3(n_481),
.B1(n_499),
.C1(n_504),
.Y(n_159)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_330),
.B(n_382),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_302),
.B(n_329),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_252),
.B(n_301),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_225),
.B(n_251),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_187),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_165),
.B(n_187),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_180),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_166),
.A2(n_180),
.B1(n_181),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_200),
.B(n_206),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g266 ( 
.A1(n_171),
.A2(n_267),
.B(n_271),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_171),
.B(n_348),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_171),
.A2(n_347),
.B(n_348),
.Y(n_368)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_215),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_188),
.B(n_216),
.C(n_224),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_200),
.B(n_206),
.Y(n_188)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_195),
.Y(n_324)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_199),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_200),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_200),
.A2(n_353),
.B1(n_389),
.B2(n_392),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_200),
.A2(n_392),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_209),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_201),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_201),
.A2(n_280),
.B1(n_321),
.B2(n_326),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_201),
.A2(n_355),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_207),
.Y(n_353)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_223),
.B2(n_224),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_241),
.B(n_250),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_240),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_239),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B(n_238),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_279),
.B(n_285),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_248),
.Y(n_250)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_254),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_277),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_264),
.B2(n_265),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_264),
.C(n_277),
.Y(n_303)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_267),
.Y(n_412)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_270),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_289),
.A3(n_291),
.B1(n_294),
.B2(n_297),
.Y(n_288)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_288),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_288),
.Y(n_308)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_304),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_328),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_308),
.C(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_318),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_319),
.C(n_320),
.Y(n_362)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_324),
.Y(n_361)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_331),
.B(n_332),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_365),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_333)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_350),
.B2(n_351),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_336),
.B(n_350),
.Y(n_477)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_362),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_362),
.B(n_363),
.C(n_365),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_372),
.B2(n_381),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_366),
.B(n_373),
.C(n_377),
.Y(n_490)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_377),
.Y(n_372)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_374),
.Y(n_479)
);

INVx6_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_467),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_SL g499 ( 
.A1(n_384),
.A2(n_467),
.B(n_500),
.C(n_503),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_442),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_385),
.B(n_442),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_418),
.C(n_430),
.Y(n_385)
);

FAx1_ASAP7_75t_SL g480 ( 
.A(n_386),
.B(n_418),
.CI(n_430),
.CON(n_480),
.SN(n_480)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_404),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_387),
.B(n_405),
.C(n_413),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_396),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_388),
.B(n_396),
.Y(n_473)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_389),
.Y(n_435)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_413),
.Y(n_404)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_406),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_425),
.B2(n_429),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_425),
.Y(n_459)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_425),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_425),
.A2(n_429),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_425),
.A2(n_459),
.B(n_462),
.Y(n_508)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_428),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_437),
.C(n_440),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_432),
.B(n_434),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_437),
.A2(n_438),
.B1(n_440),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_446),
.C(n_457),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_457),
.B2(n_458),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_453),
.B(n_456),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_454),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

FAx1_ASAP7_75t_SL g507 ( 
.A(n_456),
.B(n_508),
.CI(n_509),
.CON(n_507),
.SN(n_507)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_456),
.B(n_508),
.C(n_509),
.Y(n_529)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_480),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_468),
.B(n_480),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_473),
.C(n_474),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_469),
.A2(n_470),
.B1(n_473),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_492),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.C(n_478),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_475),
.A2(n_476),
.B1(n_478),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_478),
.Y(n_487)
);

BUFx24_ASAP7_75t_SL g547 ( 
.A(n_480),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_494),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_483),
.A2(n_501),
.B(n_502),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_491),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_491),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_488),
.C(n_490),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_497),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_488),
.A2(n_489),
.B1(n_490),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_496),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_519),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_518),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_518),
.Y(n_531)
);

BUFx24_ASAP7_75t_SL g548 ( 
.A(n_507),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_513),
.B2(n_517),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_510),
.A2(n_511),
.B1(n_525),
.B2(n_526),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_510),
.B(n_521),
.C(n_525),
.Y(n_537)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_513),
.Y(n_517)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_531),
.B(n_532),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_520),
.B(n_529),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_529),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_522),
.B1(n_523),
.B2(n_524),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_537),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_534),
.B(n_537),
.Y(n_538)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx8_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx13_ASAP7_75t_L g544 ( 
.A(n_541),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_545),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);


endmodule