module fake_jpeg_28648_n_484 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_484);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_484;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_63),
.Y(n_100)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_51),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_20),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_25),
.B1(n_47),
.B2(n_46),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_69),
.Y(n_105)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_73),
.Y(n_121)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_16),
.B(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_78),
.B(n_84),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_88),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_4),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_87),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_4),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_92),
.B(n_52),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_10),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_40),
.B1(n_20),
.B2(n_36),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_99),
.A2(n_107),
.B1(n_112),
.B2(n_115),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_40),
.B1(n_36),
.B2(n_49),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_63),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_43),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_114),
.A2(n_124),
.B1(n_136),
.B2(n_41),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_53),
.A2(n_40),
.B1(n_49),
.B2(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_25),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_126),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_49),
.B1(n_33),
.B2(n_29),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_120),
.A2(n_132),
.B1(n_54),
.B2(n_61),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_56),
.B1(n_83),
.B2(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_30),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_65),
.A2(n_33),
.B1(n_47),
.B2(n_30),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_134),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_60),
.A2(n_27),
.B1(n_46),
.B2(n_44),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_70),
.A2(n_27),
.B1(n_46),
.B2(n_44),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_30),
.B1(n_47),
.B2(n_44),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_52),
.Y(n_156)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_154),
.Y(n_204)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_158),
.Y(n_220)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_159),
.B(n_160),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_74),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_74),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_163),
.Y(n_210)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_164),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_122),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_178),
.Y(n_216)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_168),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_186),
.Y(n_217)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g175 ( 
.A(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_184),
.B1(n_193),
.B2(n_195),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_51),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_102),
.A2(n_97),
.B1(n_77),
.B2(n_72),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_191),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_55),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_55),
.B(n_106),
.C(n_143),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_179),
.B(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_138),
.A2(n_66),
.B1(n_62),
.B2(n_96),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_192),
.B1(n_198),
.B2(n_41),
.Y(n_207)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_86),
.A3(n_89),
.B1(n_27),
.B2(n_43),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_42),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_188),
.Y(n_235)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_123),
.A2(n_95),
.B1(n_43),
.B2(n_42),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_196),
.Y(n_211)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_118),
.B(n_42),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_41),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_152),
.Y(n_229)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_98),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_110),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_109),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_147),
.B1(n_117),
.B2(n_103),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_206),
.A2(n_214),
.B(n_189),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_207),
.A2(n_191),
.B1(n_172),
.B2(n_182),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_143),
.B1(n_106),
.B2(n_137),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_213),
.A2(n_239),
.B1(n_244),
.B2(n_175),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_152),
.B(n_128),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_148),
.A3(n_35),
.B1(n_34),
.B2(n_24),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_229),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_170),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_35),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_165),
.B(n_35),
.C(n_34),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_227),
.C(n_232),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_104),
.C(n_130),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_186),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_153),
.B(n_103),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_178),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_113),
.B1(n_137),
.B2(n_135),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_181),
.A2(n_135),
.B1(n_113),
.B2(n_145),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_177),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_253),
.A2(n_212),
.B1(n_231),
.B2(n_230),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_163),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_256),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_146),
.B1(n_173),
.B2(n_155),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_259),
.B1(n_265),
.B2(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_207),
.B1(n_217),
.B2(n_214),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_157),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_261),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_164),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_159),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_222),
.B1(n_208),
.B2(n_216),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_269),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_268),
.A2(n_223),
.B(n_224),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_270),
.A2(n_277),
.B1(n_283),
.B2(n_231),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_211),
.B(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_275),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_167),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_225),
.C(n_209),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_210),
.B(n_34),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_209),
.C(n_242),
.Y(n_296)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_220),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_146),
.B1(n_193),
.B2(n_190),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_211),
.B(n_229),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_204),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_240),
.A2(n_171),
.B1(n_147),
.B2(n_154),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_224),
.B(n_204),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_216),
.A2(n_166),
.B1(n_127),
.B2(n_130),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_175),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_212),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_219),
.A2(n_127),
.B1(n_203),
.B2(n_200),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_300),
.C(n_301),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_291),
.B(n_312),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_259),
.A2(n_257),
.B1(n_250),
.B2(n_275),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_293),
.A2(n_309),
.B1(n_277),
.B2(n_288),
.Y(n_331)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_260),
.A2(n_254),
.B(n_274),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_296),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_298),
.B(n_183),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_215),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_299),
.B(n_311),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_255),
.C(n_261),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_245),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_242),
.B(n_245),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_304),
.A2(n_318),
.B(n_282),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_305),
.A2(n_315),
.B1(n_253),
.B2(n_281),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_272),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_307),
.B(n_266),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_243),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_252),
.A2(n_218),
.B(n_234),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_276),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_226),
.B1(n_231),
.B2(n_218),
.Y(n_315)
);

OR2x6_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_183),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_316),
.A2(n_267),
.B(n_234),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_265),
.A2(n_250),
.B(n_280),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_321),
.B(n_322),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_271),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_323),
.A2(n_342),
.B(n_317),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_256),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_324),
.B(n_327),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_334),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_287),
.B(n_286),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_264),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_330),
.C(n_336),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_249),
.Y(n_329)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_251),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_331),
.A2(n_289),
.B1(n_297),
.B2(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_248),
.C(n_247),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_263),
.C(n_258),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_320),
.C(n_322),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_318),
.B(n_297),
.Y(n_342)
);

AND2x2_ASAP7_75t_SL g343 ( 
.A(n_316),
.B(n_243),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_343),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_283),
.Y(n_344)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_345),
.B(n_348),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_347),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_303),
.B(n_194),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_230),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_350),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_351),
.A2(n_290),
.B1(n_292),
.B2(n_294),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_347),
.A2(n_305),
.B1(n_287),
.B2(n_315),
.Y(n_357)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_358),
.A2(n_377),
.B1(n_350),
.B2(n_343),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_340),
.A2(n_316),
.B1(n_293),
.B2(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_364),
.C(n_369),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_288),
.C(n_304),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g366 ( 
.A1(n_346),
.A2(n_316),
.B1(n_291),
.B2(n_294),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_10),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_332),
.A2(n_337),
.B(n_343),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_368),
.A2(n_128),
.B(n_1),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_312),
.C(n_314),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_292),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_10),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_341),
.C(n_336),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_372),
.C(n_338),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_317),
.C(n_314),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_375),
.A2(n_332),
.B(n_334),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_331),
.A2(n_344),
.B1(n_342),
.B2(n_333),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_380),
.A2(n_402),
.B(n_353),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_394),
.B1(n_352),
.B2(n_354),
.Y(n_417)
);

A2O1A1O1Ixp25_ASAP7_75t_L g383 ( 
.A1(n_375),
.A2(n_326),
.B(n_335),
.C(n_329),
.D(n_349),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_400),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_363),
.B(n_327),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_384),
.B(n_388),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_335),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_365),
.Y(n_407)
);

FAx1_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_324),
.CI(n_325),
.CON(n_386),
.SN(n_386)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_363),
.B(n_351),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_339),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_393),
.C(n_370),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_226),
.C(n_195),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_377),
.A2(n_202),
.B1(n_162),
.B2(n_169),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_395),
.A2(n_373),
.B(n_402),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_379),
.A2(n_183),
.B1(n_24),
.B2(n_0),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_397),
.A2(n_356),
.B1(n_355),
.B2(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_398),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_374),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_399)
);

AOI322xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_354),
.A3(n_355),
.B1(n_356),
.B2(n_353),
.C1(n_379),
.C2(n_358),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_372),
.Y(n_411)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_1),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_369),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_397),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_405),
.B(n_420),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_373),
.B(n_368),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_406),
.A2(n_395),
.B(n_391),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_419),
.Y(n_429)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_408),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_400),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_371),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_421),
.Y(n_426)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_396),
.B1(n_394),
.B2(n_393),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_359),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_366),
.B(n_359),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_437),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g424 ( 
.A(n_410),
.B(n_382),
.CI(n_386),
.CON(n_424),
.SN(n_424)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_430),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_409),
.A2(n_401),
.B(n_383),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_425),
.A2(n_433),
.B(n_424),
.Y(n_450)
);

OAI221xp5_ASAP7_75t_L g427 ( 
.A1(n_416),
.A2(n_392),
.B1(n_389),
.B2(n_403),
.C(n_387),
.Y(n_427)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_406),
.A2(n_366),
.B(n_386),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_428),
.B(n_408),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_435),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_366),
.B1(n_2),
.B2(n_3),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_3),
.Y(n_437)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_438),
.Y(n_439)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_410),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_446),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_443),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_420),
.C(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_445),
.B(n_447),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_R g446 ( 
.A(n_424),
.B(n_422),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_414),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_414),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_11),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_452),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_438),
.A2(n_404),
.B1(n_417),
.B2(n_419),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_433),
.C(n_431),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

AO22x1_ASAP7_75t_L g454 ( 
.A1(n_450),
.A2(n_428),
.B1(n_423),
.B2(n_431),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_460),
.C(n_442),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_460),
.C(n_453),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_440),
.A2(n_412),
.B(n_432),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_458),
.B(n_459),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_429),
.C(n_407),
.Y(n_459)
);

AOI21x1_ASAP7_75t_SL g460 ( 
.A1(n_444),
.A2(n_413),
.B(n_429),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_461),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_449),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_466),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

AO21x1_ASAP7_75t_L g475 ( 
.A1(n_467),
.A2(n_470),
.B(n_11),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_452),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_471),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_456),
.B(n_11),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_469),
.A2(n_12),
.B(n_15),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_467),
.A2(n_454),
.B1(n_453),
.B2(n_12),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_474),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_475),
.A2(n_15),
.B(n_0),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_476),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_479),
.A2(n_472),
.B(n_473),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_477),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g482 ( 
.A1(n_480),
.A2(n_481),
.B(n_465),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_482),
.A2(n_478),
.B(n_0),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_0),
.B(n_475),
.Y(n_484)
);


endmodule