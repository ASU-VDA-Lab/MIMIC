module fake_jpeg_23802_n_46 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx4_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_29),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_12),
.B1(n_18),
.B2(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_30),
.B1(n_19),
.B2(n_7),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_1),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_22),
.B1(n_24),
.B2(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_33),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_32),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_37),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_6),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_15),
.Y(n_46)
);


endmodule