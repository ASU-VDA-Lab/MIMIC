module real_jpeg_3469_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_57),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_24),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_4),
.A2(n_85),
.B(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_51),
.C(n_62),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_31),
.B1(n_33),
.B2(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_48),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_106),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_24),
.B(n_74),
.Y(n_168)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_31),
.B1(n_33),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_67),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_12),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_14),
.A2(n_35),
.B1(n_85),
.B2(n_86),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_19),
.B(n_80),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.C(n_71),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_20),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_21),
.B(n_39),
.C(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_22),
.A2(n_30),
.B1(n_34),
.B2(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_43),
.C(n_86),
.Y(n_120)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_25),
.B(n_29),
.C(n_33),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_44),
.B(n_89),
.C(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_31),
.B(n_73),
.C(n_75),
.Y(n_72)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_31),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_31),
.B(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_84),
.B1(n_91),
.B2(n_93),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_92),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_43),
.A2(n_44),
.B1(n_85),
.B2(n_86),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_55),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_47),
.B(n_78),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_47),
.A2(n_77),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_48),
.A2(n_58),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_58),
.B1(n_90),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_48),
.A2(n_58),
.B1(n_149),
.B2(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_51),
.B(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_58),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_71),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_60),
.A2(n_106),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_60),
.A2(n_106),
.B1(n_134),
.B2(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_66),
.A2(n_103),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_72),
.B(n_76),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_107),
.B2(n_108),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_94),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_90),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_173),
.B(n_177),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_162),
.B(n_172),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_143),
.B(n_161),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_140),
.C(n_142),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_155),
.B(n_160),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_150),
.B(n_154),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_153),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_159),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_176),
.Y(n_177)
);


endmodule