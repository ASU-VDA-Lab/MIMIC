module fake_jpeg_14990_n_349 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_48),
.Y(n_63)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_24),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_36),
.B1(n_24),
.B2(n_34),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_74),
.Y(n_94)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_34),
.B1(n_46),
.B2(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_45),
.B1(n_36),
.B2(n_18),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_81),
.B1(n_84),
.B2(n_91),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_39),
.C(n_47),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_85),
.C(n_52),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_45),
.B1(n_32),
.B2(n_26),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_39),
.C(n_47),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_99),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_46),
.B1(n_34),
.B2(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_50),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_104),
.Y(n_120)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_50),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_31),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_25),
.B1(n_35),
.B2(n_33),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_30),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_50),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_31),
.C(n_20),
.Y(n_163)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_133),
.B1(n_137),
.B2(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_67),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_35),
.B(n_25),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_62),
.Y(n_130)
);

FAx1_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_58),
.CI(n_77),
.CON(n_131),
.SN(n_131)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_27),
.A3(n_21),
.B1(n_22),
.B2(n_28),
.Y(n_156)
);

NOR2xp67_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_82),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_0),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_56),
.C(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_23),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_25),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_135),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_0),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_29),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_29),
.B1(n_33),
.B2(n_86),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_140),
.B(n_28),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_93),
.B1(n_54),
.B2(n_88),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_149),
.B1(n_162),
.B2(n_133),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_156),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_136),
.B1(n_88),
.B2(n_115),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_152),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_86),
.B1(n_56),
.B2(n_99),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_105),
.B(n_73),
.C(n_69),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_133),
.B(n_129),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_92),
.B1(n_91),
.B2(n_105),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_92),
.B1(n_29),
.B2(n_20),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_86),
.B1(n_73),
.B2(n_52),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_134),
.C(n_120),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_128),
.B1(n_124),
.B2(n_130),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_126),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_162),
.Y(n_165)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_173),
.B1(n_178),
.B2(n_184),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_109),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_171),
.C(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_174),
.B(n_176),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_163),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_172),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_114),
.B1(n_110),
.B2(n_113),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_185),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_125),
.B(n_123),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_95),
.C(n_118),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_112),
.B(n_111),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_31),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_148),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_117),
.B(n_105),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_147),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_147),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_206),
.B(n_210),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_171),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_184),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_147),
.B1(n_141),
.B2(n_158),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_186),
.B1(n_173),
.B2(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_217),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_190),
.B1(n_166),
.B2(n_189),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_164),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_211),
.C(n_28),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_150),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_154),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_154),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_214),
.B(n_218),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_142),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_142),
.C(n_13),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_196),
.B1(n_192),
.B2(n_198),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_223),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_188),
.C(n_181),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_174),
.B1(n_167),
.B2(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_235),
.B1(n_238),
.B2(n_240),
.Y(n_257)
);

XOR2x2_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_176),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_229),
.A2(n_241),
.B(n_23),
.Y(n_261)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_193),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_95),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_201),
.C(n_202),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_212),
.B(n_31),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_205),
.A2(n_28),
.B(n_27),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_228),
.Y(n_266)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_246),
.B(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_192),
.B1(n_204),
.B2(n_197),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_254),
.B1(n_259),
.B2(n_266),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_201),
.B1(n_197),
.B2(n_210),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_222),
.C(n_242),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_228),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_195),
.B1(n_215),
.B2(n_1),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_219),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_207),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_235),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_246),
.B(n_223),
.CI(n_232),
.CON(n_274),
.SN(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_236),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_275),
.B(n_277),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_239),
.B(n_5),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_261),
.B(n_5),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_27),
.C(n_22),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_258),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_22),
.C(n_21),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_248),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_247),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_21),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_20),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_283),
.A2(n_264),
.B(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_277),
.Y(n_306)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_268),
.A2(n_253),
.B1(n_250),
.B2(n_257),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_274),
.B1(n_285),
.B2(n_4),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_R g297 ( 
.A(n_284),
.B(n_248),
.C(n_245),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_11),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_294),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_251),
.B(n_5),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_300),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_271),
.A2(n_251),
.B(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_270),
.B1(n_284),
.B2(n_269),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_20),
.C(n_4),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_290),
.C(n_292),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_287),
.B(n_17),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_11),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_314),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_299),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_12),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_295),
.B(n_11),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_10),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_313),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_304),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_301),
.C(n_290),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_325),
.C(n_309),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_SL g335 ( 
.A(n_326),
.B(n_8),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_4),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_9),
.C(n_12),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_303),
.B1(n_308),
.B2(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_331),
.A2(n_332),
.B(n_333),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_298),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_321),
.A2(n_10),
.B(n_7),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_318),
.B(n_9),
.Y(n_338)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_319),
.B(n_317),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_337),
.A2(n_329),
.B(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_340),
.C(n_9),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_330),
.A2(n_320),
.B(n_323),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_13),
.B(n_14),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_342),
.Y(n_345)
);

O2A1O1Ixp33_ASAP7_75t_SL g346 ( 
.A1(n_345),
.A2(n_344),
.B(n_336),
.C(n_341),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_343),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_14),
.C(n_16),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_4),
.Y(n_349)
);


endmodule