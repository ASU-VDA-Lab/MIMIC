module fake_jpeg_15712_n_38 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_21),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_1),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_16),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_21),
.B(n_14),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_15),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_15),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_30),
.B(n_29),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_23),
.B(n_7),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_18),
.C(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_1),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_35),
.C2(n_29),
.Y(n_38)
);


endmodule