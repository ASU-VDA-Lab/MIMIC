module fake_jpeg_13158_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_62),
.Y(n_70)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_40),
.B1(n_52),
.B2(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_22),
.Y(n_93)
);

AOI22x1_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_54),
.B1(n_42),
.B2(n_47),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_59),
.B1(n_57),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_48),
.B1(n_41),
.B2(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_1),
.Y(n_79)
);

FAx1_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_0),
.CI(n_1),
.CON(n_78),
.SN(n_78)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_2),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_91),
.B1(n_20),
.B2(n_9),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_85),
.Y(n_105)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_3),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_3),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_88),
.B(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_4),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_93),
.B(n_27),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_37),
.Y(n_115)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_30),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_97),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_32),
.Y(n_113)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_34),
.B(n_36),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_123),
.B(n_118),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_121),
.A3(n_105),
.B1(n_115),
.B2(n_112),
.C1(n_95),
.C2(n_108),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_113),
.Y(n_129)
);


endmodule