module fake_netlist_5_270_n_1027 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1027);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1027;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_607;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_699;
wire n_632;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_49),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_82),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_127),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_45),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_117),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_29),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_148),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_77),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_69),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_132),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_213),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_101),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_86),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_115),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_30),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_114),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_196),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_56),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_32),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_120),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_68),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_40),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_3),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_9),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_152),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_16),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_150),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_143),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_121),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_119),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_6),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_60),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_75),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_79),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_102),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_100),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_178),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_164),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_85),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_171),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_61),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_149),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_36),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_70),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_95),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_74),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_38),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_23),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_138),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_34),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_20),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_11),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_26),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_108),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_103),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_39),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_124),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_97),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_163),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_36),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_99),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_57),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_33),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_71),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_35),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_184),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_105),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_187),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_123),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_176),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_153),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_31),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_32),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_47),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_225),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_0),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_232),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_265),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_258),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_234),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_247),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_247),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_0),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_237),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_290),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_290),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_261),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_253),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_223),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_239),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_248),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_241),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_242),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_258),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_245),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_229),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_235),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_249),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_265),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_252),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_251),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_318),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_240),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_281),
.B(n_1),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_275),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_259),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_281),
.B(n_2),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_260),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_275),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_264),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_228),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_233),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_270),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_292),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_256),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_297),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_236),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_238),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_285),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_338),
.A2(n_307),
.B1(n_308),
.B2(n_304),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_303),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_285),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_340),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_326),
.B(n_329),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_334),
.B(n_341),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_342),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_360),
.B(n_267),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_343),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_336),
.B(n_267),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_254),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_353),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_254),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_349),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_267),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_305),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_356),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_374),
.B(n_337),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_324),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_362),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_362),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_350),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_R g428 ( 
.A(n_369),
.B(n_230),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_R g429 ( 
.A(n_372),
.B(n_257),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_330),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_381),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_350),
.Y(n_437)
);

BUFx4f_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_317),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_380),
.A2(n_305),
.B1(n_243),
.B2(n_255),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_410),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_403),
.B(n_401),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_250),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_403),
.B(n_303),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_403),
.B(n_303),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_378),
.A2(n_272),
.B1(n_276),
.B2(n_244),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_230),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_231),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_435),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_429),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_380),
.A2(n_287),
.B1(n_288),
.B2(n_283),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_411),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_293),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_385),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_408),
.B(n_298),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_382),
.B(n_419),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_303),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

INVx4_ASAP7_75t_SL g478 ( 
.A(n_380),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_415),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_412),
.B(n_306),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_380),
.B(n_263),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_319),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_409),
.B(n_224),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_398),
.B(n_266),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_380),
.B(n_391),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_413),
.B(n_379),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_351),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_413),
.B(n_268),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_392),
.B(n_269),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_399),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_381),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_399),
.B(n_351),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_381),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_424),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_380),
.B(n_271),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_386),
.B(n_231),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_407),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

OAI221xp5_ASAP7_75t_L g508 ( 
.A1(n_400),
.A2(n_316),
.B1(n_315),
.B2(n_273),
.C(n_278),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_404),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_448),
.A2(n_279),
.B(n_274),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_448),
.B(n_465),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_434),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_486),
.A2(n_418),
.B1(n_423),
.B2(n_331),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_473),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_486),
.A2(n_289),
.B1(n_314),
.B2(n_311),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_460),
.B(n_388),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_457),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_483),
.A2(n_277),
.B1(n_312),
.B2(n_309),
.Y(n_521)
);

INVx8_ASAP7_75t_L g522 ( 
.A(n_480),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_280),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_474),
.A2(n_301),
.B1(n_284),
.B2(n_299),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_441),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_474),
.B(n_431),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_479),
.B(n_434),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_505),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_282),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_475),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_388),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_502),
.A2(n_348),
.B1(n_328),
.B2(n_435),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_397),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_505),
.B(n_302),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_507),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_313),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_460),
.B(n_397),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_472),
.B(n_315),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_501),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_472),
.B(n_483),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_468),
.B(n_432),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_434),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_483),
.B(n_316),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_506),
.B(n_277),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_480),
.A2(n_277),
.B1(n_309),
.B2(n_312),
.Y(n_547)
);

NOR2x1p5_ASAP7_75t_L g548 ( 
.A(n_509),
.B(n_430),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_506),
.B(n_309),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_506),
.B(n_312),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_458),
.B(n_433),
.C(n_432),
.Y(n_552)
);

A2O1A1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_458),
.A2(n_433),
.B(n_430),
.C(n_434),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_508),
.B(n_424),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_485),
.B(n_444),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_446),
.B(n_46),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_447),
.A2(n_434),
.B1(n_430),
.B2(n_425),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_422),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_438),
.A2(n_426),
.B(n_427),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_488),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_463),
.B(n_48),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_451),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_461),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_466),
.A2(n_469),
.B1(n_439),
.B2(n_484),
.Y(n_567)
);

AND2x6_ASAP7_75t_SL g568 ( 
.A(n_499),
.B(n_328),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_440),
.B(n_50),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_444),
.B(n_51),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_462),
.B(n_54),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_462),
.B(n_58),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_480),
.A2(n_427),
.B1(n_348),
.B2(n_425),
.Y(n_575)
);

O2A1O1Ixp5_ASAP7_75t_L g576 ( 
.A1(n_450),
.A2(n_128),
.B(n_222),
.C(n_221),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_L g577 ( 
.A(n_480),
.B(n_59),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_509),
.B(n_2),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_450),
.B(n_62),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_453),
.B(n_63),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_453),
.B(n_64),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_484),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_509),
.B(n_4),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_461),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_471),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_477),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_502),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_504),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_480),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_482),
.A2(n_492),
.B1(n_504),
.B2(n_481),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_471),
.B(n_65),
.Y(n_591)
);

NAND2x1p5_ASAP7_75t_L g592 ( 
.A(n_440),
.B(n_66),
.Y(n_592)
);

NAND2x1_ASAP7_75t_L g593 ( 
.A(n_436),
.B(n_67),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_510),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_487),
.B(n_72),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_445),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_482),
.A2(n_134),
.B1(n_220),
.B2(n_218),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_528),
.B(n_482),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_528),
.B(n_482),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_544),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_R g601 ( 
.A(n_587),
.B(n_511),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_513),
.A2(n_482),
.B1(n_492),
.B2(n_503),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_535),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_517),
.B(n_445),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_513),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_517),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_517),
.B(n_478),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_589),
.A2(n_455),
.B1(n_476),
.B2(n_487),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_530),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_596),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_568),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_544),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_560),
.Y(n_614)
);

BUFx4f_ASAP7_75t_L g615 ( 
.A(n_544),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_522),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_523),
.B(n_467),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_526),
.B(n_495),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_563),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_522),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_540),
.B(n_467),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_565),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_566),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_555),
.B(n_464),
.Y(n_627)
);

AO22x1_ASAP7_75t_L g628 ( 
.A1(n_554),
.A2(n_495),
.B1(n_459),
.B2(n_476),
.Y(n_628)
);

BUFx12f_ASAP7_75t_L g629 ( 
.A(n_548),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_550),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_520),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_582),
.A2(n_476),
.B1(n_498),
.B2(n_491),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_541),
.B(n_442),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_584),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_594),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_532),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_545),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_SL g638 ( 
.A(n_552),
.B(n_489),
.C(n_7),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_514),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_596),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_572),
.Y(n_641)
);

AND3x1_ASAP7_75t_SL g642 ( 
.A(n_543),
.B(n_8),
.C(n_9),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_539),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_542),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_561),
.B(n_464),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_SL g648 ( 
.A(n_553),
.B(n_533),
.C(n_531),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_558),
.B(n_442),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_562),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_586),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_572),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_577),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_519),
.B(n_442),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_546),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_591),
.Y(n_656)
);

AND2x2_ASAP7_75t_SL g657 ( 
.A(n_573),
.B(n_438),
.Y(n_657)
);

AND3x1_ASAP7_75t_L g658 ( 
.A(n_516),
.B(n_498),
.C(n_491),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_575),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_578),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_549),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_557),
.Y(n_662)
);

INVx3_ASAP7_75t_SL g663 ( 
.A(n_583),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_624),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_641),
.A2(n_590),
.B(n_534),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_605),
.B(n_567),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_654),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_627),
.A2(n_569),
.B(n_591),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_618),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_641),
.A2(n_529),
.B(n_579),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_579),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_648),
.B(n_524),
.C(n_521),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_661),
.B(n_538),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_615),
.Y(n_674)
);

AO31x2_ASAP7_75t_L g675 ( 
.A1(n_656),
.A2(n_580),
.A3(n_581),
.B(n_595),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_641),
.A2(n_581),
.B(n_580),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_603),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_656),
.B(n_556),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_660),
.A2(n_573),
.B(n_574),
.C(n_518),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_657),
.A2(n_571),
.B(n_576),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_657),
.A2(n_571),
.B(n_574),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_629),
.B(n_559),
.Y(n_682)
);

BUFx4_ASAP7_75t_SL g683 ( 
.A(n_651),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_598),
.A2(n_595),
.B(n_593),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_599),
.A2(n_592),
.B(n_564),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_647),
.A2(n_592),
.B(n_500),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_660),
.A2(n_536),
.B(n_547),
.C(n_512),
.Y(n_687)
);

AO31x2_ASAP7_75t_L g688 ( 
.A1(n_633),
.A2(n_551),
.A3(n_436),
.B(n_476),
.Y(n_688)
);

AOI21x1_ASAP7_75t_L g689 ( 
.A1(n_621),
.A2(n_527),
.B(n_436),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_651),
.B(n_537),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_606),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_610),
.B(n_452),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_633),
.B(n_452),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_641),
.A2(n_490),
.B(n_452),
.Y(n_694)
);

INVx6_ASAP7_75t_SL g695 ( 
.A(n_608),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_611),
.A2(n_500),
.B(n_597),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_650),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_611),
.A2(n_478),
.B(n_452),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_634),
.Y(n_699)
);

NOR2x1_ASAP7_75t_SL g700 ( 
.A(n_620),
.B(n_490),
.Y(n_700)
);

AOI21x1_ASAP7_75t_L g701 ( 
.A1(n_617),
.A2(n_478),
.B(n_490),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_640),
.A2(n_643),
.B(n_634),
.Y(n_702)
);

NOR2x1_ASAP7_75t_SL g703 ( 
.A(n_620),
.B(n_490),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_645),
.B(n_476),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_628),
.B(n_497),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_645),
.B(n_497),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_659),
.A2(n_497),
.B1(n_12),
.B2(n_13),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_640),
.A2(n_497),
.B(n_76),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_631),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_601),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_602),
.A2(n_137),
.B(n_216),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_653),
.A2(n_135),
.B(n_215),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_624),
.Y(n_714)
);

AO21x1_ASAP7_75t_L g715 ( 
.A1(n_622),
.A2(n_10),
.B(n_12),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_677),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_674),
.B(n_604),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_699),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_672),
.A2(n_659),
.B1(n_662),
.B2(n_669),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_702),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_691),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_706),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_697),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_683),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_669),
.B(n_638),
.Y(n_726)
);

OAI21x1_ASAP7_75t_SL g727 ( 
.A1(n_712),
.A2(n_622),
.B(n_632),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_667),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_695),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_692),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_698),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_695),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_712),
.A2(n_662),
.B1(n_663),
.B2(n_636),
.Y(n_733)
);

AO31x2_ASAP7_75t_L g734 ( 
.A1(n_679),
.A2(n_643),
.A3(n_619),
.B(n_625),
.Y(n_734)
);

OA21x2_ASAP7_75t_L g735 ( 
.A1(n_681),
.A2(n_632),
.B(n_609),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_686),
.A2(n_658),
.B(n_646),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_690),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_674),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_666),
.B(n_663),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_673),
.B(n_614),
.Y(n_740)
);

AOI21xp33_ASAP7_75t_SL g741 ( 
.A1(n_711),
.A2(n_636),
.B(n_635),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_709),
.A2(n_646),
.B(n_644),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_671),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_696),
.A2(n_644),
.B(n_623),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_684),
.A2(n_652),
.B(n_609),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_671),
.B(n_600),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_701),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_681),
.A2(n_653),
.B(n_615),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_685),
.A2(n_652),
.B(n_649),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_674),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_680),
.A2(n_653),
.B(n_604),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_687),
.A2(n_604),
.B(n_653),
.Y(n_752)
);

CKINVDCx11_ASAP7_75t_R g753 ( 
.A(n_664),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_678),
.B(n_639),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_690),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_714),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_708),
.A2(n_613),
.B1(n_600),
.B2(n_639),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_665),
.A2(n_620),
.B(n_626),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_670),
.A2(n_620),
.B(n_626),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_682),
.Y(n_760)
);

AO21x2_ASAP7_75t_L g761 ( 
.A1(n_680),
.A2(n_654),
.B(n_645),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_678),
.A2(n_626),
.B(n_608),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_675),
.Y(n_763)
);

AOI21x1_ASAP7_75t_L g764 ( 
.A1(n_689),
.A2(n_608),
.B(n_645),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_708),
.B(n_607),
.Y(n_765)
);

INVx6_ASAP7_75t_L g766 ( 
.A(n_682),
.Y(n_766)
);

AO21x1_ASAP7_75t_L g767 ( 
.A1(n_693),
.A2(n_642),
.B(n_607),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_733),
.A2(n_682),
.B1(n_629),
.B2(n_705),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_720),
.A2(n_715),
.B1(n_612),
.B2(n_601),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_728),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_SL g771 ( 
.A(n_756),
.B(n_612),
.C(n_713),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_739),
.A2(n_707),
.B1(n_704),
.B2(n_616),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_726),
.B(n_645),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_726),
.A2(n_642),
.B1(n_624),
.B2(n_676),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_740),
.B(n_645),
.Y(n_775)
);

OA21x2_ASAP7_75t_L g776 ( 
.A1(n_744),
.A2(n_668),
.B(n_693),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_716),
.B(n_675),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_743),
.B(n_675),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_723),
.Y(n_779)
);

CKINVDCx11_ASAP7_75t_R g780 ( 
.A(n_753),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_725),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_716),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_743),
.B(n_688),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_735),
.A2(n_704),
.B1(n_616),
.B2(n_694),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_757),
.A2(n_616),
.B1(n_703),
.B2(n_700),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_724),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_SL g787 ( 
.A(n_741),
.B(n_10),
.C(n_13),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_766),
.A2(n_760),
.B1(n_765),
.B2(n_755),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_724),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_718),
.B(n_688),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_717),
.B(n_616),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_735),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_766),
.A2(n_688),
.B1(n_15),
.B2(n_17),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_738),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_718),
.B(n_14),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_741),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_722),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_765),
.B(n_18),
.C(n_20),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_722),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_735),
.A2(n_727),
.B1(n_766),
.B2(n_767),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_746),
.B(n_21),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_723),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_752),
.A2(n_21),
.B(n_22),
.Y(n_803)
);

AOI21xp33_ASAP7_75t_L g804 ( 
.A1(n_727),
.A2(n_22),
.B(n_24),
.Y(n_804)
);

BUFx12f_ASAP7_75t_L g805 ( 
.A(n_729),
.Y(n_805)
);

AOI221xp5_ASAP7_75t_L g806 ( 
.A1(n_755),
.A2(n_737),
.B1(n_767),
.B2(n_748),
.C(n_746),
.Y(n_806)
);

AOI221xp5_ASAP7_75t_L g807 ( 
.A1(n_737),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_748),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_722),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_719),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_719),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_718),
.B(n_73),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_735),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_730),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_766),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_763),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_738),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_718),
.B(n_35),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_754),
.B(n_37),
.Y(n_819)
);

AO22x2_ASAP7_75t_L g820 ( 
.A1(n_763),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_754),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_821)
);

AOI221xp5_ASAP7_75t_L g822 ( 
.A1(n_730),
.A2(n_729),
.B1(n_732),
.B2(n_751),
.C(n_762),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_786),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_789),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_768),
.A2(n_732),
.B1(n_750),
.B2(n_738),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_803),
.A2(n_761),
.B1(n_751),
.B2(n_738),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_774),
.A2(n_762),
.B(n_758),
.C(n_759),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_787),
.A2(n_761),
.B1(n_738),
.B2(n_750),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_769),
.A2(n_750),
.B1(n_738),
.B2(n_747),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_775),
.B(n_750),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_769),
.A2(n_736),
.B(n_749),
.Y(n_831)
);

AOI21xp33_ASAP7_75t_L g832 ( 
.A1(n_808),
.A2(n_761),
.B(n_736),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_777),
.B(n_734),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_810),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_798),
.A2(n_750),
.B1(n_763),
.B2(n_745),
.Y(n_835)
);

AOI221xp5_ASAP7_75t_L g836 ( 
.A1(n_796),
.A2(n_750),
.B1(n_721),
.B2(n_747),
.C(n_731),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_815),
.A2(n_747),
.B1(n_721),
.B2(n_764),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_802),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_811),
.Y(n_839)
);

OAI221xp5_ASAP7_75t_L g840 ( 
.A1(n_821),
.A2(n_721),
.B1(n_747),
.B2(n_764),
.C(n_731),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_794),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_L g842 ( 
.A1(n_821),
.A2(n_731),
.B1(n_734),
.B2(n_43),
.C(n_44),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_782),
.B(n_734),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_793),
.A2(n_734),
.B1(n_42),
.B2(n_44),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_819),
.B(n_734),
.Y(n_845)
);

OAI33xp33_ASAP7_75t_L g846 ( 
.A1(n_801),
.A2(n_41),
.A3(n_45),
.B1(n_734),
.B2(n_744),
.B3(n_745),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_807),
.A2(n_742),
.B1(n_749),
.B2(n_81),
.Y(n_847)
);

AOI211xp5_ASAP7_75t_L g848 ( 
.A1(n_804),
.A2(n_742),
.B(n_80),
.C(n_83),
.Y(n_848)
);

AO31x2_ASAP7_75t_L g849 ( 
.A1(n_816),
.A2(n_78),
.A3(n_84),
.B(n_88),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_773),
.B(n_89),
.Y(n_850)
);

OAI221xp5_ASAP7_75t_L g851 ( 
.A1(n_792),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.C(n_93),
.Y(n_851)
);

OAI22xp33_ASAP7_75t_L g852 ( 
.A1(n_788),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_779),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_781),
.A2(n_770),
.B1(n_822),
.B2(n_805),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_797),
.Y(n_855)
);

AOI222xp33_ASAP7_75t_L g856 ( 
.A1(n_792),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.C1(n_112),
.C2(n_113),
.Y(n_856)
);

OAI211xp5_ASAP7_75t_L g857 ( 
.A1(n_813),
.A2(n_116),
.B(n_118),
.C(n_122),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_814),
.Y(n_858)
);

AOI33xp33_ASAP7_75t_L g859 ( 
.A1(n_813),
.A2(n_126),
.A3(n_129),
.B1(n_130),
.B2(n_131),
.B3(n_133),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_785),
.A2(n_139),
.B(n_140),
.Y(n_860)
);

AOI222xp33_ASAP7_75t_L g861 ( 
.A1(n_820),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.C1(n_145),
.C2(n_146),
.Y(n_861)
);

OAI22xp33_ASAP7_75t_L g862 ( 
.A1(n_781),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_862)
);

INVx3_ASAP7_75t_SL g863 ( 
.A(n_795),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_820),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_818),
.B(n_159),
.Y(n_865)
);

NAND4xp25_ASAP7_75t_L g866 ( 
.A(n_806),
.B(n_160),
.C(n_161),
.D(n_162),
.Y(n_866)
);

OAI21xp33_ASAP7_75t_SL g867 ( 
.A1(n_800),
.A2(n_166),
.B(n_167),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_799),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_845),
.B(n_800),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_833),
.B(n_783),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_823),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_843),
.B(n_778),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_855),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_858),
.B(n_797),
.Y(n_874)
);

INVx8_ASAP7_75t_L g875 ( 
.A(n_841),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_824),
.B(n_790),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_834),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_868),
.B(n_809),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_839),
.B(n_809),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_830),
.B(n_820),
.Y(n_881)
);

NOR2x1p5_ASAP7_75t_L g882 ( 
.A(n_866),
.B(n_812),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_838),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_854),
.B(n_816),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_849),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_831),
.Y(n_886)
);

NAND2x1p5_ASAP7_75t_L g887 ( 
.A(n_841),
.B(n_776),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_849),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_826),
.B(n_776),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_863),
.B(n_776),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_840),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_827),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_829),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_861),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_837),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_832),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_835),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_864),
.B(n_784),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_861),
.B(n_825),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_828),
.B(n_784),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_892),
.B(n_780),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_877),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_871),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_871),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_894),
.A2(n_856),
.B1(n_842),
.B2(n_844),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_894),
.A2(n_856),
.B1(n_851),
.B2(n_857),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_SL g907 ( 
.A1(n_899),
.A2(n_862),
.B(n_852),
.Y(n_907)
);

NAND4xp25_ASAP7_75t_SL g908 ( 
.A(n_899),
.B(n_859),
.C(n_848),
.D(n_836),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_883),
.B(n_850),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_870),
.B(n_772),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_894),
.A2(n_860),
.B(n_847),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_871),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_892),
.A2(n_853),
.B(n_865),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_894),
.A2(n_846),
.B1(n_867),
.B2(n_812),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_883),
.B(n_817),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_SL g916 ( 
.A(n_882),
.B(n_771),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_878),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_881),
.B(n_794),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_881),
.B(n_805),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_903),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_904),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_912),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_918),
.B(n_890),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_919),
.B(n_890),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_917),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_915),
.B(n_896),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_902),
.B(n_878),
.Y(n_927)
);

NAND4xp25_ASAP7_75t_L g928 ( 
.A(n_905),
.B(n_896),
.C(n_886),
.D(n_897),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_910),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_909),
.B(n_869),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_902),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_902),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_902),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_911),
.A2(n_891),
.B(n_886),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_920),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_921),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_930),
.B(n_869),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_921),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_930),
.B(n_876),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_922),
.Y(n_940)
);

NAND5xp2_ASAP7_75t_L g941 ( 
.A(n_934),
.B(n_907),
.C(n_905),
.D(n_906),
.E(n_913),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_922),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_937),
.B(n_901),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_941),
.B(n_780),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_937),
.B(n_924),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_939),
.B(n_928),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_935),
.B(n_908),
.C(n_916),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_939),
.B(n_901),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_938),
.B(n_924),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_942),
.A2(n_926),
.B(n_929),
.Y(n_950)
);

O2A1O1Ixp5_ASAP7_75t_L g951 ( 
.A1(n_943),
.A2(n_926),
.B(n_932),
.C(n_933),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_948),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_949),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_947),
.B(n_923),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_SL g955 ( 
.A1(n_944),
.A2(n_946),
.B1(n_898),
.B2(n_893),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_955),
.B(n_945),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_953),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_954),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_SL g959 ( 
.A(n_952),
.B(n_950),
.C(n_931),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_951),
.A2(n_882),
.B1(n_898),
.B2(n_897),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_L g961 ( 
.A(n_959),
.B(n_914),
.C(n_895),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_923),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_958),
.B(n_936),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_956),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_960),
.B(n_927),
.Y(n_965)
);

NOR2x1_ASAP7_75t_L g966 ( 
.A(n_961),
.B(n_932),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_963),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_964),
.B(n_962),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_914),
.C(n_895),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_964),
.B(n_891),
.C(n_936),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_961),
.B(n_927),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_891),
.C(n_940),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_963),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_968),
.Y(n_974)
);

AOI33xp33_ASAP7_75t_L g975 ( 
.A1(n_967),
.A2(n_927),
.A3(n_900),
.B1(n_925),
.B2(n_878),
.B3(n_888),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_971),
.B(n_925),
.Y(n_976)
);

AOI221x1_ASAP7_75t_L g977 ( 
.A1(n_973),
.A2(n_812),
.B1(n_888),
.B2(n_884),
.C(n_877),
.Y(n_977)
);

NAND4xp25_ASAP7_75t_L g978 ( 
.A(n_966),
.B(n_791),
.C(n_884),
.D(n_900),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_972),
.B(n_970),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_969),
.B(n_876),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_968),
.B(n_874),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_974),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_976),
.Y(n_983)
);

NAND4xp25_ASAP7_75t_SL g984 ( 
.A(n_977),
.B(n_889),
.C(n_872),
.D(n_885),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_R g985 ( 
.A(n_979),
.B(n_981),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_978),
.B(n_872),
.Y(n_986)
);

XNOR2xp5_ASAP7_75t_L g987 ( 
.A(n_980),
.B(n_887),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_975),
.Y(n_988)
);

OAI332xp33_ASAP7_75t_L g989 ( 
.A1(n_974),
.A2(n_889),
.A3(n_885),
.B1(n_817),
.B2(n_870),
.B3(n_880),
.C1(n_879),
.C2(n_175),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_979),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_982),
.B(n_874),
.Y(n_991)
);

NAND4xp75_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_880),
.C(n_879),
.D(n_885),
.Y(n_992)
);

NOR2x1_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_877),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_985),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_988),
.B(n_887),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_986),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_987),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_L g998 ( 
.A(n_984),
.B(n_877),
.C(n_873),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_983),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_999),
.Y(n_1000)
);

OAI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_994),
.A2(n_887),
.B1(n_873),
.B2(n_875),
.C(n_172),
.Y(n_1001)
);

NAND4xp25_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_873),
.C(n_169),
.D(n_170),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_996),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_995),
.A2(n_875),
.B1(n_873),
.B2(n_174),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_L g1005 ( 
.A(n_991),
.B(n_168),
.C(n_173),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_998),
.A2(n_993),
.B1(n_992),
.B2(n_875),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_1000),
.B(n_1003),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_1004),
.Y(n_1008)
);

AND4x1_ASAP7_75t_L g1009 ( 
.A(n_1005),
.B(n_179),
.C(n_180),
.D(n_181),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1002),
.Y(n_1010)
);

NAND4xp25_ASAP7_75t_SL g1011 ( 
.A(n_1006),
.B(n_875),
.C(n_183),
.D(n_185),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_1007),
.Y(n_1012)
);

AOI31xp33_ASAP7_75t_L g1013 ( 
.A1(n_1010),
.A2(n_1001),
.A3(n_186),
.B(n_188),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1008),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_1009),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_1012),
.A2(n_1011),
.B(n_189),
.Y(n_1016)
);

XNOR2x1_ASAP7_75t_L g1017 ( 
.A(n_1014),
.B(n_182),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1017),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_1016),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1018),
.B(n_1015),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_1019),
.A2(n_1013),
.B1(n_191),
.B2(n_192),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1020),
.A2(n_190),
.B(n_193),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1021),
.A2(n_875),
.B1(n_195),
.B2(n_197),
.Y(n_1023)
);

OAI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_1023),
.A2(n_875),
.B1(n_199),
.B2(n_200),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_1022),
.A2(n_194),
.B1(n_201),
.B2(n_203),
.Y(n_1025)
);

AOI221xp5_ASAP7_75t_L g1026 ( 
.A1(n_1024),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.C(n_208),
.Y(n_1026)
);

AOI211xp5_ASAP7_75t_L g1027 ( 
.A1(n_1026),
.A2(n_1025),
.B(n_210),
.C(n_212),
.Y(n_1027)
);


endmodule