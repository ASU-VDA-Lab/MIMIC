module fake_jpeg_12876_n_390 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_0),
.B(n_7),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_55),
.B(n_57),
.Y(n_138)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_59),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_53),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_63),
.B(n_64),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_22),
.B(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_66),
.B(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_69),
.B(n_72),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_27),
.B(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_75),
.B(n_77),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_29),
.B(n_9),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_34),
.B(n_12),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

NAND2x1_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_0),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_35),
.Y(n_149)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_106),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_37),
.B(n_1),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_95),
.Y(n_137)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_2),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_101),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_48),
.Y(n_105)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_40),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_39),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_41),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_113),
.B(n_143),
.Y(n_220)
);

OA22x2_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_17),
.B1(n_31),
.B2(n_48),
.Y(n_116)
);

OR2x4_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_174),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_31),
.B1(n_51),
.B2(n_18),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_121),
.A2(n_134),
.B1(n_148),
.B2(n_151),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_71),
.A2(n_49),
.B1(n_51),
.B2(n_18),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_124),
.A2(n_136),
.B(n_142),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_41),
.B1(n_50),
.B2(n_45),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_49),
.B1(n_36),
.B2(n_47),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_36),
.B1(n_47),
.B2(n_46),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_89),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_101),
.B1(n_81),
.B2(n_70),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_67),
.A2(n_78),
.B1(n_107),
.B2(n_103),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_163),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_74),
.A2(n_53),
.B1(n_50),
.B2(n_45),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_61),
.A2(n_105),
.B(n_91),
.C(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_165),
.Y(n_190)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_111),
.B(n_108),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_105),
.A2(n_25),
.B(n_3),
.C(n_2),
.Y(n_165)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_87),
.B(n_2),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_57),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_94),
.B(n_96),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_178),
.B(n_185),
.Y(n_263)
);

AO22x2_ASAP7_75t_L g179 ( 
.A1(n_116),
.A2(n_102),
.B1(n_84),
.B2(n_70),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_35),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_194),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_197),
.Y(n_249)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_43),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_136),
.Y(n_243)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_33),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_191),
.B(n_193),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_121),
.A2(n_25),
.B1(n_113),
.B2(n_28),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_33),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_2),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_195),
.Y(n_251)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_139),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx4_ASAP7_75t_SL g199 ( 
.A(n_173),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_215),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_137),
.A2(n_3),
.B1(n_153),
.B2(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_203),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_202),
.B(n_205),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_137),
.B(n_132),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_138),
.B(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_138),
.B(n_119),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_207),
.B(n_210),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_119),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_216),
.Y(n_252)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_120),
.B(n_128),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_142),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_168),
.B(n_144),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_219),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_117),
.B(n_127),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_225),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_145),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_117),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_122),
.B(n_147),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_141),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_131),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_152),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_140),
.B(n_176),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_161),
.C(n_141),
.Y(n_248)
);

AND2x4_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_135),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_248),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_258),
.B1(n_272),
.B2(n_246),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_208),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_124),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_246),
.C(n_254),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_130),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_255),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_204),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_181),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_146),
.C(n_161),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_180),
.B(n_146),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_194),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_256),
.B(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_190),
.A2(n_221),
.B1(n_217),
.B2(n_189),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_221),
.A2(n_208),
.B1(n_189),
.B2(n_179),
.Y(n_272)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_179),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_277),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_255),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_279),
.B(n_283),
.Y(n_312)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_280),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_237),
.C(n_244),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_296),
.C(n_297),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_285),
.Y(n_314)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_179),
.B1(n_231),
.B2(n_228),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_236),
.B1(n_248),
.B2(n_250),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_265),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_286),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_182),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_288),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_231),
.B(n_182),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_298),
.B(n_299),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_263),
.B(n_183),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_295),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_209),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_187),
.C(n_195),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_199),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_233),
.A2(n_215),
.B(n_184),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_232),
.B(n_206),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_303),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_233),
.A2(n_213),
.B1(n_188),
.B2(n_177),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_301),
.A2(n_270),
.B1(n_251),
.B2(n_262),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_214),
.C(n_254),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_278),
.C(n_273),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_241),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_261),
.B(n_236),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_304),
.A2(n_298),
.B(n_290),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_240),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_319),
.C(n_315),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_313),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_297),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_234),
.B1(n_252),
.B2(n_267),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_259),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_324),
.C(n_302),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_321),
.A2(n_277),
.B(n_282),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_234),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_289),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_328),
.A2(n_337),
.B1(n_339),
.B2(n_341),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_285),
.Y(n_329)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_340),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_332),
.C(n_336),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_287),
.C(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_322),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_309),
.B1(n_313),
.B2(n_306),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_287),
.C(n_294),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_299),
.A3(n_284),
.B1(n_301),
.B2(n_287),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_235),
.Y(n_338)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_239),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_275),
.B(n_293),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_323),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_305),
.C(n_310),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_349),
.B1(n_352),
.B2(n_327),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_333),
.A2(n_320),
.B1(n_312),
.B2(n_308),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_328),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_332),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_335),
.B1(n_340),
.B2(n_312),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_342),
.C(n_331),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_356),
.A2(n_362),
.B1(n_311),
.B2(n_308),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_347),
.B(n_330),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_365),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_304),
.B(n_335),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_361),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_351),
.C(n_337),
.Y(n_370)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_346),
.Y(n_360)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

OA21x2_ASAP7_75t_SL g361 ( 
.A1(n_345),
.A2(n_323),
.B(n_322),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_317),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_317),
.B1(n_321),
.B2(n_325),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_363),
.A2(n_364),
.B1(n_353),
.B2(n_354),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_355),
.B(n_336),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_362),
.A2(n_348),
.B1(n_344),
.B2(n_343),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_366),
.B(n_274),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_354),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_369),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_362),
.C(n_365),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_371),
.A2(n_239),
.B(n_245),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_372),
.B(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_376),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_378),
.C(n_373),
.Y(n_382)
);

AOI322xp5_ASAP7_75t_L g376 ( 
.A1(n_366),
.A2(n_358),
.A3(n_280),
.B1(n_247),
.B2(n_292),
.C1(n_283),
.C2(n_300),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_270),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_377),
.A2(n_370),
.B(n_371),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_382),
.B(n_380),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_379),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_385),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_368),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_367),
.B(n_245),
.C(n_260),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_387),
.A2(n_251),
.B(n_262),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_388),
.Y(n_390)
);


endmodule