module fake_jpeg_9976_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_18),
.B1(n_19),
.B2(n_13),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_63),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_31),
.A3(n_34),
.B1(n_19),
.B2(n_17),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_62),
.B1(n_26),
.B2(n_23),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_61),
.B1(n_49),
.B2(n_43),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_16),
.B1(n_13),
.B2(n_17),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_16),
.B1(n_26),
.B2(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_43),
.B1(n_42),
.B2(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_68),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_31),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_73),
.B(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_48),
.C(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_48),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_35),
.B(n_15),
.C(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_64),
.B1(n_68),
.B2(n_38),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_88),
.B(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_38),
.B(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_54),
.B1(n_29),
.B2(n_24),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_69),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_88),
.C(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_103),
.B(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_65),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_73),
.B1(n_66),
.B2(n_71),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_102),
.B1(n_80),
.B2(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_76),
.B1(n_74),
.B2(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_11),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_92),
.C(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_80),
.B1(n_39),
.B2(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_121)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_24),
.B1(n_20),
.B2(n_11),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_20),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_116),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_102),
.B(n_94),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_2),
.C(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_126),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_108),
.C(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_112),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_126),
.A2(n_115),
.B1(n_108),
.B2(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_114),
.C(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_125),
.C(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_7),
.Y(n_134)
);

OAI321xp33_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.A3(n_130),
.B1(n_9),
.B2(n_10),
.C(n_8),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_130),
.C(n_9),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_9),
.C(n_10),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);


endmodule