module fake_jpeg_1729_n_105 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_7),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_33),
.Y(n_54)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_39),
.B(n_40),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_14),
.B(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_25),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_26),
.C(n_24),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_49),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_53),
.B1(n_56),
.B2(n_32),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_53)
);

NOR2x1_ASAP7_75t_R g55 ( 
.A(n_39),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_23),
.B1(n_20),
.B2(n_0),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_63),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_36),
.B1(n_30),
.B2(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_35),
.B1(n_13),
.B2(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_1),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_68),
.B1(n_50),
.B2(n_60),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_52),
.C(n_55),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_76),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_58),
.C(n_57),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_2),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_52),
.C(n_48),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_43),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_62),
.B(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_83),
.C(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_61),
.B(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_74),
.C(n_85),
.Y(n_93)
);

XNOR2x1_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_96),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_77),
.B(n_85),
.C(n_72),
.D(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_91),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_75),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_94),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_92),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_87),
.A3(n_13),
.B1(n_11),
.B2(n_10),
.C1(n_9),
.C2(n_75),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_10),
.C(n_11),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_13),
.Y(n_105)
);


endmodule