module fake_jpeg_13637_n_509 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_63),
.Y(n_103)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_32),
.B(n_16),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_92),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g116 ( 
.A(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_16),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_15),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_71),
.B(n_86),
.Y(n_134)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_14),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_25),
.B(n_14),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

CKINVDCx6p67_ASAP7_75t_R g153 ( 
.A(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_91),
.B(n_39),
.CON(n_143),
.SN(n_143)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_28),
.B(n_13),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_94),
.B(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_28),
.B(n_29),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_96),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_98),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_29),
.B(n_0),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_37),
.B(n_31),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_38),
.B1(n_35),
.B2(n_50),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_101),
.A2(n_102),
.B1(n_125),
.B2(n_129),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_53),
.A2(n_38),
.B1(n_35),
.B2(n_41),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_105),
.B(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_73),
.A2(n_21),
.B1(n_35),
.B2(n_38),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_57),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_35),
.B1(n_21),
.B2(n_30),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_51),
.A2(n_21),
.B1(n_22),
.B2(n_43),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_131),
.A2(n_137),
.B1(n_141),
.B2(n_144),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_78),
.A2(n_21),
.B1(n_30),
.B2(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_58),
.B(n_37),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_40),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_31),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_87),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_141)
);

NAND2x1_ASAP7_75t_SL g185 ( 
.A(n_143),
.B(n_40),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_55),
.A2(n_46),
.B1(n_19),
.B2(n_42),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_19),
.B1(n_42),
.B2(n_40),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_22),
.C(n_24),
.Y(n_158)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_54),
.B(n_46),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_139),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_180),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_33),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_166),
.B(n_172),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_167),
.A2(n_178),
.B(n_203),
.Y(n_249)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_170),
.Y(n_258)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_33),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_175),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_176),
.B(n_182),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_115),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_177),
.B(n_153),
.C(n_107),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_54),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_110),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_123),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_190),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_186),
.B(n_188),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_192),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_112),
.B(n_72),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_125),
.A2(n_59),
.B1(n_56),
.B2(n_93),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_193),
.B1(n_207),
.B2(n_142),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_128),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_131),
.A2(n_76),
.B1(n_81),
.B2(n_84),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_209),
.B1(n_118),
.B2(n_104),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_106),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_197),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_147),
.B(n_88),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_196),
.B(n_205),
.Y(n_256)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_143),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_199),
.Y(n_232)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_27),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_204),
.Y(n_235)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_202),
.Y(n_245)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

OR2x4_ASAP7_75t_L g203 ( 
.A(n_124),
.B(n_39),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_27),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_116),
.B(n_39),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_149),
.B(n_88),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_206),
.B(n_213),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_120),
.A2(n_82),
.B1(n_27),
.B2(n_24),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_210),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_116),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_24),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_122),
.Y(n_237)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_39),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_137),
.B(n_129),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_214),
.A2(n_225),
.B(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_119),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_221),
.C(n_238),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_174),
.A2(n_102),
.B1(n_104),
.B2(n_118),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_218),
.A2(n_248),
.B1(n_251),
.B2(n_195),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_167),
.B(n_153),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_161),
.A2(n_132),
.B(n_153),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_241),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_132),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_122),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_253),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_178),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_190),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_180),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_174),
.A2(n_140),
.B1(n_52),
.B2(n_96),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_197),
.B(n_123),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_0),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_0),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_160),
.B(n_66),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_0),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_208),
.A2(n_66),
.B1(n_106),
.B2(n_100),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_159),
.B(n_100),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_269),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_178),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_275),
.C(n_280),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_204),
.B(n_203),
.Y(n_266)
);

AOI21x1_ASAP7_75t_SL g332 ( 
.A1(n_266),
.A2(n_258),
.B(n_229),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_183),
.B1(n_163),
.B2(n_171),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_272),
.B1(n_285),
.B2(n_234),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_236),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_270),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_235),
.A2(n_241),
.B1(n_214),
.B2(n_219),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_239),
.B(n_187),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_236),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_278),
.Y(n_336)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_169),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_244),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_224),
.B1(n_250),
.B2(n_247),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_230),
.B(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_183),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_288),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_217),
.B(n_184),
.C(n_201),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_298),
.C(n_258),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_281),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_242),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_296),
.B1(n_223),
.B2(n_215),
.Y(n_333)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_199),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_299),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_168),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_257),
.B(n_202),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_244),
.B(n_170),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_212),
.B1(n_180),
.B2(n_175),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_198),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_223),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_107),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_234),
.B(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_33),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_240),
.B(n_209),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_181),
.Y(n_342)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_142),
.B1(n_149),
.B2(n_194),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_306),
.A2(n_296),
.B1(n_304),
.B2(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_311),
.A2(n_316),
.B1(n_317),
.B2(n_344),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_234),
.B1(n_251),
.B2(n_225),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_272),
.A2(n_250),
.B1(n_252),
.B2(n_222),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_289),
.A2(n_259),
.B1(n_261),
.B2(n_221),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_319),
.A2(n_324),
.B1(n_333),
.B2(n_304),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_226),
.B1(n_222),
.B2(n_227),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_245),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_326),
.B(n_328),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_264),
.A2(n_232),
.B(n_227),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_293),
.B(n_265),
.Y(n_358)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_297),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_330),
.B(n_347),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_335),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_229),
.C(n_233),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_338),
.C(n_286),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_233),
.C(n_260),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_346),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_343),
.A2(n_295),
.B1(n_306),
.B2(n_267),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_264),
.A2(n_142),
.B1(n_149),
.B2(n_181),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_273),
.B(n_1),
.Y(n_346)
);

AOI322xp5_ASAP7_75t_L g347 ( 
.A1(n_273),
.A2(n_48),
.A3(n_106),
.B1(n_68),
.B2(n_75),
.C1(n_83),
.C2(n_39),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_348),
.A2(n_363),
.B1(n_374),
.B2(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_375),
.C(n_377),
.Y(n_390)
);

A2O1A1O1Ixp25_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_274),
.B(n_283),
.C(n_266),
.D(n_293),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_358),
.B(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

XOR2x1_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_298),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_354),
.B(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_345),
.Y(n_356)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_345),
.Y(n_357)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_271),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_360),
.B(n_361),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_329),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_319),
.A2(n_292),
.B1(n_274),
.B2(n_297),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_334),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_364),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_310),
.B(n_283),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_366),
.B(n_371),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_339),
.B(n_313),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_370),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_346),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_291),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_311),
.A2(n_306),
.B1(n_277),
.B2(n_276),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_379),
.B1(n_314),
.B2(n_321),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_295),
.C(n_279),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_324),
.A2(n_301),
.B1(n_48),
.B2(n_4),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_335),
.C(n_337),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_378),
.B(n_380),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_316),
.A2(n_48),
.B1(n_2),
.B2(n_5),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_1),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_2),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_2),
.C(n_6),
.Y(n_410)
);

BUFx8_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_358),
.A2(n_327),
.B(n_344),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_398),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_309),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_386),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_338),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_381),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_373),
.A2(n_379),
.B1(n_350),
.B2(n_367),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_393),
.A2(n_403),
.B1(n_376),
.B2(n_368),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_329),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_395),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_308),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_399),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_363),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_348),
.A2(n_342),
.B1(n_336),
.B2(n_318),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_405),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_359),
.A2(n_314),
.B1(n_321),
.B2(n_323),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_325),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_407),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_331),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_331),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_375),
.C(n_359),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_6),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_417),
.C(n_411),
.Y(n_438)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_354),
.C(n_350),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_387),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_428),
.B1(n_430),
.B2(n_432),
.Y(n_441)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_421),
.B(n_385),
.Y(n_451)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_391),
.Y(n_423)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

HAxp5_ASAP7_75t_SL g424 ( 
.A(n_383),
.B(n_352),
.CON(n_424),
.SN(n_424)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_427),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_426),
.B(n_410),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_384),
.B(n_368),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_371),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_429),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_403),
.A2(n_365),
.B1(n_370),
.B2(n_380),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_392),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_7),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_434),
.C(n_400),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_7),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_436),
.Y(n_460)
);

OAI321xp33_ASAP7_75t_L g437 ( 
.A1(n_419),
.A2(n_399),
.A3(n_382),
.B1(n_389),
.B2(n_401),
.C(n_395),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_440),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_416),
.C(n_413),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_431),
.B(n_419),
.Y(n_439)
);

XOR2x2_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_451),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_390),
.C(n_407),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_412),
.A2(n_431),
.B1(n_417),
.B2(n_427),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_10),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_390),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_443),
.B(n_446),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_430),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_412),
.A2(n_404),
.B1(n_382),
.B2(n_405),
.Y(n_447)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_447),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_414),
.B(n_397),
.Y(n_450)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_450),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_424),
.A2(n_395),
.B(n_386),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_453),
.A2(n_432),
.B(n_428),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_444),
.A2(n_421),
.B1(n_413),
.B2(n_423),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_445),
.B1(n_451),
.B2(n_448),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_411),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_458),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_459),
.A2(n_470),
.B(n_441),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_404),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_464),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_422),
.C(n_420),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_8),
.C(n_9),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_11),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_449),
.A2(n_9),
.B(n_10),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_467),
.A2(n_459),
.B(n_470),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_9),
.Y(n_469)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_469),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_471),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_462),
.B(n_445),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_472),
.B(n_479),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_444),
.C(n_449),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_475),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_437),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_466),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_460),
.B(n_448),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_452),
.C(n_454),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_481),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_456),
.A2(n_452),
.B1(n_454),
.B2(n_11),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_483),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_468),
.C(n_478),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_486),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_461),
.C(n_458),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_455),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_492),
.Y(n_499)
);

OAI321xp33_ASAP7_75t_L g493 ( 
.A1(n_477),
.A2(n_12),
.A3(n_465),
.B1(n_466),
.B2(n_469),
.C(n_471),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_493),
.A2(n_485),
.B1(n_490),
.B2(n_489),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_480),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_487),
.A2(n_474),
.B(n_469),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_497),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_485),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_498),
.A2(n_499),
.B(n_494),
.Y(n_503)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_496),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_500),
.B(n_502),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_503),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_504),
.Y(n_506)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_506),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_507),
.B(n_501),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_505),
.Y(n_509)
);


endmodule