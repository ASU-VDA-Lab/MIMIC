module fake_jpeg_25415_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_22),
.Y(n_44)
);

NOR2x1_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_10),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_28),
.B(n_20),
.C(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_12),
.B1(n_11),
.B2(n_13),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_37),
.B1(n_27),
.B2(n_20),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_12),
.B1(n_18),
.B2(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_12),
.B1(n_24),
.B2(n_18),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_36),
.B(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_30),
.C(n_35),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_35),
.C(n_36),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_39),
.B(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_23),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_68),
.C(n_31),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_65),
.B(n_67),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_32),
.B(n_34),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_14),
.B(n_33),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_49),
.C(n_56),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_52),
.C(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_49),
.C(n_14),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_48),
.B1(n_45),
.B2(n_58),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_75),
.B(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_53),
.B1(n_38),
.B2(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_62),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_63),
.C(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_85),
.C(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_83),
.B1(n_74),
.B2(n_71),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_19),
.Y(n_82)
);

OA21x2_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_19),
.B(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_29),
.C(n_19),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_72),
.B(n_78),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_92),
.Y(n_96)
);

OAI31xp33_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_29),
.A3(n_2),
.B(n_3),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_81),
.B1(n_79),
.B2(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_1),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_29),
.C(n_13),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_1),
.B(n_2),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_92),
.C(n_88),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_87),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.C(n_100),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_8),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_9),
.B(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_102),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_105),
.Y(n_107)
);


endmodule