module fake_jpeg_3794_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_18),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.C(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_4),
.C(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_23),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_10),
.B(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_12),
.B1(n_11),
.B2(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_15),
.B1(n_14),
.B2(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_26),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_34),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_27),
.B(n_28),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_37),
.C(n_34),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_46),
.B(n_39),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_38),
.Y(n_50)
);

OA21x2_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_10),
.B(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_51),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_47),
.B1(n_4),
.B2(n_5),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_55),
.B(n_52),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_6),
.B(n_2),
.Y(n_60)
);


endmodule