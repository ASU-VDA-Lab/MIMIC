module fake_jpeg_29500_n_431 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_47),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_42),
.B(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_70),
.Y(n_123)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_23),
.B(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

CKINVDCx6p67_ASAP7_75t_R g125 ( 
.A(n_74),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_76),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_79),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_28),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_83),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g136 ( 
.A(n_82),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_46),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_36),
.B(n_7),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_41),
.B1(n_45),
.B2(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_94),
.A2(n_97),
.B1(n_100),
.B2(n_62),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_22),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_95),
.B(n_99),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_37),
.B1(n_45),
.B2(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_38),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_44),
.B1(n_38),
.B2(n_29),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_18),
.B1(n_26),
.B2(n_34),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_27),
.B1(n_34),
.B2(n_68),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_110),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_43),
.B1(n_29),
.B2(n_44),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_118),
.B1(n_142),
.B2(n_124),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_43),
.B1(n_34),
.B2(n_27),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_17),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_128),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_17),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_47),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_12),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_34),
.B1(n_27),
.B2(n_17),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_158),
.Y(n_194)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_144),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_63),
.B1(n_77),
.B2(n_73),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_76),
.C(n_84),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_161),
.C(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_151),
.Y(n_209)
);

BUFx2_ASAP7_75t_SL g149 ( 
.A(n_125),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_149),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_99),
.B(n_91),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_152),
.A2(n_162),
.B1(n_169),
.B2(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_79),
.B1(n_69),
.B2(n_67),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_119),
.B1(n_104),
.B2(n_125),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_155),
.A2(n_177),
.B1(n_183),
.B2(n_186),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_109),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_156),
.A2(n_173),
.B1(n_180),
.B2(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_163),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_30),
.B(n_27),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_107),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_103),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_11),
.B(n_15),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_168),
.B(n_174),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_11),
.B(n_15),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_107),
.A2(n_10),
.B1(n_13),
.B2(n_4),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_185),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_46),
.B1(n_10),
.B2(n_4),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_46),
.B1(n_11),
.B2(n_5),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_129),
.A2(n_46),
.B1(n_11),
.B2(n_5),
.Y(n_174)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_98),
.A2(n_46),
.B1(n_1),
.B2(n_0),
.Y(n_175)
);

AO21x2_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_125),
.B(n_149),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

BUFx2_ASAP7_75t_SL g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_113),
.A2(n_135),
.B1(n_130),
.B2(n_111),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_12),
.B1(n_13),
.B2(n_0),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_188),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_0),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_129),
.A2(n_1),
.B1(n_130),
.B2(n_127),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_1),
.B1(n_133),
.B2(n_127),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_104),
.B1(n_133),
.B2(n_114),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_198),
.A2(n_215),
.B1(n_216),
.B2(n_219),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_201),
.B1(n_211),
.B2(n_180),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_122),
.B1(n_121),
.B2(n_93),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_131),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_218),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_152),
.B(n_169),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_121),
.B1(n_122),
.B2(n_105),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_148),
.A2(n_115),
.B1(n_117),
.B2(n_102),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_155),
.A2(n_115),
.B1(n_119),
.B2(n_117),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_137),
.Y(n_218)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_136),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_229),
.C(n_190),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_174),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_136),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_230),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_102),
.B(n_137),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_210),
.B(n_215),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_170),
.B(n_103),
.C(n_105),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_151),
.B(n_103),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_161),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_232),
.B(n_252),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_171),
.B(n_184),
.C(n_146),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_233),
.B(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_145),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_245),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_213),
.B(n_182),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_168),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_239),
.B(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_163),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_246),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_217),
.A2(n_179),
.B1(n_189),
.B2(n_165),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_150),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_196),
.B(n_173),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_248),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_191),
.B(n_187),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_253),
.C(n_256),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_178),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_203),
.A2(n_153),
.B1(n_175),
.B2(n_144),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_254),
.A2(n_210),
.B1(n_207),
.B2(n_225),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_175),
.B1(n_162),
.B2(n_166),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_255),
.A2(n_260),
.B1(n_264),
.B2(n_199),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_175),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_209),
.B(n_181),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_154),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_251),
.C(n_252),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_203),
.A2(n_165),
.B(n_176),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_214),
.A2(n_1),
.B1(n_176),
.B2(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_197),
.B(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_204),
.B(n_194),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_268),
.B(n_204),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_201),
.B(n_211),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_212),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_271),
.A2(n_246),
.B(n_259),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_282),
.B(n_266),
.C(n_239),
.D(n_232),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_210),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_280),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_241),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_278),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_240),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_231),
.B(n_210),
.C(n_200),
.D(n_202),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_255),
.A2(n_210),
.B1(n_231),
.B2(n_200),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_291),
.B1(n_268),
.B2(n_264),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_274),
.C(n_245),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_207),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_293),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_292),
.A2(n_296),
.B1(n_254),
.B2(n_257),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_219),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_241),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_295),
.B(n_301),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_260),
.A2(n_202),
.B1(n_225),
.B2(n_228),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_205),
.B1(n_228),
.B2(n_193),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_308),
.B1(n_313),
.B2(n_315),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_307),
.C(n_324),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_253),
.C(n_245),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_234),
.B1(n_267),
.B2(n_256),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_309),
.A2(n_325),
.B1(n_293),
.B2(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_248),
.B1(n_234),
.B2(n_238),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_234),
.B1(n_258),
.B2(n_246),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_320),
.B(n_327),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_318),
.Y(n_332)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_236),
.B(n_235),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_262),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_310),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_233),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_294),
.A2(n_244),
.B1(n_265),
.B2(n_262),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_193),
.B(n_249),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_287),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_333),
.A2(n_341),
.B1(n_342),
.B2(n_352),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_334),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_310),
.B(n_277),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_344),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_269),
.B(n_289),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_350),
.B(n_275),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_269),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_347),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_309),
.A2(n_298),
.B1(n_273),
.B2(n_269),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_311),
.A2(n_298),
.B1(n_278),
.B2(n_282),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_303),
.B(n_270),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_279),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_275),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_321),
.B(n_270),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_351),
.B(n_314),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_298),
.B1(n_282),
.B2(n_280),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_279),
.C(n_290),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_308),
.C(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_372),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_305),
.B1(n_321),
.B2(n_315),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_357),
.A2(n_359),
.B1(n_331),
.B2(n_350),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_341),
.A2(n_320),
.B1(n_319),
.B2(n_328),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_325),
.B1(n_290),
.B2(n_288),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_366),
.B1(n_373),
.B2(n_342),
.Y(n_386)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_363),
.Y(n_379)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_296),
.B1(n_319),
.B2(n_322),
.Y(n_366)
);

XOR2x1_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_312),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_370),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_297),
.C(n_284),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_371),
.C(n_338),
.Y(n_377)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_284),
.C(n_318),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_364),
.B(n_353),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_382),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_377),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_357),
.A2(n_340),
.B1(n_350),
.B2(n_337),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_358),
.A2(n_330),
.B1(n_347),
.B2(n_345),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_352),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_385),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_332),
.C(n_335),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_360),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_335),
.B1(n_332),
.B2(n_345),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_387),
.Y(n_389)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_388),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_390),
.B(n_385),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_368),
.B(n_383),
.Y(n_393)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_379),
.A2(n_367),
.B(n_356),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_394),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_369),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_399),
.Y(n_405)
);

AO22x1_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_359),
.B1(n_372),
.B2(n_358),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_376),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_389),
.A2(n_396),
.B1(n_397),
.B2(n_400),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_406),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_404),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_396),
.A2(n_380),
.B1(n_382),
.B2(n_378),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_391),
.A2(n_378),
.B1(n_374),
.B2(n_379),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_361),
.C(n_286),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_361),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_275),
.C(n_208),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_392),
.A2(n_374),
.B(n_354),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_409),
.A2(n_302),
.B(n_300),
.Y(n_413)
);

AOI322xp5_ASAP7_75t_L g412 ( 
.A1(n_410),
.A2(n_398),
.A3(n_355),
.B1(n_370),
.B2(n_363),
.C1(n_362),
.C2(n_304),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_413),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g414 ( 
.A1(n_405),
.A2(n_301),
.A3(n_300),
.B1(n_299),
.B2(n_329),
.C1(n_377),
.C2(n_275),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_416),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_418),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_402),
.A2(n_205),
.B(n_208),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_411),
.A2(n_403),
.B(n_401),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_419),
.A2(n_420),
.B(n_415),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_417),
.A2(n_409),
.B(n_408),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_421),
.B(n_407),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_424),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_415),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_428),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_427),
.B1(n_426),
.B2(n_422),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_430),
.B(n_406),
.Y(n_431)
);


endmodule