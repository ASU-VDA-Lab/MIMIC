module fake_jpeg_2662_n_217 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_217);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_0),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_1),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_53),
.C(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_74),
.Y(n_105)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_64),
.B1(n_65),
.B2(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_97),
.B1(n_73),
.B2(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_68),
.B1(n_57),
.B2(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_60),
.B1(n_57),
.B2(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_64),
.B1(n_65),
.B2(n_58),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_79),
.B1(n_74),
.B2(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_111),
.B1(n_79),
.B2(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_91),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_89),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_72),
.B1(n_73),
.B2(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_87),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_91),
.B1(n_92),
.B2(n_85),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_100),
.B1(n_109),
.B2(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_129),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_89),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_49),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_49),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_71),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_131),
.B1(n_117),
.B2(n_118),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_46),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_100),
.B1(n_92),
.B2(n_104),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_103),
.B1(n_52),
.B2(n_50),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_155),
.B1(n_153),
.B2(n_143),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_63),
.B(n_70),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_153),
.B(n_69),
.Y(n_163)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_67),
.B(n_50),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_161),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_69),
.A3(n_59),
.B1(n_5),
.B2(n_6),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_171),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_154),
.B(n_142),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_176),
.B(n_180),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_176),
.B1(n_168),
.B2(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_168),
.B1(n_159),
.B2(n_144),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_10),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_174),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_11),
.B(n_12),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_44),
.B(n_43),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_138),
.B(n_29),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_14),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_187),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_192),
.B1(n_167),
.B2(n_166),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_42),
.C(n_40),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_193),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_21),
.C2(n_22),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_162),
.A3(n_182),
.B1(n_25),
.B2(n_23),
.C1(n_24),
.C2(n_32),
.Y(n_202)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.C(n_22),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_170),
.B1(n_175),
.B2(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_182),
.B1(n_178),
.B2(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_199),
.Y(n_206)
);

AOI321xp33_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_163),
.A3(n_179),
.B1(n_172),
.B2(n_169),
.C(n_180),
.Y(n_198)
);

AOI31xp67_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_203),
.A3(n_194),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_189),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_35),
.B(n_37),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_195),
.B(n_184),
.C(n_187),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_207),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_209),
.B(n_38),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_192),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_208),
.C(n_198),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_39),
.C(n_24),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_215),
.B(n_23),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_25),
.Y(n_217)
);


endmodule