module fake_jpeg_11616_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp33_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g16 ( 
.A(n_12),
.B(n_7),
.C(n_8),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_14),
.B1(n_10),
.B2(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_21),
.B1(n_0),
.B2(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_8),
.B1(n_7),
.B2(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_13),
.B1(n_10),
.B2(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_29),
.C(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_30),
.C(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_21),
.B1(n_15),
.B2(n_17),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_27),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_30),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_28),
.C(n_26),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_42),
.C(n_28),
.Y(n_49)
);

OAI321xp33_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_46),
.A3(n_45),
.B1(n_35),
.B2(n_6),
.C(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_50),
.Y(n_52)
);


endmodule