module real_jpeg_11934_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_249, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_249;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_59),
.B1(n_62),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_78),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_29),
.B1(n_37),
.B2(n_78),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_29),
.B1(n_37),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_4),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_7),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_8),
.A2(n_29),
.B1(n_37),
.B2(n_68),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_10),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_10),
.A2(n_59),
.B1(n_62),
.B2(n_109),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_109),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_29),
.B1(n_37),
.B2(n_109),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_43),
.B1(n_59),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_11),
.A2(n_29),
.B1(n_37),
.B2(n_43),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_12),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_14),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_14),
.A2(n_29),
.B1(n_37),
.B2(n_70),
.Y(n_194)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_15),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_15),
.B(n_62),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_15),
.A2(n_64),
.B(n_166),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_99),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_15),
.A2(n_45),
.B(n_49),
.C(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_15),
.B(n_105),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_15),
.B(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_15),
.B(n_85),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_15),
.A2(n_62),
.B(n_157),
.Y(n_220)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_17),
.A2(n_29),
.B1(n_37),
.B2(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_17),
.A2(n_53),
.B1(n_59),
.B2(n_62),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_131),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_21),
.B(n_113),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_22),
.A2(n_23),
.B1(n_80),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_26),
.B(n_40),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_27),
.A2(n_32),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_28),
.A2(n_33),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_28),
.A2(n_33),
.B(n_88),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_28),
.A2(n_33),
.B1(n_95),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_33),
.B1(n_147),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_28),
.A2(n_33),
.B1(n_160),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_28),
.A2(n_33),
.B1(n_99),
.B2(n_206),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_28),
.A2(n_33),
.B1(n_199),
.B2(n_206),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_29),
.B(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_37),
.A2(n_50),
.B(n_99),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_42),
.A2(n_47),
.B1(n_85),
.B2(n_151),
.Y(n_169)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_45),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_44),
.A2(n_62),
.A3(n_74),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_45),
.B(n_75),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_46),
.A2(n_51),
.B1(n_150),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_47),
.A2(n_84),
.B1(n_85),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_47),
.A2(n_85),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_47),
.A2(n_85),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_47),
.A2(n_85),
.B1(n_185),
.B2(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_57),
.A2(n_58),
.B1(n_108),
.B2(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_62),
.Y(n_97)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_99),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_76),
.B1(n_79),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_72),
.A2(n_76),
.B1(n_102),
.B2(n_143),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_72),
.A2(n_76),
.B1(n_141),
.B2(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_80),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_91),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_100),
.C(n_106),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_92),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_100),
.B(n_106),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_105),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_233),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_177),
.B(n_232),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_161),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_137),
.B(n_161),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.C(n_152),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_138),
.B(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_144),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_145),
.C(n_146),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_172),
.B2(n_176),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_162),
.B(n_173),
.C(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_168),
.C(n_171),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_226),
.B(n_231),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_215),
.B(n_225),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_195),
.B(n_214),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_191),
.C(n_193),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_203),
.B(n_213),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_201),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_209),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_221),
.C(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);


endmodule