module real_aes_11867_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g209 ( .A(n_0), .B(n_182), .Y(n_209) );
XOR2xp5_ASAP7_75t_L g712 ( .A(n_1), .B(n_474), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_2), .B(n_62), .Y(n_501) );
AND2x2_ASAP7_75t_L g580 ( .A(n_2), .B(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_2), .Y(n_612) );
INVx1_ASAP7_75t_L g654 ( .A(n_2), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_3), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_4), .B(n_143), .Y(n_207) );
INVx2_ASAP7_75t_L g487 ( .A(n_5), .Y(n_487) );
OR2x2_ASAP7_75t_L g670 ( .A(n_5), .B(n_485), .Y(n_670) );
BUFx2_ASAP7_75t_L g481 ( .A(n_6), .Y(n_481) );
BUFx2_ASAP7_75t_L g496 ( .A(n_6), .Y(n_496) );
INVx1_ASAP7_75t_L g563 ( .A(n_6), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_7), .B(n_192), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_8), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_9), .A2(n_50), .B1(n_565), .B2(n_572), .Y(n_564) );
INVx1_ASAP7_75t_L g664 ( .A(n_9), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_10), .B(n_138), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_11), .B(n_117), .Y(n_236) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_11), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_12), .B(n_138), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_13), .A2(n_23), .B1(n_550), .B2(n_552), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_13), .A2(n_23), .B1(n_578), .B2(n_586), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_14), .B(n_124), .Y(n_163) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_15), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_16), .B(n_138), .Y(n_144) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_17), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_18), .B(n_192), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_19), .A2(n_46), .B1(n_529), .B2(n_533), .Y(n_528) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_19), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_20), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_21), .B(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g685 ( .A(n_22), .Y(n_685) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_25), .B(n_117), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_26), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g485 ( .A(n_27), .Y(n_485) );
INVx1_ASAP7_75t_L g514 ( .A(n_27), .Y(n_514) );
NAND2xp33_ASAP7_75t_SL g162 ( .A(n_28), .B(n_89), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_28), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_28), .Y(n_681) );
INVx1_ASAP7_75t_L g544 ( .A(n_29), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_29), .A2(n_595), .B1(n_598), .B2(n_614), .C(n_627), .Y(n_594) );
INVx1_ASAP7_75t_L g642 ( .A(n_30), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_30), .A2(n_40), .B1(n_668), .B2(n_671), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_31), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_32), .B(n_122), .Y(n_239) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_33), .A2(n_55), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_34), .B(n_147), .Y(n_194) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_35), .A2(n_40), .B1(n_644), .B2(n_647), .C(n_650), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_35), .A2(n_59), .B1(n_673), .B2(n_675), .Y(n_672) );
AND2x6_ASAP7_75t_L g82 ( .A(n_36), .B(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_36), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_36), .B(n_698), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_37), .B(n_154), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_38), .B(n_154), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_39), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_41), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_42), .Y(n_203) );
INVx1_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_43), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_44), .B(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_45), .Y(n_689) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_46), .Y(n_626) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_47), .B(n_89), .Y(n_160) );
INVx1_ASAP7_75t_L g548 ( .A(n_48), .Y(n_548) );
OAI211xp5_ASAP7_75t_SL g629 ( .A1(n_48), .A2(n_630), .B(n_635), .C(n_655), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_49), .Y(n_478) );
INVx1_ASAP7_75t_L g660 ( .A(n_50), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_51), .B(n_124), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_52), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_53), .B(n_179), .Y(n_216) );
INVx2_ASAP7_75t_L g505 ( .A(n_54), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_56), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_57), .B(n_173), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_58), .B(n_147), .Y(n_241) );
INVx1_ASAP7_75t_L g639 ( .A(n_59), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_60), .Y(n_688) );
BUFx10_ASAP7_75t_L g707 ( .A(n_61), .Y(n_707) );
INVx2_ASAP7_75t_L g581 ( .A(n_62), .Y(n_581) );
INVx1_ASAP7_75t_L g613 ( .A(n_62), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_63), .B(n_117), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_64), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_65), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_66), .B(n_138), .Y(n_188) );
INVx2_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_68), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_69), .B(n_114), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_70), .B(n_192), .Y(n_220) );
INVx2_ASAP7_75t_L g506 ( .A(n_71), .Y(n_506) );
INVx1_ASAP7_75t_L g522 ( .A(n_72), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_73), .Y(n_141) );
INVx1_ASAP7_75t_L g527 ( .A(n_74), .Y(n_527) );
BUFx3_ASAP7_75t_L g490 ( .A(n_75), .Y(n_490) );
INVx1_ASAP7_75t_L g519 ( .A(n_75), .Y(n_519) );
BUFx3_ASAP7_75t_L g492 ( .A(n_76), .Y(n_492) );
INVx1_ASAP7_75t_L g521 ( .A(n_76), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_472), .Y(n_77) );
AND2x2_ASAP7_75t_L g78 ( .A(n_79), .B(n_84), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx8_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx2_ASAP7_75t_SL g145 ( .A(n_81), .Y(n_145) );
INVx8_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OAI21x1_ASAP7_75t_L g186 ( .A1(n_82), .A2(n_187), .B(n_190), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_82), .A2(n_125), .B(n_202), .C(n_205), .Y(n_201) );
OAI21x1_ASAP7_75t_SL g213 ( .A1(n_82), .A2(n_214), .B(n_217), .Y(n_213) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
AO21x1_ASAP7_75t_L g723 ( .A1(n_85), .A2(n_724), .B(n_725), .Y(n_723) );
NAND2xp33_ASAP7_75t_L g85 ( .A(n_86), .B(n_91), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx2_ASAP7_75t_L g219 ( .A(n_89), .Y(n_219) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_90), .Y(n_117) );
INVx2_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
INVx1_ASAP7_75t_L g180 ( .A(n_90), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_L g140 ( .A1(n_91), .A2(n_141), .B(n_142), .C(n_144), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_91), .A2(n_188), .B(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_91), .A2(n_192), .B(n_215), .C(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_91), .A2(n_239), .B(n_240), .Y(n_238) );
INVx5_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx5_ASAP7_75t_L g118 ( .A(n_92), .Y(n_118) );
BUFx12f_ASAP7_75t_L g208 ( .A(n_92), .Y(n_208) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND4xp75_ASAP7_75t_L g96 ( .A(n_97), .B(n_356), .C(n_400), .D(n_447), .Y(n_96) );
NOR2x1_ASAP7_75t_L g97 ( .A(n_98), .B(n_306), .Y(n_97) );
NAND2xp5_ASAP7_75t_SL g98 ( .A(n_99), .B(n_273), .Y(n_98) );
AOI321xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_165), .A3(n_195), .B1(n_223), .B2(n_242), .C(n_253), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NOR2x1_ASAP7_75t_L g102 ( .A(n_103), .B(n_129), .Y(n_102) );
AND2x4_ASAP7_75t_SL g349 ( .A(n_103), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g355 ( .A(n_103), .Y(n_355) );
INVx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g276 ( .A(n_104), .B(n_130), .Y(n_276) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_104), .Y(n_288) );
AND2x4_ASAP7_75t_L g324 ( .A(n_104), .B(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g281 ( .A(n_105), .Y(n_281) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g293 ( .A(n_106), .Y(n_293) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_111), .B(n_127), .Y(n_106) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_107), .A2(n_133), .B(n_146), .Y(n_132) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_107), .A2(n_201), .B(n_209), .Y(n_200) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_107), .A2(n_234), .B(n_241), .Y(n_233) );
BUFx5_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_108), .Y(n_128) );
INVx1_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g149 ( .A(n_109), .Y(n_149) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_119), .B(n_126), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_118), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g124 ( .A(n_115), .Y(n_124) );
INVx2_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
INVx2_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_117), .A2(n_122), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx2_ASAP7_75t_SL g125 ( .A(n_118), .Y(n_125) );
INVx2_ASAP7_75t_SL g139 ( .A(n_118), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_118), .A2(n_158), .B(n_159), .C(n_160), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_118), .A2(n_172), .B(n_174), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B(n_125), .Y(n_119) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_125), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21x1_ASAP7_75t_L g175 ( .A1(n_125), .A2(n_176), .B(n_177), .Y(n_175) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_126), .A2(n_235), .B(n_238), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_150), .Y(n_129) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_130), .A2(n_254), .B1(n_258), .B2(n_266), .Y(n_253) );
AND2x4_ASAP7_75t_SL g330 ( .A(n_130), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_131), .B(n_292), .Y(n_313) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g230 ( .A(n_132), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_145), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B(n_139), .Y(n_134) );
INVx5_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_139), .A2(n_191), .B(n_193), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_139), .A2(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_145), .A2(n_157), .B(n_161), .Y(n_156) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_145), .A2(n_171), .B(n_175), .Y(n_170) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
INVx1_ASAP7_75t_L g300 ( .A(n_150), .Y(n_300) );
INVx1_ASAP7_75t_L g386 ( .A(n_150), .Y(n_386) );
INVx1_ASAP7_75t_L g404 ( .A(n_150), .Y(n_404) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g331 ( .A(n_151), .B(n_293), .Y(n_331) );
AND2x2_ASAP7_75t_L g410 ( .A(n_151), .B(n_352), .Y(n_410) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_152), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_152), .B(n_293), .Y(n_398) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g286 ( .A(n_153), .B(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_153), .Y(n_373) );
OAI21x1_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_164), .Y(n_153) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_154), .A2(n_186), .B(n_194), .Y(n_185) );
INVx2_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g470 ( .A(n_167), .B(n_245), .Y(n_470) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g317 ( .A(n_168), .Y(n_317) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_184), .Y(n_168) );
AND2x2_ASAP7_75t_L g250 ( .A(n_169), .B(n_185), .Y(n_250) );
BUFx2_ASAP7_75t_L g271 ( .A(n_169), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_181), .B(n_183), .Y(n_169) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_170), .A2(n_181), .B(n_183), .Y(n_265) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g192 ( .A(n_180), .Y(n_192) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_182), .A2(n_213), .B(n_221), .Y(n_212) );
AND2x2_ASAP7_75t_L g247 ( .A(n_184), .B(n_211), .Y(n_247) );
INVx1_ASAP7_75t_L g261 ( .A(n_184), .Y(n_261) );
INVx1_ASAP7_75t_L g269 ( .A(n_184), .Y(n_269) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_184), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g343 ( .A(n_184), .Y(n_343) );
AND2x2_ASAP7_75t_L g443 ( .A(n_184), .B(n_210), .Y(n_443) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_196), .A2(n_466), .B1(n_467), .B2(n_468), .C(n_469), .Y(n_465) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x6_ASAP7_75t_L g316 ( .A(n_197), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g411 ( .A(n_198), .B(n_250), .Y(n_411) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_199), .B(n_211), .Y(n_252) );
AND2x2_ASAP7_75t_L g263 ( .A(n_199), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g268 ( .A(n_199), .Y(n_268) );
AND2x2_ASAP7_75t_L g303 ( .A(n_199), .B(n_281), .Y(n_303) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g246 ( .A(n_200), .Y(n_246) );
AND2x2_ASAP7_75t_L g347 ( .A(n_200), .B(n_264), .Y(n_347) );
AND2x2_ASAP7_75t_L g367 ( .A(n_200), .B(n_212), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_208), .A2(n_218), .B(n_220), .Y(n_217) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
INVxp67_ASAP7_75t_SL g260 ( .A(n_211), .Y(n_260) );
INVx1_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
INVx1_ASAP7_75t_L g296 ( .A(n_211), .Y(n_296) );
AND2x2_ASAP7_75t_L g344 ( .A(n_211), .B(n_268), .Y(n_344) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_211), .Y(n_394) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
AND2x4_ASAP7_75t_L g318 ( .A(n_225), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g362 ( .A(n_225), .Y(n_362) );
AND2x2_ASAP7_75t_L g446 ( .A(n_225), .B(n_279), .Y(n_446) );
OR2x2_ASAP7_75t_L g471 ( .A(n_225), .B(n_320), .Y(n_471) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_226), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g351 ( .A(n_226), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g354 ( .A(n_228), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g365 ( .A(n_228), .B(n_280), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_228), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g464 ( .A(n_228), .B(n_256), .Y(n_464) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g257 ( .A(n_229), .B(n_232), .Y(n_257) );
INVx1_ASAP7_75t_L g335 ( .A(n_229), .Y(n_335) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g279 ( .A(n_230), .B(n_232), .Y(n_279) );
INVx1_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
BUFx2_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g287 ( .A(n_232), .Y(n_287) );
INVx1_ASAP7_75t_L g372 ( .A(n_232), .Y(n_372) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_248), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g282 ( .A(n_244), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_245), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_245), .B(n_250), .Y(n_337) );
OR2x2_ASAP7_75t_L g379 ( .A(n_245), .B(n_380), .Y(n_379) );
INVx4_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x4_ASAP7_75t_L g305 ( .A(n_247), .B(n_283), .Y(n_305) );
INVx1_ASAP7_75t_L g380 ( .A(n_247), .Y(n_380) );
AND2x2_ASAP7_75t_L g405 ( .A(n_247), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_249), .A2(n_289), .B1(n_349), .B2(n_376), .C1(n_378), .C2(n_381), .Y(n_375) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_250), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_251), .B(n_261), .Y(n_359) );
AND2x2_ASAP7_75t_L g412 ( .A(n_251), .B(n_389), .Y(n_412) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g299 ( .A(n_257), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
INVx1_ASAP7_75t_L g314 ( .A(n_258), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_258), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_258), .B(n_432), .Y(n_456) );
OR2x6_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g417 ( .A(n_260), .B(n_406), .Y(n_417) );
INVx1_ASAP7_75t_L g440 ( .A(n_261), .Y(n_440) );
INVx1_ASAP7_75t_L g381 ( .A(n_262), .Y(n_381) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g429 ( .A(n_263), .B(n_295), .Y(n_429) );
AND2x2_ASAP7_75t_L g442 ( .A(n_263), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g283 ( .A(n_264), .Y(n_283) );
AND2x4_ASAP7_75t_L g342 ( .A(n_264), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_R g406 ( .A(n_265), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g424 ( .A(n_271), .Y(n_424) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_271), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_282), .B(n_284), .C(n_297), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g289 ( .A(n_279), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g403 ( .A(n_279), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g419 ( .A(n_280), .Y(n_419) );
BUFx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_281), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g387 ( .A(n_281), .B(n_367), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_282), .A2(n_417), .B1(n_418), .B2(n_420), .Y(n_416) );
INVx2_ASAP7_75t_L g389 ( .A(n_283), .Y(n_389) );
AND2x2_ASAP7_75t_L g445 ( .A(n_283), .B(n_367), .Y(n_445) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B(n_294), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_286), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_286), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_286), .B(n_369), .Y(n_377) );
INVx2_ASAP7_75t_L g432 ( .A(n_286), .Y(n_432) );
INVx1_ASAP7_75t_L g352 ( .A(n_287), .Y(n_352) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g409 ( .A(n_292), .Y(n_409) );
INVx2_ASAP7_75t_L g437 ( .A(n_292), .Y(n_437) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_296), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_301), .C(n_304), .Y(n_297) );
AO21x1_ASAP7_75t_L g457 ( .A1(n_298), .A2(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g418 ( .A(n_299), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g433 ( .A(n_302), .B(n_405), .Y(n_433) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_304), .A2(n_346), .B1(n_348), .B2(n_353), .Y(n_345) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_332), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_314), .B1(n_315), .B2(n_318), .C(n_322), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_311), .B(n_437), .Y(n_451) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI22xp5_ASAP7_75t_SL g322 ( .A1(n_316), .A2(n_323), .B1(n_326), .B2(n_329), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_SL g363 ( .A1(n_317), .A2(n_364), .B(n_366), .C(n_368), .Y(n_363) );
INVx2_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g325 ( .A(n_321), .Y(n_325) );
INVx1_ASAP7_75t_L g467 ( .A(n_327), .Y(n_467) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI32xp33_ASAP7_75t_L g444 ( .A1(n_328), .A2(n_370), .A3(n_387), .B1(n_445), .B2(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI211x1_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .B(n_338), .C(n_345), .Y(n_332) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_335), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_339), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g427 ( .A(n_340), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_341), .A2(n_391), .B1(n_395), .B2(n_399), .Y(n_390) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx2_ASAP7_75t_L g455 ( .A(n_342), .Y(n_455) );
INVx1_ASAP7_75t_L g468 ( .A(n_342), .Y(n_468) );
AND2x2_ASAP7_75t_L g423 ( .A(n_344), .B(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g466 ( .A(n_344), .Y(n_466) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR3x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_374), .C(n_382), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g399 ( .A(n_362), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_364), .A2(n_435), .B1(n_438), .B2(n_441), .C(n_444), .Y(n_434) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g459 ( .A(n_366), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_367), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_371), .B(n_396), .Y(n_420) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_388), .B(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_397), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g415 ( .A(n_398), .Y(n_415) );
NOR3x1_ASAP7_75t_L g400 ( .A(n_401), .B(n_421), .C(n_434), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_416), .Y(n_401) );
AOI222xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_407), .B2(n_411), .C1(n_412), .C2(n_413), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
BUFx2_ASAP7_75t_L g428 ( .A(n_410), .Y(n_428) );
NAND2xp67_ASAP7_75t_SL g436 ( .A(n_410), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g458 ( .A(n_411), .Y(n_458) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_430), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_428), .B2(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_461), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_449), .B(n_457), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B(n_456), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_458), .A2(n_462), .B1(n_465), .B2(n_471), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_694), .B1(n_712), .B2(n_713), .C(n_717), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_678), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
XOR2xp5_ASAP7_75t_L g720 ( .A(n_475), .B(n_721), .Y(n_720) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND4x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_507), .C(n_576), .D(n_666), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_493), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x4_ASAP7_75t_L g539 ( .A(n_481), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_488), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g561 ( .A(n_483), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g710 ( .A(n_483), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g540 ( .A(n_486), .B(n_514), .Y(n_540) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g513 ( .A(n_487), .B(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g575 ( .A(n_489), .Y(n_575) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g532 ( .A(n_490), .B(n_521), .Y(n_532) );
AND2x2_ASAP7_75t_L g559 ( .A(n_490), .B(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g570 ( .A(n_491), .Y(n_570) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g537 ( .A(n_492), .B(n_519), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
INVx2_ASAP7_75t_L g665 ( .A(n_494), .Y(n_665) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x6_ASAP7_75t_L g511 ( .A(n_495), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
AND2x2_ASAP7_75t_L g657 ( .A(n_498), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g627 ( .A(n_499), .B(n_628), .Y(n_627) );
OR2x6_ASAP7_75t_L g662 ( .A(n_499), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_504), .Y(n_597) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g585 ( .A(n_505), .Y(n_585) );
INVx2_ASAP7_75t_L g593 ( .A(n_505), .Y(n_593) );
INVx1_ASAP7_75t_L g602 ( .A(n_505), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_505), .B(n_506), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_505), .B(n_583), .Y(n_619) );
INVx1_ASAP7_75t_L g659 ( .A(n_505), .Y(n_659) );
INVx2_ASAP7_75t_L g583 ( .A(n_506), .Y(n_583) );
AND2x4_ASAP7_75t_L g592 ( .A(n_506), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g603 ( .A(n_506), .Y(n_603) );
INVx1_ASAP7_75t_L g634 ( .A(n_506), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_554), .C(n_564), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_515), .B1(n_538), .B2(n_541), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_SL g703 ( .A(n_513), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_522), .B1(n_523), .B2(n_527), .C(n_528), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g543 ( .A(n_517), .Y(n_543) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x2_ASAP7_75t_L g526 ( .A(n_518), .B(n_520), .Y(n_526) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_522), .A2(n_527), .B1(n_599), .B2(n_604), .C(n_608), .Y(n_598) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g547 ( .A(n_526), .Y(n_547) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g551 ( .A(n_532), .Y(n_551) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_532), .Y(n_677) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g553 ( .A(n_537), .Y(n_553) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_544), .B1(n_545), .B2(n_548), .C(n_549), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g674 ( .A(n_543), .Y(n_674) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x6_ASAP7_75t_L g671 ( .A(n_547), .B(n_669), .Y(n_671) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x6_ASAP7_75t_L g668 ( .A(n_553), .B(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g571 ( .A(n_561), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_561), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g669 ( .A(n_563), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g705 ( .A(n_568), .Y(n_705) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g711 ( .A(n_569), .Y(n_711) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI31xp33_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_594), .A3(n_629), .B(n_665), .Y(n_576) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx2_ASAP7_75t_L g589 ( .A(n_580), .Y(n_589) );
AND2x4_ASAP7_75t_L g596 ( .A(n_580), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g653 ( .A(n_581), .Y(n_653) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g663 ( .A(n_583), .Y(n_663) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
AND2x4_ASAP7_75t_L g631 ( .A(n_588), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx3_ASAP7_75t_L g625 ( .A(n_592), .Y(n_625) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_592), .Y(n_641) );
AND2x4_ASAP7_75t_L g633 ( .A(n_593), .B(n_634), .Y(n_633) );
CKINVDCx6p67_ASAP7_75t_R g595 ( .A(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_597), .Y(n_649) );
BUFx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g628 ( .A(n_601), .Y(n_628) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_620), .B1(n_621), .B2(n_626), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g638 ( .A(n_618), .Y(n_638) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx8_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_633), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .B1(n_640), .B2(n_642), .C(n_643), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_660), .B1(n_661), .B2(n_664), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
CKINVDCx11_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_672), .Y(n_666) );
OR2x2_ASAP7_75t_L g673 ( .A(n_669), .B(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g675 ( .A(n_669), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_683), .B1(n_692), .B2(n_693), .Y(n_678) );
INVx1_ASAP7_75t_L g692 ( .A(n_679), .Y(n_692) );
INVx1_ASAP7_75t_L g682 ( .A(n_680), .Y(n_682) );
INVx1_ASAP7_75t_L g693 ( .A(n_683), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_688), .Y(n_691) );
INVx1_ASAP7_75t_L g690 ( .A(n_689), .Y(n_690) );
INVx8_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OR2x6_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
OR2x4_ASAP7_75t_L g719 ( .A(n_697), .B(n_701), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_698), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g724 ( .A(n_698), .Y(n_724) );
INVx1_ASAP7_75t_L g716 ( .A(n_699), .Y(n_716) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI31xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .A3(n_706), .B(n_708), .Y(n_701) );
BUFx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx6_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
endmodule