module fake_jpeg_31234_n_513 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_513);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_513;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_8),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_94),
.Y(n_117)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_47),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_69),
.Y(n_159)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_27),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_78),
.Y(n_128)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_85),
.Y(n_122)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_30),
.B(n_7),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_101),
.Y(n_136)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_33),
.B(n_9),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_98),
.Y(n_142)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_100),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_112),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_48),
.B1(n_49),
.B2(n_35),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_107),
.A2(n_123),
.B1(n_115),
.B2(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_47),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_48),
.B1(n_39),
.B2(n_49),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_113),
.A2(n_126),
.B1(n_39),
.B2(n_18),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_115),
.A2(n_129),
.B1(n_147),
.B2(n_39),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_59),
.A2(n_26),
.B1(n_43),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_45),
.B1(n_33),
.B2(n_46),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_45),
.B1(n_33),
.B2(n_49),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_46),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_53),
.A2(n_21),
.B1(n_42),
.B2(n_37),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_20),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_100),
.B(n_20),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_32),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_100),
.B(n_20),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_160),
.B(n_168),
.Y(n_219)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g226 ( 
.A(n_164),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_54),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_165),
.B(n_172),
.Y(n_240)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_167),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_102),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_37),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_19),
.Y(n_230)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_171),
.Y(n_233)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_177),
.Y(n_224)
);

BUFx2_ASAP7_75t_SL g176 ( 
.A(n_102),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_181),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g179 ( 
.A(n_102),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_179),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_61),
.B1(n_95),
.B2(n_78),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_180),
.A2(n_205),
.B1(n_209),
.B2(n_210),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_111),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_21),
.B(n_42),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_186),
.Y(n_228)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_143),
.B1(n_147),
.B2(n_154),
.Y(n_214)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_193),
.Y(n_239)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_194),
.B(n_196),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_158),
.B1(n_149),
.B2(n_127),
.Y(n_220)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_107),
.A2(n_63),
.B1(n_96),
.B2(n_66),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_201),
.B1(n_204),
.B2(n_123),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_117),
.B(n_101),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_43),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_21),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_113),
.A2(n_87),
.B1(n_88),
.B2(n_77),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_106),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_121),
.A2(n_83),
.B1(n_67),
.B2(n_76),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_26),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_207),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_65),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_19),
.Y(n_244)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_159),
.A2(n_95),
.B1(n_28),
.B2(n_35),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_43),
.Y(n_249)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_214),
.A2(n_251),
.B1(n_254),
.B2(n_38),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_215),
.A2(n_221),
.B1(n_231),
.B2(n_236),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_222),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_110),
.B1(n_69),
.B2(n_74),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_172),
.A2(n_144),
.B1(n_156),
.B2(n_121),
.Y(n_222)
);

AOI22x1_ASAP7_75t_SL g229 ( 
.A1(n_198),
.A2(n_151),
.B1(n_127),
.B2(n_158),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_229),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_230),
.B(n_0),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_68),
.B1(n_149),
.B2(n_144),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_170),
.A2(n_26),
.B(n_18),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_235),
.A2(n_38),
.B(n_34),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_192),
.A2(n_139),
.B1(n_132),
.B2(n_153),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_166),
.B(n_162),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_238),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_24),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_139),
.B1(n_153),
.B2(n_151),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_165),
.A2(n_209),
.B1(n_185),
.B2(n_161),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_165),
.A2(n_28),
.B1(n_37),
.B2(n_24),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_163),
.B(n_35),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_196),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_263),
.Y(n_304)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_262),
.B(n_264),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_224),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_164),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_265),
.B(n_272),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_214),
.A2(n_173),
.B1(n_174),
.B2(n_182),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_267),
.A2(n_279),
.B1(n_296),
.B2(n_233),
.Y(n_326)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_213),
.C(n_169),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_282),
.C(n_293),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_202),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_273),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_252),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_276),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_229),
.A2(n_189),
.B1(n_193),
.B2(n_183),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_181),
.Y(n_276)
);

AO22x1_ASAP7_75t_SL g277 ( 
.A1(n_229),
.A2(n_220),
.B1(n_240),
.B2(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_223),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_278),
.B(n_281),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_212),
.B1(n_210),
.B2(n_205),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_219),
.B(n_167),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_171),
.C(n_19),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_19),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_223),
.B(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_228),
.B(n_19),
.Y(n_286)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_36),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_19),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_256),
.A3(n_237),
.B1(n_225),
.B2(n_239),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_252),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_292),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_226),
.B1(n_217),
.B2(n_241),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_SL g295 ( 
.A1(n_220),
.A2(n_32),
.B(n_36),
.Y(n_295)
);

AOI32xp33_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_239),
.A3(n_220),
.B1(n_237),
.B2(n_258),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_298),
.B(n_235),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_235),
.A2(n_38),
.B(n_34),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_220),
.B1(n_215),
.B2(n_221),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_300),
.A2(n_302),
.B1(n_310),
.B2(n_316),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_301),
.A2(n_307),
.B(n_273),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_323),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_247),
.B(n_256),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_308),
.A2(n_273),
.B(n_281),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_298),
.B(n_297),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_309),
.A2(n_280),
.B(n_270),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_268),
.B1(n_271),
.B2(n_277),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_243),
.B1(n_231),
.B2(n_236),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_225),
.B1(n_226),
.B2(n_258),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_319),
.A2(n_326),
.B1(n_328),
.B2(n_232),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_277),
.A2(n_250),
.B1(n_218),
.B2(n_242),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_324),
.B1(n_332),
.B2(n_335),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_234),
.C(n_245),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_329),
.C(n_32),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_247),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_271),
.A2(n_218),
.B1(n_248),
.B2(n_255),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_271),
.A2(n_234),
.B1(n_245),
.B2(n_242),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_261),
.B(n_282),
.C(n_272),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_276),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_263),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_261),
.A2(n_248),
.B1(n_233),
.B2(n_246),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_265),
.A2(n_246),
.B1(n_227),
.B2(n_258),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_306),
.A2(n_285),
.B(n_278),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_336),
.A2(n_339),
.B1(n_350),
.B2(n_312),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_337),
.A2(n_349),
.B(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_292),
.B(n_274),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_347),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_262),
.Y(n_342)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_342),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_264),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_354),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_320),
.B(n_284),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_345),
.B(n_351),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_331),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_359),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_259),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_348),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_327),
.A2(n_314),
.B1(n_330),
.B2(n_283),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_289),
.C(n_291),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_363),
.Y(n_389)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_293),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_327),
.A2(n_294),
.B1(n_296),
.B2(n_279),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_356),
.B1(n_358),
.B2(n_302),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_269),
.B1(n_260),
.B2(n_266),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_309),
.A2(n_301),
.B(n_334),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_310),
.A2(n_232),
.B(n_269),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_311),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_300),
.A2(n_227),
.B1(n_216),
.B2(n_38),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_362),
.A2(n_366),
.B1(n_315),
.B2(n_313),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_31),
.B(n_10),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_0),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_311),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_316),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_333),
.A2(n_10),
.B(n_2),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_367),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_303),
.C(n_322),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_396),
.B1(n_355),
.B2(n_356),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_374),
.C(n_379),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_303),
.C(n_325),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_376),
.B(n_388),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_325),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_384),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_318),
.C(n_315),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_381),
.A2(n_340),
.B1(n_360),
.B2(n_352),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_318),
.A3(n_333),
.B1(n_323),
.B2(n_307),
.Y(n_382)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_328),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_337),
.B(n_305),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_394),
.C(n_395),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_342),
.B(n_324),
.Y(n_393)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_332),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_348),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_340),
.A2(n_312),
.B1(n_317),
.B2(n_1),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_418)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_398),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_364),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_402),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_400),
.A2(n_403),
.B1(n_414),
.B2(n_370),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_386),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_409),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_386),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_349),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_412),
.B(n_411),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_416),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_371),
.A2(n_359),
.B1(n_358),
.B2(n_341),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_422),
.B1(n_424),
.B2(n_389),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_418),
.Y(n_431)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_366),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_373),
.B(n_345),
.C(n_317),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_423),
.C(n_394),
.Y(n_430)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_32),
.C(n_1),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_380),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_401),
.A2(n_382),
.B(n_389),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_426),
.B(n_432),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_383),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_428),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_383),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_434),
.Y(n_458)
);

AOI21xp33_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_419),
.B(n_387),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_397),
.Y(n_434)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_435),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_403),
.A2(n_381),
.B1(n_385),
.B2(n_391),
.Y(n_436)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_406),
.A2(n_385),
.B1(n_396),
.B2(n_370),
.Y(n_437)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_377),
.C(n_384),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_423),
.C(n_404),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_409),
.A2(n_414),
.B(n_422),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_407),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_410),
.B1(n_424),
.B2(n_5),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_32),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_443),
.B(n_6),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_445),
.B(n_411),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_452),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_431),
.A2(n_404),
.B1(n_400),
.B2(n_412),
.Y(n_450)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_455),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_416),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_431),
.A2(n_420),
.B(n_407),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_456),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_457),
.A2(n_459),
.B1(n_433),
.B2(n_440),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_442),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_460)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_460),
.Y(n_467)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_6),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_430),
.C(n_438),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_469),
.C(n_470),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_425),
.Y(n_465)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_465),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_471),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_434),
.C(n_445),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_428),
.C(n_443),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_429),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_454),
.A2(n_439),
.B1(n_433),
.B2(n_426),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_32),
.C(n_10),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_459),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_479),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_464),
.A2(n_446),
.B1(n_457),
.B2(n_456),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_467),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_481),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_450),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_452),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_490),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_453),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_486),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_463),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_453),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_447),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_494),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_455),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_477),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_497),
.Y(n_500)
);

AOI21xp33_ASAP7_75t_L g497 ( 
.A1(n_484),
.A2(n_476),
.B(n_474),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_487),
.A2(n_476),
.B(n_11),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_499),
.B(n_6),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_485),
.Y(n_501)
);

AO21x1_ASAP7_75t_L g507 ( 
.A1(n_501),
.A2(n_502),
.B(n_503),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_488),
.Y(n_503)
);

AOI31xp33_ASAP7_75t_L g505 ( 
.A1(n_500),
.A2(n_488),
.A3(n_490),
.B(n_492),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_505),
.B(n_501),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_504),
.A2(n_491),
.B(n_492),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_494),
.Y(n_509)
);

OAI321xp33_ASAP7_75t_L g510 ( 
.A1(n_508),
.A2(n_509),
.A3(n_507),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_6),
.B(n_12),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_14),
.B(n_16),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_512),
.A2(n_14),
.B(n_502),
.Y(n_513)
);


endmodule