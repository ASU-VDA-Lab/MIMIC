module fake_netlist_1_4380_n_27 (n_1, n_2, n_4, n_3, n_5, n_0, n_27);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
INVx1_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_4), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_1), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_0), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
NAND2xp33_ASAP7_75t_L g12 ( .A(n_6), .B(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
OR2x6_ASAP7_75t_L g15 ( .A(n_11), .B(n_7), .Y(n_15) );
BUFx4f_ASAP7_75t_SL g16 ( .A(n_13), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_14), .B(n_9), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_15), .B(n_14), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_SL g20 ( .A1(n_18), .A2(n_16), .B(n_12), .C(n_15), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_19), .B(n_15), .Y(n_21) );
NAND3xp33_ASAP7_75t_SL g22 ( .A(n_21), .B(n_10), .C(n_19), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_16), .B1(n_18), .B2(n_12), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_2), .Y(n_25) );
OAI31xp33_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_2), .A3(n_3), .B(n_5), .Y(n_26) );
AOI22xp33_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_24), .B1(n_3), .B2(n_5), .Y(n_27) );
endmodule