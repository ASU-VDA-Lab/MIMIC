module fake_jpeg_18949_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_45),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_22),
.B1(n_30),
.B2(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_54),
.A2(n_92),
.B1(n_20),
.B2(n_3),
.Y(n_133)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_58),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_75),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_16),
.Y(n_62)
);

OA22x2_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_26),
.B1(n_33),
.B2(n_19),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_29),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_68),
.Y(n_117)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_49),
.B1(n_48),
.B2(n_22),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_66),
.A2(n_70),
.B1(n_80),
.B2(n_98),
.Y(n_131)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_37),
.B1(n_17),
.B2(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_42),
.A2(n_37),
.B1(n_21),
.B2(n_32),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_21),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_38),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_41),
.B(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_95),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_44),
.A2(n_32),
.B1(n_23),
.B2(n_31),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_39),
.B(n_25),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_16),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_33),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_31),
.B1(n_24),
.B2(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_101),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_33),
.B1(n_26),
.B2(n_18),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_115),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_57),
.B1(n_70),
.B2(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_66),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g123 ( 
.A1(n_62),
.A2(n_19),
.B1(n_20),
.B2(n_4),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_124),
.B1(n_82),
.B2(n_57),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_20),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_55),
.Y(n_129)
);

CKINVDCx11_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_80),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_58),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_141),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_136),
.A2(n_106),
.B(n_67),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_139),
.B1(n_150),
.B2(n_81),
.Y(n_191)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_53),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_147),
.Y(n_175)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_78),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_78),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_71),
.A3(n_83),
.B1(n_76),
.B2(n_72),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_73),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_109),
.C(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_73),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_170),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_101),
.B1(n_84),
.B2(n_81),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_165),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_77),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_118),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

FAx1_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_120),
.CI(n_123),
.CON(n_172),
.SN(n_172)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_150),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_105),
.C(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_199),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_123),
.B1(n_83),
.B2(n_71),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_189),
.B1(n_190),
.B2(n_193),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_180),
.B(n_184),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_13),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_113),
.B1(n_130),
.B2(n_56),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_129),
.B1(n_119),
.B2(n_126),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_137),
.B1(n_140),
.B2(n_146),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_130),
.B1(n_126),
.B2(n_122),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_198),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_106),
.B1(n_127),
.B2(n_84),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_201),
.B(n_161),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_67),
.B1(n_127),
.B2(n_96),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_140),
.A2(n_1),
.B(n_4),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_143),
.A2(n_96),
.B1(n_93),
.B2(n_118),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_138),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_144),
.A2(n_10),
.B(n_14),
.Y(n_205)
);

NOR2x1_ASAP7_75t_R g233 ( 
.A(n_205),
.B(n_7),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_209),
.A2(n_216),
.B1(n_232),
.B2(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_215),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_213),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_149),
.B1(n_151),
.B2(n_163),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_220),
.B(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_157),
.C(n_158),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_230),
.C(n_196),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_233),
.B1(n_213),
.B2(n_186),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_162),
.B(n_145),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_166),
.Y(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_147),
.C(n_93),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_182),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_1),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_186),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_183),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_237),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_171),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_187),
.A3(n_171),
.B1(n_195),
.B2(n_178),
.C1(n_172),
.C2(n_193),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_229),
.C(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_182),
.B1(n_200),
.B2(n_201),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_242),
.B1(n_216),
.B2(n_218),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_227),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_203),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_255),
.C(n_256),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_248),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_210),
.B(n_173),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_251),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_172),
.C(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_172),
.C(n_180),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_210),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_228),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_259),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_212),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_217),
.B1(n_215),
.B2(n_224),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_247),
.B(n_241),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_270),
.B1(n_255),
.B2(n_243),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_257),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_273),
.C(n_240),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_211),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_234),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_208),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_189),
.B1(n_190),
.B2(n_220),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_207),
.B1(n_177),
.B2(n_233),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_248),
.Y(n_286)
);

AOI221xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_232),
.B1(n_184),
.B2(n_222),
.C(n_206),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_279),
.B1(n_264),
.B2(n_267),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_256),
.B1(n_243),
.B2(n_241),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_251),
.B(n_246),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_291),
.Y(n_299)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_231),
.B1(n_221),
.B2(n_246),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_194),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_251),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_261),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_245),
.B(n_249),
.Y(n_292)
);

OA21x2_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_275),
.B(n_272),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_303),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.Y(n_309)
);

AOI31xp33_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_221),
.A3(n_192),
.B(n_194),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_275),
.C(n_268),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_302),
.C(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_287),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_281),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_272),
.C(n_265),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_231),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_279),
.B(n_185),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_288),
.C(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_311),
.C(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_284),
.C(n_290),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_301),
.Y(n_316)
);

FAx1_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_283),
.CI(n_299),
.CON(n_310),
.SN(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_204),
.B(n_5),
.C(n_6),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_277),
.Y(n_311)
);

OAI21x1_ASAP7_75t_SL g319 ( 
.A1(n_312),
.A2(n_313),
.B(n_295),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_305),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_320),
.C(n_306),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_300),
.B(n_304),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_318),
.B(n_319),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_185),
.B(n_192),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_317),
.B(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_311),
.C(n_310),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_329),
.B(n_330),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_310),
.B(n_204),
.C(n_12),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.C(n_327),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_333),
.Y(n_334)
);


endmodule