module fake_aes_12659_n_521 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_521);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_521;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g65 ( .A(n_24), .Y(n_65) );
INVx2_ASAP7_75t_L g66 ( .A(n_13), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_43), .Y(n_67) );
CKINVDCx5p33_ASAP7_75t_R g68 ( .A(n_32), .Y(n_68) );
INVx2_ASAP7_75t_SL g69 ( .A(n_5), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_22), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_36), .Y(n_71) );
INVx2_ASAP7_75t_L g72 ( .A(n_17), .Y(n_72) );
INVx2_ASAP7_75t_L g73 ( .A(n_16), .Y(n_73) );
INVxp33_ASAP7_75t_SL g74 ( .A(n_21), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_39), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_52), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_7), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_56), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_20), .Y(n_79) );
OR2x2_ASAP7_75t_L g80 ( .A(n_26), .B(n_64), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_51), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_29), .Y(n_83) );
INVx3_ASAP7_75t_L g84 ( .A(n_47), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_10), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_0), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_60), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_11), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_42), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_49), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_40), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_12), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_28), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_41), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_9), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_55), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_34), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_84), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_84), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_69), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_91), .B(n_0), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_84), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_66), .Y(n_110) );
AND2x6_ASAP7_75t_L g111 ( .A(n_83), .B(n_30), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_103), .B(n_1), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_75), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_77), .B(n_1), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_66), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_85), .B(n_2), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_72), .B(n_2), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_88), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_100), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_98), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_98), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_73), .Y(n_125) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_85), .B(n_86), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_86), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_73), .Y(n_128) );
BUFx8_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_102), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_65), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_115), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_111), .Y(n_138) );
INVx2_ASAP7_75t_SL g139 ( .A(n_131), .Y(n_139) );
OAI21xp33_ASAP7_75t_L g140 ( .A1(n_133), .A2(n_79), .B(n_74), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_104), .B(n_99), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_107), .B(n_68), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_128), .Y(n_144) );
BUFx4_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_128), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_122), .B(n_78), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_122), .B(n_102), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_128), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_117), .B(n_101), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_115), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_131), .B(n_101), .Y(n_154) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_119), .A2(n_96), .B(n_65), .Y(n_155) );
NAND3x1_ASAP7_75t_L g156 ( .A(n_108), .B(n_96), .C(n_67), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_130), .B(n_82), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_114), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_105), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_111), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_114), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_129), .Y(n_170) );
AO22x2_ASAP7_75t_L g171 ( .A1(n_108), .A2(n_82), .B1(n_94), .B2(n_70), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_129), .B(n_81), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_105), .B(n_71), .Y(n_173) );
INVxp67_ASAP7_75t_SL g174 ( .A(n_106), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_139), .B(n_126), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_154), .B(n_111), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_139), .B(n_127), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_174), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_154), .B(n_111), .Y(n_180) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_154), .B(n_80), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_168), .B(n_112), .Y(n_182) );
AOI22xp33_ASAP7_75t_SL g183 ( .A1(n_157), .A2(n_127), .B1(n_95), .B2(n_111), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_168), .A2(n_109), .B(n_106), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_145), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_152), .B(n_135), .Y(n_186) );
NOR2x1_ASAP7_75t_L g187 ( .A(n_147), .B(n_135), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_164), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_137), .B(n_111), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_163), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_148), .B(n_110), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_143), .B(n_109), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_171), .A2(n_121), .B1(n_113), .B2(n_125), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_141), .B(n_140), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_172), .B(n_116), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_153), .B(n_113), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_158), .B(n_125), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
INVx1_ASAP7_75t_SL g205 ( .A(n_145), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_142), .A2(n_92), .B(n_70), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_155), .A2(n_121), .B1(n_132), .B2(n_134), .Y(n_210) );
CKINVDCx11_ASAP7_75t_R g211 ( .A(n_164), .Y(n_211) );
INVx5_ASAP7_75t_L g212 ( .A(n_173), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_155), .A2(n_121), .B1(n_132), .B2(n_134), .Y(n_213) );
AND2x6_ASAP7_75t_L g214 ( .A(n_149), .B(n_92), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_170), .B(n_124), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_169), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_190), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_203), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_194), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_204), .A2(n_156), .B1(n_169), .B2(n_161), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_181), .B(n_156), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_206), .B(n_155), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_216), .A2(n_123), .B1(n_71), .B2(n_76), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_206), .B(n_67), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_178), .B(n_93), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_181), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_214), .B(n_173), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_192), .B(n_76), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_215), .B(n_81), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_177), .Y(n_232) );
AOI222xp33_ASAP7_75t_L g233 ( .A1(n_211), .A2(n_89), .B1(n_90), .B2(n_94), .C1(n_173), .C2(n_134), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_214), .B(n_173), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_185), .B(n_90), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_189), .A2(n_166), .B(n_136), .Y(n_236) );
INVxp67_ASAP7_75t_L g237 ( .A(n_205), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_177), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_214), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_195), .B(n_166), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_214), .B(n_173), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_183), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_201), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_201), .Y(n_248) );
NOR2x1_ASAP7_75t_SL g249 ( .A(n_176), .B(n_89), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_244), .B(n_207), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_220), .A2(n_209), .B1(n_214), .B2(n_199), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_246), .A2(n_198), .B1(n_199), .B2(n_175), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_228), .B(n_175), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_217), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_220), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_226), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_230), .A2(n_186), .B1(n_208), .B2(n_197), .C(n_193), .Y(n_257) );
AOI222xp33_ASAP7_75t_L g258 ( .A1(n_246), .A2(n_200), .B1(n_202), .B2(n_193), .C1(n_179), .C2(n_176), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_222), .A2(n_180), .B1(n_202), .B2(n_187), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_240), .A2(n_180), .B1(n_210), .B2(n_213), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_223), .A2(n_189), .B1(n_182), .B2(n_195), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_236), .A2(n_184), .B(n_159), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_217), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_235), .B(n_201), .Y(n_265) );
OAI21x1_ASAP7_75t_SL g266 ( .A1(n_249), .A2(n_165), .B(n_136), .Y(n_266) );
OAI221xp5_ASAP7_75t_L g267 ( .A1(n_227), .A2(n_165), .B1(n_121), .B2(n_134), .C(n_151), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_224), .A2(n_146), .B(n_150), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_229), .A2(n_159), .B(n_150), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_235), .B(n_212), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_264), .B(n_235), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_252), .A2(n_239), .B1(n_225), .B2(n_231), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_254), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_252), .A2(n_239), .B1(n_218), .B2(n_243), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_258), .A2(n_245), .B(n_234), .Y(n_279) );
AOI222xp33_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_221), .B1(n_242), .B2(n_173), .C1(n_241), .C2(n_238), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_250), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g282 ( .A1(n_260), .A2(n_221), .B1(n_242), .B2(n_238), .Y(n_282) );
AOI21xp33_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_233), .B(n_241), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_260), .B(n_248), .Y(n_284) );
AO31x2_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_146), .A3(n_151), .B(n_248), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_269), .A2(n_247), .B(n_232), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_253), .A2(n_247), .B1(n_232), .B2(n_219), .C(n_162), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g289 ( .A1(n_255), .A2(n_256), .B1(n_268), .B2(n_265), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_256), .A2(n_247), .B1(n_232), .B2(n_219), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_251), .B(n_247), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_269), .A2(n_247), .B(n_232), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_287), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_273), .A2(n_268), .B1(n_257), .B2(n_265), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_278), .B(n_250), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
OAI321xp33_ASAP7_75t_L g297 ( .A1(n_277), .A2(n_259), .A3(n_267), .B1(n_261), .B2(n_262), .C(n_271), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
INVx6_ASAP7_75t_L g299 ( .A(n_284), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_272), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_281), .B(n_269), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_281), .B(n_259), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_274), .B(n_270), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_289), .B(n_271), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_283), .B(n_3), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_275), .B(n_3), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_275), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_276), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_276), .B(n_4), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_286), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_284), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_279), .B(n_4), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_282), .B(n_5), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_285), .B(n_6), .Y(n_319) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_280), .B(n_219), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_309), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_298), .B(n_291), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_303), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_314), .B(n_280), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_299), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_304), .B(n_219), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_296), .B(n_285), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_296), .B(n_285), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_308), .B(n_285), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_301), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_308), .B(n_285), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_312), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_304), .B(n_292), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_290), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_312), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_304), .B(n_6), .Y(n_339) );
AO21x2_ASAP7_75t_L g340 ( .A1(n_318), .A2(n_270), .B(n_266), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_318), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_306), .B(n_288), .C(n_160), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_312), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_304), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_302), .B(n_7), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_319), .B(n_8), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_314), .B(n_9), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_319), .B(n_10), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_307), .B(n_14), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_317), .B(n_162), .C(n_160), .Y(n_351) );
INVx5_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_300), .B(n_266), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
NAND2x1_ASAP7_75t_L g355 ( .A(n_303), .B(n_232), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_294), .B(n_219), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_316), .B(n_162), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_316), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_316), .B(n_293), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_341), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_333), .B(n_293), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_341), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_333), .B(n_307), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_348), .B(n_305), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_320), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_359), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_322), .B(n_295), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_352), .B(n_320), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_359), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_320), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_330), .B(n_311), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_330), .B(n_295), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_347), .B(n_313), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_331), .B(n_299), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_337), .B(n_310), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_349), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_349), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
NOR3xp33_ASAP7_75t_L g383 ( .A(n_346), .B(n_297), .C(n_263), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_352), .B(n_15), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_352), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_335), .Y(n_387) );
AOI322xp5_ASAP7_75t_L g388 ( .A1(n_326), .A2(n_297), .A3(n_162), .B1(n_160), .B2(n_144), .C1(n_299), .C2(n_35), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_337), .B(n_162), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_352), .Y(n_391) );
AOI33xp33_ASAP7_75t_L g392 ( .A1(n_360), .A2(n_299), .A3(n_23), .B1(n_25), .B2(n_27), .B3(n_31), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_327), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_331), .B(n_160), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_345), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_345), .B(n_160), .Y(n_396) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_342), .B(n_144), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_334), .B(n_144), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_346), .B(n_144), .C(n_212), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_353), .A2(n_144), .B1(n_212), .B2(n_38), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_352), .B(n_18), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_351), .B(n_212), .C(n_44), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_334), .B(n_37), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_354), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_327), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_352), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_338), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_367), .Y(n_409) );
AOI21xp33_ASAP7_75t_SL g410 ( .A1(n_380), .A2(n_342), .B(n_350), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_367), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_363), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_379), .B(n_360), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_380), .A2(n_332), .B1(n_350), .B2(n_360), .Y(n_416) );
NOR2xp33_ASAP7_75t_SL g417 ( .A(n_386), .B(n_344), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_373), .B(n_360), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_373), .B(n_332), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_376), .B(n_332), .Y(n_422) );
NAND4xp25_ASAP7_75t_L g423 ( .A(n_365), .B(n_351), .C(n_356), .D(n_332), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_370), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_381), .B(n_354), .Y(n_425) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_407), .A2(n_324), .B(n_336), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_368), .B(n_321), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_386), .B(n_336), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_376), .B(n_324), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_368), .B(n_323), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_386), .B(n_324), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_372), .B(n_324), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_372), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_362), .Y(n_438) );
NOR2x1_ASAP7_75t_L g439 ( .A(n_399), .B(n_397), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_407), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_387), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_377), .B(n_324), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_366), .B(n_338), .Y(n_443) );
OAI211xp5_ASAP7_75t_L g444 ( .A1(n_383), .A2(n_355), .B(n_358), .C(n_325), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_362), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_391), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_377), .B(n_325), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_364), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_375), .B(n_323), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_364), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_423), .A2(n_369), .B1(n_366), .B2(n_371), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_446), .Y(n_452) );
AOI221x1_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_401), .B1(n_385), .B2(n_402), .C(n_403), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_442), .A2(n_374), .B1(n_371), .B2(n_378), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_439), .A2(n_392), .B(n_388), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_442), .A2(n_369), .B1(n_406), .B2(n_393), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_444), .B(n_392), .C(n_403), .D(n_391), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_448), .B(n_394), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
AOI21xp33_ASAP7_75t_SL g460 ( .A1(n_426), .A2(n_385), .B(n_401), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_SL g461 ( .A1(n_420), .A2(n_394), .B(n_398), .C(n_400), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_433), .B(n_408), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_413), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_417), .A2(n_369), .B1(n_401), .B2(n_385), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_421), .A2(n_398), .B(n_389), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_416), .A2(n_408), .B1(n_404), .B2(n_389), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_446), .A2(n_396), .B(n_355), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_433), .B(n_404), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_428), .A2(n_396), .B1(n_358), .B2(n_328), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_450), .B(n_357), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_428), .A2(n_340), .B1(n_357), .B2(n_328), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_437), .B(n_340), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_447), .B(n_328), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_425), .A2(n_340), .B(n_46), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_428), .B(n_45), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_409), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_418), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_440), .A2(n_48), .B1(n_50), .B2(n_53), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_452), .B(n_419), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_451), .B(n_419), .Y(n_480) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_461), .A2(n_414), .B(n_431), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_460), .A2(n_434), .B(n_421), .C(n_443), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_455), .A2(n_430), .B(n_429), .C(n_427), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_459), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_457), .A2(n_434), .B(n_435), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_472), .B(n_445), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_463), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_475), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_476), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_477), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_470), .Y(n_491) );
NOR2xp67_ASAP7_75t_SL g492 ( .A(n_455), .B(n_435), .Y(n_492) );
OAI31xp33_ASAP7_75t_SL g493 ( .A1(n_464), .A2(n_434), .A3(n_422), .B(n_443), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_462), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_483), .A2(n_457), .B1(n_465), .B2(n_458), .C(n_438), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_481), .A2(n_454), .B1(n_467), .B2(n_471), .C(n_469), .Y(n_497) );
OAI21xp5_ASAP7_75t_SL g498 ( .A1(n_493), .A2(n_453), .B(n_475), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_491), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_473), .B(n_466), .C(n_474), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_482), .A2(n_468), .B(n_478), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_488), .B(n_432), .Y(n_502) );
OAI32xp33_ASAP7_75t_L g503 ( .A1(n_488), .A2(n_422), .A3(n_449), .B1(n_432), .B2(n_412), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_495), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_494), .B(n_409), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_496), .B(n_485), .C(n_482), .Y(n_506) );
OAI32xp33_ASAP7_75t_L g507 ( .A1(n_502), .A2(n_488), .A3(n_480), .B1(n_495), .B2(n_486), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_498), .A2(n_480), .B1(n_487), .B2(n_484), .C(n_490), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g509 ( .A1(n_501), .A2(n_489), .B(n_479), .Y(n_509) );
OAI211xp5_ASAP7_75t_L g510 ( .A1(n_497), .A2(n_479), .B(n_412), .C(n_415), .Y(n_510) );
NAND4xp75_ASAP7_75t_L g511 ( .A(n_508), .B(n_505), .C(n_499), .D(n_504), .Y(n_511) );
NOR3x2_ASAP7_75t_L g512 ( .A(n_509), .B(n_503), .C(n_500), .Y(n_512) );
NOR3x1_ASAP7_75t_L g513 ( .A(n_506), .B(n_57), .C(n_58), .Y(n_513) );
NOR3xp33_ASAP7_75t_SL g514 ( .A(n_511), .B(n_510), .C(n_507), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_512), .B(n_415), .C(n_436), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_515), .Y(n_516) );
XOR2xp5_ASAP7_75t_L g517 ( .A(n_516), .B(n_513), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_517), .A2(n_514), .B1(n_424), .B2(n_436), .Y(n_518) );
AOI222xp33_ASAP7_75t_SL g519 ( .A1(n_518), .A2(n_424), .B1(n_441), .B2(n_62), .C1(n_63), .C2(n_59), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_519), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_520), .A2(n_441), .B(n_61), .Y(n_521) );
endmodule