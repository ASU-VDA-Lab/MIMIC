module fake_jpeg_27065_n_310 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

NAND2xp67_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_23),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_50),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_19),
.C(n_26),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_37),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_39),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_29),
.C(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_60),
.B1(n_67),
.B2(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_35),
.B1(n_27),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_26),
.B1(n_17),
.B2(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_23),
.B1(n_27),
.B2(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_75),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_15),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_62),
.C(n_34),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_51),
.B1(n_41),
.B2(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_75),
.B1(n_72),
.B2(n_70),
.Y(n_106)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_95),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_8),
.Y(n_122)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_89),
.B1(n_63),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_26),
.B1(n_17),
.B2(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_14),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_53),
.B(n_20),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_18),
.B(n_14),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_20),
.B1(n_22),
.B2(n_13),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_56),
.B1(n_71),
.B2(n_20),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_108),
.B1(n_90),
.B2(n_94),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_122),
.B1(n_88),
.B2(n_86),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_88),
.B1(n_95),
.B2(n_77),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_62),
.B1(n_65),
.B2(n_69),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_115),
.C(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_100),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_84),
.B(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_33),
.C(n_31),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_33),
.C(n_31),
.Y(n_116)
);

AOI22x1_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_29),
.B1(n_13),
.B2(n_25),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_6),
.B(n_11),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_13),
.C(n_25),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_82),
.C(n_78),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_22),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_125),
.Y(n_141)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_22),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_0),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_137),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_87),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_108),
.B(n_122),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_157),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_134),
.A2(n_156),
.B(n_5),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_88),
.B1(n_78),
.B2(n_94),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_143),
.B1(n_147),
.B2(n_152),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_90),
.B1(n_81),
.B2(n_100),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_102),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_18),
.C(n_82),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_105),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_98),
.B1(n_93),
.B2(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_98),
.C(n_93),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_153),
.C(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_113),
.B(n_5),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_8),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_169),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_109),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_166),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_144),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_182),
.B1(n_158),
.B2(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_188),
.C(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_177),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_183),
.B(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx4_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_118),
.B1(n_111),
.B2(n_102),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_191),
.B1(n_160),
.B2(n_183),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_102),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_111),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_111),
.C(n_7),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_195),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_207),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_132),
.B(n_137),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_175),
.B(n_192),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_149),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_149),
.B1(n_141),
.B2(n_131),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_191),
.B1(n_184),
.B2(n_167),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_152),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_212),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_174),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_211),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_151),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_161),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_148),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_218),
.B1(n_176),
.B2(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_223),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_185),
.C(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_208),
.C(n_209),
.Y(n_239)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_180),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_181),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_229),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_177),
.B(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_196),
.B1(n_193),
.B2(n_198),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_186),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_245),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_202),
.CI(n_205),
.CON(n_243),
.SN(n_243)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_202),
.C(n_237),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_208),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_210),
.B1(n_199),
.B2(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_252),
.B1(n_238),
.B2(n_220),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_204),
.C(n_207),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_233),
.C(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_261),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_249),
.B1(n_244),
.B2(n_231),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_267),
.B1(n_262),
.B2(n_265),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_248),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_234),
.B(n_203),
.C(n_226),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_245),
.B(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_229),
.B(n_193),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_196),
.B(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_253),
.Y(n_276)
);

FAx1_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_216),
.CI(n_235),
.CON(n_265),
.SN(n_265)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_243),
.B1(n_7),
.B2(n_8),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_223),
.B1(n_167),
.B2(n_164),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_225),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_276),
.B(n_280),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_279),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_239),
.C(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_256),
.C(n_259),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_0),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_283),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_265),
.B(n_259),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_281),
.A2(n_9),
.B(n_1),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_288),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_271),
.B1(n_272),
.B2(n_4),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_0),
.C(n_1),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_2),
.C(n_3),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_2),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_2),
.B(n_3),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_3),
.Y(n_302)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_303),
.B1(n_296),
.B2(n_293),
.C(n_290),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_291),
.B(n_282),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_289),
.B(n_294),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.C(n_300),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_290),
.C(n_4),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_4),
.C(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);


endmodule