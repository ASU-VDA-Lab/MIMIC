module fake_ariane_1559_n_1782 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1782);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1782;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1759;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_45),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_17),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_89),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_52),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_13),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_1),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_69),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_2),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_107),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_41),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_29),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_151),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_123),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_0),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_3),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_21),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_33),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_55),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_60),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_83),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_25),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_32),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_56),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_3),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_11),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_41),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_47),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_43),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_68),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_104),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_9),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_82),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_105),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_140),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_57),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_24),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_99),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_84),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_50),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_101),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_81),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_98),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_44),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_59),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_73),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_154),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_64),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_4),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_33),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_37),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_58),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_46),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_47),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_10),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_14),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_130),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_40),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_20),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_27),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_36),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_110),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_29),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_112),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_21),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_62),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_120),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_46),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_78),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_65),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_137),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_49),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_124),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_31),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_15),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_17),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_80),
.Y(n_265)
);

BUFx2_ASAP7_75t_SL g266 ( 
.A(n_115),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_27),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_118),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_32),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_22),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_44),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_54),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_2),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_106),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_134),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_30),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_19),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_143),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_36),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_39),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_54),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_86),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_113),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_30),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_19),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_94),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_93),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_142),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_146),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_91),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_18),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_61),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_24),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_87),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_31),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_127),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_18),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_51),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_92),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_67),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_135),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_119),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_111),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_72),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_35),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_158),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_158),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_161),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_161),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_163),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_221),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_226),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_285),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_225),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_251),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_229),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_165),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_254),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_265),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_214),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_172),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_169),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_160),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_203),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_162),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_170),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_167),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_187),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_199),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_170),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_R g347 ( 
.A(n_190),
.B(n_152),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_190),
.B(n_5),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_291),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_219),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_243),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_262),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_168),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_197),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_173),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_170),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_258),
.B(n_5),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_174),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_177),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_188),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_291),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_201),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_202),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_205),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_204),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_204),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_264),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_282),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_207),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_216),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_211),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_234),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_211),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_235),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_217),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_185),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_236),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_217),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_284),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_214),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_224),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_258),
.B(n_6),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_237),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_238),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_224),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_378),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_313),
.A2(n_244),
.B(n_227),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_330),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_316),
.B(n_179),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_157),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_323),
.B(n_324),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_227),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_329),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_244),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_348),
.B(n_170),
.Y(n_419)
);

OR2x6_ASAP7_75t_L g420 ( 
.A(n_348),
.B(n_237),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_357),
.B(n_170),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_342),
.B(n_275),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_343),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_331),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_354),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_354),
.B(n_361),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_366),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_179),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_367),
.B(n_274),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

AND3x1_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_192),
.C(n_191),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_375),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_357),
.B(n_242),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_377),
.A2(n_279),
.B(n_275),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_380),
.B(n_383),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_344),
.A2(n_250),
.B1(n_274),
.B2(n_263),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_387),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_334),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_339),
.B(n_191),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_340),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_333),
.B(n_246),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_453),
.B(n_328),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_391),
.B(n_392),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_420),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

BUFx6f_ASAP7_75t_SL g464 ( 
.A(n_453),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g466 ( 
.A1(n_448),
.A2(n_420),
.B1(n_328),
.B2(n_451),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g468 ( 
.A1(n_451),
.A2(n_335),
.B1(n_346),
.B2(n_293),
.Y(n_468)
);

NOR2x1p5_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_359),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_420),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_453),
.B(n_454),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_349),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_420),
.A2(n_337),
.B1(n_183),
.B2(n_200),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_399),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_453),
.B(n_363),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_362),
.Y(n_483)
);

CKINVDCx6p67_ASAP7_75t_R g484 ( 
.A(n_427),
.Y(n_484)
);

BUFx4f_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_420),
.B(n_183),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_420),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_392),
.B(n_321),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_427),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_420),
.A2(n_200),
.B1(n_270),
.B2(n_280),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_399),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_453),
.B(n_364),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_L g499 ( 
.A(n_453),
.B(n_365),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_414),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_436),
.A2(n_347),
.B1(n_252),
.B2(n_273),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_453),
.B(n_370),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_434),
.A2(n_222),
.B1(n_228),
.B2(n_270),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_436),
.A2(n_271),
.B1(n_286),
.B2(n_247),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_R g511 ( 
.A(n_400),
.B(n_326),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_406),
.B(n_192),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_426),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_434),
.B(n_222),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_429),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

AND3x2_ASAP7_75t_L g524 ( 
.A(n_413),
.B(n_358),
.C(n_355),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_426),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_454),
.B(n_371),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_413),
.B(n_376),
.C(n_372),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_434),
.A2(n_280),
.B1(n_228),
.B2(n_272),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_395),
.B(n_379),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_437),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_406),
.B(n_360),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_448),
.A2(n_213),
.B1(n_239),
.B2(n_272),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_374),
.C(n_269),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_454),
.B(n_386),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_437),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_411),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_395),
.B(n_166),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_413),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_437),
.Y(n_545)
);

INVx11_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_437),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_406),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

BUFx8_ASAP7_75t_SL g551 ( 
.A(n_446),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_409),
.B(n_434),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_396),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_437),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_388),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_388),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_388),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_394),
.Y(n_558)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_434),
.B(n_178),
.Y(n_559)
);

AND2x2_ASAP7_75t_SL g560 ( 
.A(n_454),
.B(n_178),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_454),
.B(n_159),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_396),
.B(n_231),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_394),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_409),
.B(n_281),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_388),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_419),
.A2(n_196),
.B1(n_241),
.B2(n_240),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_409),
.B(n_279),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_419),
.A2(n_241),
.B1(n_240),
.B2(n_239),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_394),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_452),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_402),
.B(n_281),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_394),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_389),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_389),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_389),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_456),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_450),
.B(n_317),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_389),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_398),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_397),
.B(n_288),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_398),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_450),
.B(n_288),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_397),
.B(n_300),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_398),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_450),
.A2(n_322),
.B1(n_320),
.B2(n_327),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_398),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_403),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_402),
.B(n_193),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_401),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_403),
.Y(n_591)
);

AND2x4_ASAP7_75t_SL g592 ( 
.A(n_450),
.B(n_350),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_401),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_450),
.B(n_193),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_455),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_405),
.B(n_300),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_446),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_455),
.B(n_175),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_402),
.B(n_195),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_451),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_401),
.B(n_307),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_445),
.B(n_267),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_401),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_415),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_415),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_405),
.B(n_307),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_587),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_600),
.B(n_422),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_479),
.B(n_438),
.Y(n_609)
);

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_494),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_469),
.B(n_446),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_516),
.B(n_438),
.C(n_445),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_558),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_560),
.B(n_408),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_558),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_587),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_571),
.B(n_410),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_552),
.B(n_433),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_571),
.B(n_410),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_560),
.B(n_408),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_600),
.B(n_422),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_560),
.B(n_412),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_523),
.B(n_412),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_597),
.B(n_516),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_595),
.B(n_416),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_595),
.B(n_526),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_559),
.A2(n_421),
.B1(n_415),
.B2(n_417),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_503),
.A2(n_424),
.B1(n_407),
.B2(n_447),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_561),
.B(n_416),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_467),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_559),
.A2(n_440),
.B1(n_449),
.B2(n_447),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_494),
.B(n_351),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_564),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_559),
.B(n_418),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_549),
.B(n_418),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_551),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_539),
.B(n_407),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_523),
.B(n_423),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_549),
.B(n_423),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_473),
.B(n_440),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_544),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_552),
.B(n_433),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_523),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_553),
.B(n_425),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_553),
.B(n_425),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_473),
.B(n_428),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_527),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_565),
.B(n_433),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_484),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_511),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_552),
.B(n_473),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_520),
.B(n_538),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_527),
.B(n_428),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_589),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_552),
.B(n_430),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_565),
.B(n_456),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_604),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_SL g663 ( 
.A1(n_586),
.A2(n_352),
.B1(n_368),
.B2(n_381),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_515),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_520),
.B(n_430),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_604),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_572),
.B(n_535),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_520),
.B(n_431),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_538),
.B(n_431),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_527),
.B(n_538),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_594),
.A2(n_449),
.B1(n_444),
.B2(n_442),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_570),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_460),
.B(n_435),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_583),
.B(n_435),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_555),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_L g676 ( 
.A(n_475),
.B(n_483),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_467),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_546),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_568),
.A2(n_580),
.B(n_593),
.C(n_574),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_583),
.B(n_441),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_570),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_574),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_441),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_484),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_460),
.B(n_442),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_555),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_531),
.B(n_444),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_583),
.B(n_415),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_471),
.A2(n_487),
.B1(n_486),
.B2(n_466),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_417),
.Y(n_690)
);

AND2x6_ASAP7_75t_SL g691 ( 
.A(n_578),
.B(n_195),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_471),
.B(n_424),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_556),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_580),
.A2(n_439),
.B(n_432),
.C(n_421),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_593),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_487),
.A2(n_417),
.B1(n_421),
.B2(n_439),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_563),
.B(n_417),
.Y(n_697)
);

AOI22x1_ASAP7_75t_L g698 ( 
.A1(n_573),
.A2(n_421),
.B1(n_432),
.B2(n_439),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_536),
.A2(n_468),
.B1(n_583),
.B2(n_509),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_495),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_495),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_536),
.A2(n_439),
.B1(n_432),
.B2(n_393),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_485),
.B(n_562),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_513),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_598),
.B(n_432),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_573),
.B(n_393),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_583),
.B(n_403),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_605),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_556),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_469),
.B(n_456),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_573),
.B(n_393),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_503),
.B(n_301),
.C(n_277),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_537),
.B(n_175),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_496),
.B(n_443),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_528),
.B(n_278),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_594),
.B(n_443),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_594),
.B(n_443),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_562),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_513),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_557),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_497),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_457),
.B(n_294),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_594),
.A2(n_311),
.B1(n_289),
.B2(n_196),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_557),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_468),
.A2(n_213),
.B1(n_255),
.B2(n_260),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_566),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_535),
.B(n_369),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_490),
.B(n_281),
.Y(n_730)
);

O2A1O1Ixp5_ASAP7_75t_L g731 ( 
.A1(n_562),
.A2(n_232),
.B(n_308),
.C(n_206),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_463),
.A2(n_476),
.B(n_465),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_478),
.B(n_308),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_602),
.B(n_304),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_458),
.B(n_206),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_519),
.B(n_245),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_509),
.B(n_255),
.C(n_297),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_485),
.B(n_180),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_519),
.B(n_245),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_541),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_519),
.B(n_248),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_566),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_575),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_583),
.B(n_403),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_468),
.A2(n_289),
.B1(n_260),
.B2(n_303),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_497),
.B(n_291),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_519),
.B(n_248),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_583),
.B(n_297),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_485),
.B(n_481),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_498),
.B(n_304),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_545),
.B(n_403),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_590),
.Y(n_752)
);

BUFx5_ASAP7_75t_L g753 ( 
.A(n_463),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_590),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_486),
.A2(n_180),
.B1(n_293),
.B2(n_266),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_468),
.A2(n_299),
.B1(n_303),
.B2(n_304),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_505),
.B(n_164),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_499),
.B(n_299),
.C(n_242),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_517),
.B(n_171),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_577),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_575),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_576),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_592),
.B(n_242),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_590),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_576),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_517),
.B(n_176),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_486),
.A2(n_266),
.B1(n_310),
.B2(n_309),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_486),
.B(n_6),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_597),
.B(n_185),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_577),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_517),
.B(n_589),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_517),
.B(n_181),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_589),
.B(n_7),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_589),
.B(n_182),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_599),
.A2(n_403),
.B1(n_296),
.B2(n_298),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_579),
.Y(n_776)
);

NOR3x1_ASAP7_75t_L g777 ( 
.A(n_581),
.B(n_8),
.C(n_9),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_599),
.A2(n_242),
.B1(n_218),
.B2(n_295),
.C(n_292),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_599),
.B(n_10),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_592),
.B(n_12),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_740),
.A2(n_472),
.B(n_541),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_647),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_687),
.B(n_599),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_629),
.A2(n_464),
.B1(n_482),
.B2(n_492),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_654),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_708),
.A2(n_465),
.B(n_476),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_611),
.B(n_591),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_713),
.A2(n_510),
.B(n_512),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_684),
.B(n_584),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_687),
.B(n_641),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_613),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_667),
.B(n_590),
.Y(n_792)
);

AOI21x1_ASAP7_75t_L g793 ( 
.A1(n_718),
.A2(n_512),
.B(n_501),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_692),
.B(n_507),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_620),
.Y(n_795)
);

AOI21xp33_ASAP7_75t_L g796 ( 
.A1(n_724),
.A2(n_567),
.B(n_569),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_704),
.A2(n_488),
.B(n_491),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_656),
.B(n_590),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_647),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_704),
.A2(n_488),
.B(n_491),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_633),
.B(n_657),
.C(n_612),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_647),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_655),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_732),
.A2(n_534),
.B(n_504),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_610),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_692),
.B(n_529),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_771),
.B(n_480),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_607),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_647),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_683),
.B(n_579),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_632),
.A2(n_493),
.B(n_501),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_645),
.B(n_480),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_652),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_616),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_619),
.A2(n_493),
.B(n_504),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_652),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_730),
.B(n_480),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_621),
.A2(n_749),
.B(n_706),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_616),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_652),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_626),
.A2(n_522),
.B(n_506),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_SL g822 ( 
.A1(n_626),
.A2(n_506),
.B(n_508),
.C(n_510),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_738),
.A2(n_508),
.B(n_514),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_738),
.A2(n_514),
.B(n_522),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_653),
.B(n_582),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_661),
.B(n_524),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_631),
.B(n_582),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_719),
.A2(n_534),
.B(n_540),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_770),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_652),
.B(n_545),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_608),
.B(n_585),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_627),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_654),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_688),
.A2(n_540),
.B(n_547),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_615),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_674),
.A2(n_547),
.B(n_550),
.Y(n_836)
);

OAI321xp33_ASAP7_75t_L g837 ( 
.A1(n_756),
.A2(n_606),
.A3(n_596),
.B1(n_242),
.B2(n_603),
.C(n_585),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_680),
.A2(n_550),
.B(n_554),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_614),
.A2(n_554),
.B(n_459),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_700),
.A2(n_601),
.B1(n_603),
.B2(n_591),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_625),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_622),
.A2(n_459),
.B(n_462),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_624),
.A2(n_461),
.B(n_470),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_720),
.B(n_545),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_679),
.A2(n_502),
.B(n_461),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_628),
.A2(n_462),
.B(n_474),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_637),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_657),
.A2(n_525),
.B(n_477),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_620),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_608),
.B(n_482),
.Y(n_850)
);

AO21x2_ASAP7_75t_L g851 ( 
.A1(n_716),
.A2(n_533),
.B(n_518),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_623),
.B(n_646),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_669),
.A2(n_482),
.B(n_548),
.C(n_492),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_617),
.A2(n_525),
.B(n_477),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_617),
.A2(n_474),
.B(n_489),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_638),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_609),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_659),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_694),
.A2(n_532),
.B(n_470),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_623),
.B(n_492),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_646),
.B(n_521),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_723),
.B(n_521),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_646),
.B(n_521),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_618),
.A2(n_533),
.B(n_502),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_618),
.A2(n_543),
.B(n_518),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_644),
.A2(n_543),
.B(n_489),
.Y(n_866)
);

AOI21x1_ASAP7_75t_L g867 ( 
.A1(n_711),
.A2(n_532),
.B(n_500),
.Y(n_867)
);

NOR2x1_ASAP7_75t_L g868 ( 
.A(n_611),
.B(n_591),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_729),
.Y(n_869)
);

AOI21xp33_ASAP7_75t_L g870 ( 
.A1(n_724),
.A2(n_500),
.B(n_530),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_700),
.B(n_545),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_662),
.A2(n_530),
.B(n_548),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_727),
.A2(n_601),
.B1(n_298),
.B2(n_296),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_720),
.B(n_545),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_644),
.A2(n_548),
.B(n_530),
.C(n_218),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_678),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_646),
.B(n_601),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_760),
.B(n_588),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_778),
.B(n_249),
.C(n_198),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_646),
.B(n_601),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_651),
.B(n_601),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_651),
.A2(n_464),
.B1(n_588),
.B2(n_253),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_664),
.B(n_601),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_662),
.A2(n_464),
.B(n_259),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_682),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_666),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_678),
.B(n_601),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_665),
.B(n_186),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_730),
.A2(n_233),
.B1(n_208),
.B2(n_306),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_769),
.B(n_14),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_773),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_753),
.B(n_588),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_666),
.A2(n_668),
.B(n_665),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_753),
.B(n_671),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_668),
.A2(n_588),
.B1(n_305),
.B2(n_302),
.Y(n_895)
);

CKINVDCx16_ASAP7_75t_R g896 ( 
.A(n_636),
.Y(n_896)
);

AO21x1_ASAP7_75t_L g897 ( 
.A1(n_768),
.A2(n_157),
.B(n_230),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_660),
.B(n_189),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_663),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_689),
.A2(n_588),
.B1(n_287),
.B2(n_276),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_639),
.B(n_194),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_642),
.A2(n_256),
.B(n_209),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_643),
.B(n_212),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_676),
.B(n_215),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_699),
.B(n_634),
.Y(n_905)
);

AOI21x1_ASAP7_75t_L g906 ( 
.A1(n_728),
.A2(n_403),
.B(n_157),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_712),
.B(n_230),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_699),
.Y(n_908)
);

NAND2x1_ASAP7_75t_L g909 ( 
.A(n_754),
.B(n_403),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_658),
.A2(n_257),
.B(n_220),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_690),
.A2(n_697),
.B(n_649),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_650),
.A2(n_268),
.B(n_261),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_773),
.B(n_223),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_753),
.B(n_588),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_695),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_779),
.B(n_16),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_648),
.A2(n_230),
.B(n_157),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_779),
.B(n_16),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_733),
.B(n_20),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_672),
.A2(n_230),
.B(n_157),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_746),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_707),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_714),
.B(n_22),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_675),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_735),
.B(n_23),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_736),
.B(n_23),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_763),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_635),
.A2(n_230),
.B1(n_26),
.B2(n_28),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_725),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_768),
.A2(n_403),
.B(n_77),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_753),
.B(n_754),
.Y(n_931)
);

AND2x6_ASAP7_75t_SL g932 ( 
.A(n_712),
.B(n_34),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_681),
.A2(n_670),
.B(n_710),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_746),
.B(n_34),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_673),
.A2(n_79),
.B(n_141),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_630),
.A2(n_75),
.B(n_138),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_SL g937 ( 
.A(n_659),
.B(n_35),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_630),
.A2(n_696),
.B(n_765),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_634),
.B(n_38),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_739),
.B(n_38),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_741),
.B(n_40),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_759),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_685),
.A2(n_95),
.B(n_136),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_705),
.B(n_90),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_705),
.Y(n_945)
);

AOI21xp33_ASAP7_75t_L g946 ( 
.A1(n_734),
.A2(n_42),
.B(n_48),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_677),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_686),
.A2(n_97),
.B(n_132),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_686),
.A2(n_74),
.B(n_129),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_780),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_734),
.B(n_52),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_693),
.A2(n_103),
.B(n_128),
.Y(n_952)
);

NOR2x1p5_ASAP7_75t_SL g953 ( 
.A(n_753),
.B(n_71),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_747),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_737),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_743),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_767),
.B(n_53),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_761),
.A2(n_66),
.B(n_70),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_756),
.B(n_745),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_693),
.A2(n_108),
.B(n_117),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_722),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_722),
.A2(n_125),
.B(n_147),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_776),
.A2(n_742),
.B(n_762),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_752),
.Y(n_964)
);

CKINVDCx8_ASAP7_75t_R g965 ( 
.A(n_691),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_727),
.B(n_745),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_766),
.B(n_772),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_755),
.A2(n_748),
.B(n_731),
.C(n_774),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_857),
.B(n_712),
.Y(n_969)
);

XNOR2xp5_ASAP7_75t_L g970 ( 
.A(n_829),
.B(n_640),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_791),
.Y(n_971)
);

CKINVDCx8_ASAP7_75t_R g972 ( 
.A(n_896),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_L g973 ( 
.A1(n_951),
.A2(n_717),
.B(n_757),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_857),
.B(n_750),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_899),
.A2(n_775),
.B1(n_715),
.B2(n_726),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_893),
.A2(n_698),
.B(n_758),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_790),
.A2(n_762),
.B(n_726),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_832),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_783),
.A2(n_677),
.B(n_701),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_869),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_795),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_907),
.B(n_777),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_835),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_951),
.B(n_701),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_907),
.B(n_703),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_856),
.B(n_742),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_924),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_818),
.A2(n_807),
.B(n_881),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_782),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_858),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_891),
.A2(n_703),
.B1(n_775),
.B2(n_702),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_SL g992 ( 
.A1(n_817),
.A2(n_702),
.B(n_721),
.C(n_709),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_801),
.B(n_921),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_891),
.A2(n_721),
.B1(n_752),
.B2(n_764),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_805),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_803),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_894),
.A2(n_764),
.B(n_744),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_858),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_916),
.A2(n_918),
.B1(n_966),
.B2(n_840),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_954),
.B(n_753),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_782),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_841),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_L g1003 ( 
.A(n_876),
.B(n_751),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_847),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_894),
.A2(n_911),
.B(n_817),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_885),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_786),
.A2(n_788),
.B(n_810),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_936),
.A2(n_923),
.B(n_946),
.C(n_792),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_961),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_867),
.A2(n_963),
.B(n_828),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_915),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_856),
.B(n_959),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_782),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_852),
.B(n_806),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_808),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_795),
.B(n_849),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_923),
.A2(n_792),
.B(n_967),
.C(n_796),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_849),
.B(n_954),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_782),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_907),
.B(n_826),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_814),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_819),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_931),
.A2(n_781),
.B(n_798),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_813),
.B(n_945),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_813),
.B(n_945),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_799),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_939),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_950),
.B(n_833),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_794),
.B(n_825),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_787),
.B(n_927),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_931),
.A2(n_798),
.B(n_800),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_797),
.A2(n_834),
.B(n_811),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_807),
.A2(n_866),
.B(n_860),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_833),
.B(n_939),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_922),
.B(n_889),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_888),
.B(n_812),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_886),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_934),
.B(n_890),
.Y(n_1038)
);

OA22x2_ASAP7_75t_L g1039 ( 
.A1(n_787),
.A2(n_957),
.B1(n_928),
.B2(n_883),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_785),
.Y(n_1040)
);

INVx5_ASAP7_75t_L g1041 ( 
.A(n_787),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_929),
.A2(n_942),
.B(n_955),
.C(n_925),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_SL g1043 ( 
.A(n_937),
.B(n_913),
.C(n_812),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_789),
.B(n_799),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_868),
.B(n_887),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_901),
.A2(n_903),
.B(n_898),
.C(n_875),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_956),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_932),
.Y(n_1048)
);

NAND2x1_ASAP7_75t_L g1049 ( 
.A(n_876),
.B(n_908),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_840),
.A2(n_873),
.B1(n_827),
.B2(n_919),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_926),
.B(n_940),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_SL g1052 ( 
.A1(n_861),
.A2(n_863),
.B(n_874),
.C(n_844),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_815),
.A2(n_850),
.B(n_846),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_799),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_873),
.B(n_964),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_799),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_941),
.A2(n_938),
.B1(n_968),
.B2(n_879),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_831),
.B(n_964),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_809),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_871),
.B(n_947),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_947),
.B(n_877),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_837),
.A2(n_933),
.B(n_958),
.C(n_870),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_SL g1063 ( 
.A(n_965),
.B(n_930),
.C(n_904),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_880),
.B(n_802),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_887),
.B(n_816),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_793),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_809),
.Y(n_1067)
);

INVx5_ASAP7_75t_L g1068 ( 
.A(n_809),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_862),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_802),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_809),
.B(n_816),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_816),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_902),
.A2(n_910),
.B(n_804),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_SL g1074 ( 
.A(n_912),
.B(n_830),
.C(n_844),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_816),
.B(n_820),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_853),
.A2(n_953),
.B(n_848),
.C(n_845),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_851),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_820),
.B(n_900),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_820),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_820),
.B(n_878),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_944),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_908),
.B(n_872),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_905),
.A2(n_944),
.B1(n_830),
.B2(n_838),
.Y(n_1083)
);

OAI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_905),
.A2(n_882),
.B1(n_895),
.B2(n_909),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_SL g1085 ( 
.A1(n_874),
.A2(n_892),
.B(n_914),
.C(n_821),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_839),
.A2(n_884),
.B(n_843),
.C(n_842),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_836),
.A2(n_859),
.B1(n_784),
.B2(n_864),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_854),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_851),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_855),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_822),
.B(n_897),
.Y(n_1091)
);

BUFx10_ASAP7_75t_L g1092 ( 
.A(n_935),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_865),
.A2(n_823),
.B1(n_824),
.B2(n_892),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_914),
.B(n_917),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_943),
.A2(n_948),
.B(n_949),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_906),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_920),
.B(n_962),
.Y(n_1097)
);

BUFx8_ASAP7_75t_SL g1098 ( 
.A(n_952),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_960),
.Y(n_1099)
);

AND2x6_ASAP7_75t_SL g1100 ( 
.A(n_951),
.B(n_712),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_951),
.B(n_578),
.C(n_539),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_791),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_951),
.A2(n_790),
.B(n_946),
.C(n_783),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_783),
.A2(n_560),
.B1(n_951),
.B2(n_891),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_782),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_829),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_L g1107 ( 
.A(n_783),
.B(n_647),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_SL g1108 ( 
.A1(n_894),
.A2(n_704),
.B(n_629),
.C(n_790),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_857),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_951),
.A2(n_790),
.B(n_946),
.C(n_783),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_783),
.A2(n_560),
.B1(n_951),
.B2(n_891),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_SL g1112 ( 
.A1(n_965),
.A2(n_497),
.B1(n_586),
.B2(n_829),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_790),
.A2(n_485),
.B(n_893),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_790),
.A2(n_485),
.B(n_893),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_951),
.B(n_494),
.C(n_497),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_SL g1116 ( 
.A1(n_894),
.A2(n_704),
.B(n_629),
.C(n_790),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_783),
.A2(n_560),
.B1(n_951),
.B2(n_891),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_971),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_L g1119 ( 
.A1(n_1104),
.A2(n_1117),
.B(n_1111),
.C(n_1008),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1041),
.B(n_1065),
.Y(n_1120)
);

AOI211x1_ASAP7_75t_L g1121 ( 
.A1(n_1035),
.A2(n_1101),
.B(n_973),
.C(n_1002),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1104),
.A2(n_1117),
.B1(n_1111),
.B2(n_984),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1106),
.Y(n_1123)
);

AOI221x1_ASAP7_75t_L g1124 ( 
.A1(n_1057),
.A2(n_1017),
.B1(n_999),
.B2(n_1050),
.C(n_1073),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1018),
.B(n_1109),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1007),
.A2(n_1023),
.B(n_1031),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1068),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1093),
.A2(n_1095),
.B(n_1005),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_972),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1051),
.A2(n_1036),
.B1(n_1103),
.B2(n_1110),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1076),
.A2(n_1033),
.B(n_1077),
.Y(n_1131)
);

AOI221x1_ASAP7_75t_L g1132 ( 
.A1(n_1057),
.A2(n_999),
.B1(n_1050),
.B2(n_1063),
.C(n_1062),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1093),
.A2(n_1087),
.B(n_1094),
.Y(n_1133)
);

INVx3_ASAP7_75t_SL g1134 ( 
.A(n_995),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_991),
.A2(n_1046),
.B(n_1058),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1038),
.B(n_978),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_1089),
.A2(n_1066),
.B(n_1012),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1087),
.A2(n_1094),
.B(n_1090),
.Y(n_1138)
);

AOI221xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1042),
.A2(n_993),
.B1(n_982),
.B2(n_994),
.C(n_979),
.Y(n_1139)
);

BUFx8_ASAP7_75t_L g1140 ( 
.A(n_990),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1088),
.A2(n_988),
.B(n_1114),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_983),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1016),
.B(n_980),
.Y(n_1143)
);

AOI221x1_ASAP7_75t_L g1144 ( 
.A1(n_1091),
.A2(n_991),
.B1(n_1083),
.B2(n_1012),
.C(n_1113),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1004),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_992),
.A2(n_1082),
.B(n_1061),
.C(n_1014),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_1068),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1108),
.A2(n_1116),
.B(n_1058),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1086),
.A2(n_1082),
.B(n_1097),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_994),
.A2(n_997),
.B(n_1014),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1006),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1029),
.A2(n_1043),
.B(n_1078),
.C(n_985),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1027),
.B(n_969),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_981),
.B(n_1028),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1115),
.A2(n_1029),
.B(n_1000),
.C(n_1107),
.Y(n_1155)
);

AOI221x1_ASAP7_75t_L g1156 ( 
.A1(n_1083),
.A2(n_1060),
.B1(n_976),
.B2(n_1055),
.C(n_1081),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1099),
.A2(n_1085),
.B(n_1003),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_998),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_986),
.A2(n_1096),
.A3(n_1060),
.B(n_1064),
.Y(n_1159)
);

BUFx4_ASAP7_75t_SL g1160 ( 
.A(n_1079),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1112),
.A2(n_974),
.B1(n_1034),
.B2(n_1039),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1040),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1011),
.B(n_1102),
.Y(n_1163)
);

O2A1O1Ixp5_ASAP7_75t_L g1164 ( 
.A1(n_1084),
.A2(n_1075),
.B(n_1061),
.C(n_1064),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1068),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_986),
.A2(n_1009),
.A3(n_1037),
.B(n_1022),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1052),
.A2(n_977),
.B(n_1039),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1080),
.A2(n_1049),
.B(n_1071),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1015),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1074),
.A2(n_1047),
.B(n_975),
.C(n_1069),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_SL g1171 ( 
.A1(n_996),
.A2(n_1070),
.B1(n_1044),
.B2(n_970),
.C(n_1013),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1020),
.B(n_1100),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1021),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1065),
.B(n_1030),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1068),
.Y(n_1175)
);

AOI221x1_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_1105),
.B1(n_1026),
.B2(n_1045),
.C(n_1067),
.Y(n_1176)
);

BUFx4_ASAP7_75t_SL g1177 ( 
.A(n_1048),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1054),
.A2(n_1001),
.B(n_1013),
.Y(n_1178)
);

AO32x1_ASAP7_75t_L g1179 ( 
.A1(n_1067),
.A2(n_1072),
.A3(n_1092),
.B1(n_1098),
.B2(n_1041),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1001),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1045),
.A2(n_1092),
.B(n_1041),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1041),
.B(n_1072),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1001),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1024),
.A2(n_1025),
.B(n_1019),
.C(n_1013),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1019),
.A2(n_1056),
.B(n_1059),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1019),
.Y(n_1186)
);

AOI221xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1056),
.A2(n_951),
.B1(n_929),
.B2(n_973),
.C(n_942),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1024),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1025),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1056),
.A2(n_1005),
.B(n_1113),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1059),
.A2(n_1101),
.B1(n_951),
.B2(n_497),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_987),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1077),
.A2(n_1089),
.A3(n_1066),
.B(n_1062),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1018),
.B(n_667),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1005),
.A2(n_1114),
.B(n_1113),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1018),
.B(n_667),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_971),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_971),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1040),
.B(n_833),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1077),
.A2(n_1089),
.A3(n_1066),
.B(n_1062),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1104),
.B(n_1111),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1101),
.B(n_661),
.Y(n_1204)
);

OA22x2_ASAP7_75t_L g1205 ( 
.A1(n_1112),
.A2(n_907),
.B1(n_497),
.B2(n_509),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1104),
.A2(n_1117),
.B(n_1111),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1018),
.B(n_667),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1005),
.A2(n_1010),
.B(n_1053),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_SL g1209 ( 
.A1(n_1057),
.A2(n_946),
.B(n_1090),
.C(n_1088),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1005),
.A2(n_1114),
.B(n_1113),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1106),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_R g1212 ( 
.A(n_1043),
.B(n_655),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1005),
.A2(n_1114),
.B(n_1113),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_971),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1104),
.A2(n_1111),
.B(n_1117),
.C(n_1101),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1041),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1005),
.A2(n_1053),
.B(n_1010),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_R g1220 ( 
.A(n_990),
.B(n_494),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_981),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_987),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1077),
.A2(n_1089),
.A3(n_1066),
.B(n_1062),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1018),
.B(n_667),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1018),
.B(n_667),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_1000),
.A2(n_936),
.B(n_1104),
.Y(n_1227)
);

NOR2x1_ASAP7_75t_SL g1228 ( 
.A(n_1068),
.B(n_1041),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1068),
.Y(n_1230)
);

AOI22x1_ASAP7_75t_SL g1231 ( 
.A1(n_1048),
.A2(n_497),
.B1(n_494),
.B2(n_1106),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1077),
.A2(n_1089),
.A3(n_1066),
.B(n_1062),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1101),
.A2(n_951),
.B1(n_497),
.B2(n_511),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_987),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1101),
.A2(n_951),
.B(n_1008),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1104),
.A2(n_951),
.B(n_1111),
.C(n_1117),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_971),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1018),
.B(n_667),
.Y(n_1239)
);

CKINVDCx6p67_ASAP7_75t_R g1240 ( 
.A(n_990),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_L g1241 ( 
.A1(n_1101),
.A2(n_497),
.B1(n_503),
.B2(n_509),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1038),
.B(n_661),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1243)
);

AOI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1005),
.A2(n_1053),
.B(n_1007),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1005),
.A2(n_1114),
.B(n_1113),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_987),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1005),
.A2(n_1114),
.B(n_1113),
.Y(n_1247)
);

AO21x1_ASAP7_75t_L g1248 ( 
.A1(n_1104),
.A2(n_1117),
.B(n_1111),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1106),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_951),
.B(n_1111),
.C(n_1117),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1104),
.A2(n_1111),
.B(n_1117),
.C(n_1101),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1005),
.A2(n_1053),
.B(n_1010),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_978),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1101),
.A2(n_1111),
.B1(n_1117),
.B2(n_1104),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1109),
.B(n_857),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1104),
.A2(n_951),
.B(n_1111),
.C(n_1117),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1005),
.A2(n_1114),
.B(n_1113),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1018),
.B(n_667),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1101),
.A2(n_539),
.B(n_951),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1010),
.A2(n_1032),
.B(n_1053),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1101),
.B(n_661),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1205),
.A2(n_1206),
.B1(n_1248),
.B2(n_1204),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1138),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1123),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1147),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1140),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1183),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_1217),
.Y(n_1269)
);

CKINVDCx9p33_ASAP7_75t_R g1270 ( 
.A(n_1231),
.Y(n_1270)
);

INVx8_ASAP7_75t_L g1271 ( 
.A(n_1182),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1237),
.A2(n_1256),
.B1(n_1250),
.B2(n_1233),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1160),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1211),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1242),
.B(n_1136),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1205),
.A2(n_1262),
.B1(n_1204),
.B2(n_1203),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1262),
.A2(n_1203),
.B1(n_1254),
.B2(n_1122),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1260),
.A2(n_1132),
.B1(n_1161),
.B2(n_1124),
.Y(n_1278)
);

CKINVDCx11_ASAP7_75t_R g1279 ( 
.A(n_1240),
.Y(n_1279)
);

BUFx2_ASAP7_75t_SL g1280 ( 
.A(n_1249),
.Y(n_1280)
);

INVxp67_ASAP7_75t_SL g1281 ( 
.A(n_1149),
.Y(n_1281)
);

BUFx4f_ASAP7_75t_SL g1282 ( 
.A(n_1140),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1131),
.Y(n_1283)
);

INVx6_ASAP7_75t_L g1284 ( 
.A(n_1217),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1134),
.Y(n_1285)
);

INVx5_ASAP7_75t_L g1286 ( 
.A(n_1217),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1195),
.B(n_1197),
.Y(n_1287)
);

CKINVDCx16_ASAP7_75t_R g1288 ( 
.A(n_1129),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1130),
.A2(n_1241),
.B1(n_1236),
.B2(n_1191),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1172),
.A2(n_1226),
.B1(n_1207),
.B2(n_1258),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1135),
.A2(n_1225),
.B1(n_1239),
.B2(n_1227),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1131),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1237),
.A2(n_1256),
.B1(n_1250),
.B2(n_1215),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1163),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1215),
.A2(n_1251),
.B1(n_1152),
.B2(n_1253),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1118),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1167),
.A2(n_1154),
.B1(n_1143),
.B2(n_1119),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1134),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1251),
.A2(n_1152),
.B1(n_1253),
.B2(n_1255),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1125),
.A2(n_1144),
.B1(n_1221),
.B2(n_1212),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1142),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1145),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1160),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1158),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1133),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1162),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1221),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1167),
.A2(n_1119),
.B1(n_1153),
.B2(n_1150),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1177),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1151),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1198),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1199),
.A2(n_1214),
.B1(n_1238),
.B2(n_1174),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1173),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1153),
.A2(n_1246),
.B1(n_1169),
.B2(n_1223),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1192),
.A2(n_1234),
.B1(n_1137),
.B2(n_1181),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1177),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1212),
.A2(n_1171),
.B1(n_1187),
.B2(n_1139),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1186),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1166),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1137),
.A2(n_1181),
.B1(n_1120),
.B2(n_1149),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1220),
.Y(n_1321)
);

OAI21xp33_ASAP7_75t_L g1322 ( 
.A1(n_1170),
.A2(n_1209),
.B(n_1155),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1121),
.B(n_1170),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1166),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1200),
.A2(n_1120),
.B1(n_1188),
.B2(n_1189),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1217),
.A2(n_1180),
.B1(n_1148),
.B2(n_1182),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1228),
.A2(n_1157),
.B1(n_1148),
.B2(n_1179),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1157),
.A2(n_1175),
.B1(n_1168),
.B2(n_1147),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1175),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1168),
.A2(n_1141),
.B1(n_1127),
.B2(n_1230),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1166),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1159),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1179),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1155),
.A2(n_1165),
.B1(n_1127),
.B2(n_1230),
.Y(n_1334)
);

INVx8_ASAP7_75t_L g1335 ( 
.A(n_1165),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1185),
.A2(n_1178),
.B1(n_1210),
.B2(n_1247),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1179),
.A2(n_1164),
.B1(n_1185),
.B2(n_1128),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1185),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1178),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1213),
.B1(n_1210),
.B2(n_1245),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1164),
.A2(n_1156),
.B1(n_1213),
.B2(n_1196),
.Y(n_1341)
);

CKINVDCx6p67_ASAP7_75t_R g1342 ( 
.A(n_1184),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1184),
.Y(n_1343)
);

AOI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1146),
.A2(n_1190),
.B1(n_1252),
.B2(n_1218),
.Y(n_1344)
);

CKINVDCx12_ASAP7_75t_R g1345 ( 
.A(n_1176),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_SL g1346 ( 
.A(n_1146),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1190),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1218),
.B(n_1252),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1126),
.Y(n_1349)
);

BUFx2_ASAP7_75t_SL g1350 ( 
.A(n_1218),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1245),
.A2(n_1257),
.B1(n_1247),
.B2(n_1252),
.Y(n_1351)
);

CKINVDCx6p67_ASAP7_75t_R g1352 ( 
.A(n_1244),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1257),
.A2(n_1208),
.B(n_1193),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1208),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1194),
.A2(n_1224),
.B1(n_1232),
.B2(n_1201),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1201),
.B(n_1224),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1201),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1224),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1224),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1202),
.B(n_1216),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1219),
.A2(n_1222),
.B1(n_1229),
.B2(n_1235),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1259),
.B1(n_1261),
.B2(n_1232),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1232),
.Y(n_1363)
);

BUFx4f_ASAP7_75t_SL g1364 ( 
.A(n_1140),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1163),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1205),
.A2(n_663),
.B1(n_899),
.B2(n_320),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1237),
.A2(n_1101),
.B1(n_1256),
.B2(n_1250),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1205),
.A2(n_1206),
.B1(n_1248),
.B2(n_1262),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1163),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1205),
.A2(n_1206),
.B1(n_1248),
.B2(n_1262),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1205),
.A2(n_663),
.B1(n_899),
.B2(n_320),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1140),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1122),
.A2(n_1254),
.B1(n_1111),
.B2(n_1117),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1163),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1237),
.A2(n_1256),
.B(n_1250),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1205),
.A2(n_1206),
.B1(n_1248),
.B2(n_1262),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1205),
.A2(n_1206),
.B1(n_1248),
.B2(n_1262),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1163),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1122),
.A2(n_1254),
.B1(n_1111),
.B2(n_1117),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1195),
.B(n_1109),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1242),
.B(n_1136),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1163),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1183),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1205),
.A2(n_663),
.B1(n_899),
.B2(n_320),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1237),
.A2(n_1101),
.B1(n_1256),
.B2(n_1250),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1140),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1319),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1324),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1331),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1362),
.A2(n_1360),
.B(n_1361),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1332),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1307),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1347),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1296),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1375),
.B(n_1343),
.Y(n_1395)
);

OAI222xp33_ASAP7_75t_L g1396 ( 
.A1(n_1366),
.A2(n_1384),
.B1(n_1371),
.B2(n_1276),
.C1(n_1272),
.C2(n_1263),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1301),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1302),
.B(n_1310),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1372),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1343),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1311),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1338),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1360),
.A2(n_1361),
.B(n_1340),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1340),
.A2(n_1336),
.B(n_1344),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1353),
.A2(n_1336),
.B(n_1322),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1349),
.A2(n_1323),
.B(n_1305),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1356),
.A2(n_1281),
.B(n_1348),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1293),
.A2(n_1385),
.B1(n_1367),
.B2(n_1290),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1354),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1380),
.B(n_1294),
.Y(n_1410)
);

OAI211xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1291),
.A2(n_1277),
.B(n_1289),
.C(n_1287),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1299),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1343),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1277),
.A2(n_1278),
.B(n_1289),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1359),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1295),
.A2(n_1357),
.B1(n_1312),
.B2(n_1339),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1365),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1363),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1283),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1355),
.A2(n_1379),
.B(n_1373),
.Y(n_1420)
);

INVx4_ASAP7_75t_SL g1421 ( 
.A(n_1269),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1330),
.A2(n_1281),
.B(n_1328),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1283),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1292),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1292),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1264),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1308),
.B(n_1275),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1264),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1305),
.Y(n_1429)
);

O2A1O1Ixp5_ASAP7_75t_L g1430 ( 
.A1(n_1278),
.A2(n_1379),
.B(n_1373),
.C(n_1300),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_R g1431 ( 
.A(n_1386),
.B(n_1316),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1313),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1355),
.A2(n_1300),
.B(n_1317),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1352),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1286),
.B(n_1330),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1320),
.A2(n_1315),
.B(n_1263),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1320),
.A2(n_1315),
.B(n_1368),
.Y(n_1437)
);

INVx6_ASAP7_75t_L g1438 ( 
.A(n_1271),
.Y(n_1438)
);

BUFx4f_ASAP7_75t_SL g1439 ( 
.A(n_1298),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1369),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1381),
.B(n_1368),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1329),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1374),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1378),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1333),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1382),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1276),
.A2(n_1377),
.B1(n_1376),
.B2(n_1370),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1370),
.A2(n_1377),
.B1(n_1376),
.B2(n_1291),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1350),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1297),
.B(n_1342),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1334),
.A2(n_1325),
.B(n_1345),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1304),
.B(n_1314),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1358),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1326),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1346),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1351),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1341),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1337),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1328),
.A2(n_1266),
.B(n_1314),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1346),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1304),
.B(n_1383),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1327),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1268),
.B(n_1383),
.Y(n_1463)
);

OAI21xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1273),
.A2(n_1303),
.B(n_1285),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1284),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1268),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1439),
.B(n_1285),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1430),
.A2(n_1318),
.B(n_1306),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1409),
.B(n_1280),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1414),
.A2(n_1335),
.B(n_1271),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1417),
.B(n_1265),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1440),
.B(n_1274),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1409),
.B(n_1288),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1408),
.A2(n_1364),
.B1(n_1282),
.B2(n_1309),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1448),
.A2(n_1412),
.B(n_1411),
.C(n_1447),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1450),
.A2(n_1267),
.B(n_1270),
.Y(n_1476)
);

AND2x2_ASAP7_75t_SL g1477 ( 
.A(n_1436),
.B(n_1270),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_SL g1478 ( 
.A1(n_1396),
.A2(n_1364),
.B(n_1279),
.C(n_1321),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1435),
.B(n_1393),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1402),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1392),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_SL g1482 ( 
.A(n_1464),
.B(n_1448),
.C(n_1450),
.D(n_1427),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1395),
.A2(n_1457),
.B1(n_1416),
.B2(n_1462),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1457),
.A2(n_1458),
.B1(n_1462),
.B2(n_1433),
.C(n_1410),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1394),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1420),
.B(n_1398),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1435),
.B(n_1421),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1435),
.B(n_1421),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1404),
.A2(n_1403),
.B(n_1390),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1398),
.B(n_1407),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1392),
.B(n_1441),
.Y(n_1491)
);

AOI211xp5_ASAP7_75t_L g1492 ( 
.A1(n_1427),
.A2(n_1464),
.B(n_1458),
.C(n_1456),
.Y(n_1492)
);

INVx4_ASAP7_75t_L g1493 ( 
.A(n_1455),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1407),
.B(n_1456),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1453),
.A2(n_1454),
.B1(n_1452),
.B2(n_1432),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1433),
.A2(n_1453),
.B1(n_1437),
.B2(n_1436),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1442),
.A2(n_1413),
.B1(n_1400),
.B2(n_1466),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1443),
.B(n_1444),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1407),
.B(n_1397),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1397),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1407),
.B(n_1401),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1442),
.A2(n_1413),
.B1(n_1400),
.B2(n_1466),
.Y(n_1502)
);

AO22x2_ASAP7_75t_L g1503 ( 
.A1(n_1454),
.A2(n_1452),
.B1(n_1432),
.B2(n_1401),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1422),
.A2(n_1459),
.B(n_1449),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1405),
.B(n_1419),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1406),
.A2(n_1434),
.B(n_1460),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1460),
.A2(n_1413),
.B(n_1461),
.C(n_1405),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1405),
.B(n_1419),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1455),
.A2(n_1438),
.B1(n_1445),
.B2(n_1463),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1399),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1446),
.A2(n_1423),
.B1(n_1425),
.B2(n_1391),
.C(n_1387),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1423),
.B(n_1425),
.Y(n_1512)
);

NAND4xp25_ASAP7_75t_L g1513 ( 
.A(n_1429),
.B(n_1445),
.C(n_1428),
.D(n_1426),
.Y(n_1513)
);

AOI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1391),
.A2(n_1387),
.B1(n_1388),
.B2(n_1389),
.C(n_1424),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1451),
.A2(n_1436),
.B1(n_1437),
.B2(n_1465),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1388),
.A2(n_1389),
.B1(n_1424),
.B2(n_1415),
.C(n_1418),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1490),
.B(n_1426),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1499),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1501),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1501),
.B(n_1429),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1487),
.B(n_1402),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1449),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1505),
.B(n_1428),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1506),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1486),
.B(n_1402),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1505),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1508),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1483),
.A2(n_1437),
.B1(n_1451),
.B2(n_1418),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1508),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1494),
.B(n_1489),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1512),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1512),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1481),
.B(n_1451),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1500),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1504),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1480),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1493),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1498),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1507),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1524),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1523),
.Y(n_1542)
);

NOR2xp67_ASAP7_75t_L g1543 ( 
.A(n_1528),
.B(n_1482),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1536),
.A2(n_1515),
.B(n_1475),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1536),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1495),
.Y(n_1546)
);

INVx5_ASAP7_75t_SL g1547 ( 
.A(n_1521),
.Y(n_1547)
);

AOI33xp33_ASAP7_75t_L g1548 ( 
.A1(n_1531),
.A2(n_1478),
.A3(n_1492),
.B1(n_1484),
.B2(n_1496),
.B3(n_1473),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1525),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1523),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1523),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1526),
.B(n_1488),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1536),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1522),
.B(n_1495),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1536),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1535),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1524),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1539),
.B(n_1520),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1540),
.B(n_1473),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1522),
.B(n_1503),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1526),
.B(n_1488),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1522),
.B(n_1479),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1519),
.B(n_1524),
.Y(n_1563)
);

INVx5_ASAP7_75t_L g1564 ( 
.A(n_1537),
.Y(n_1564)
);

AND2x2_ASAP7_75t_SL g1565 ( 
.A(n_1525),
.B(n_1477),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1540),
.A2(n_1477),
.B1(n_1478),
.B2(n_1468),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1536),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1528),
.B(n_1479),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1517),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1540),
.A2(n_1475),
.B1(n_1470),
.B2(n_1474),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1520),
.B(n_1514),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1525),
.Y(n_1572)
);

NOR3xp33_ASAP7_75t_L g1573 ( 
.A(n_1534),
.B(n_1513),
.C(n_1476),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1534),
.A2(n_1516),
.B1(n_1491),
.B2(n_1469),
.C(n_1509),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1571),
.B(n_1518),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1571),
.B(n_1519),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1559),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1544),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1567),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1531),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1564),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1559),
.B(n_1431),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1546),
.B(n_1527),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.B(n_1527),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1527),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_R g1590 ( 
.A(n_1566),
.B(n_1510),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1554),
.B(n_1527),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1530),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1550),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1549),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1550),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1543),
.B(n_1538),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1551),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1568),
.B(n_1532),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1556),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1562),
.B(n_1532),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1556),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1569),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1533),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1563),
.B(n_1520),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_SL g1606 ( 
.A(n_1565),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1562),
.B(n_1533),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1590),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1597),
.B(n_1552),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1575),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1572),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1591),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1586),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1575),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1586),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1573),
.C(n_1570),
.D(n_1566),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1595),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1575),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1595),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1572),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1594),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1558),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1578),
.B(n_1558),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

NAND4xp75_ASAP7_75t_L g1627 ( 
.A(n_1597),
.B(n_1565),
.C(n_1543),
.D(n_1574),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1578),
.B(n_1431),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1581),
.A2(n_1565),
.B1(n_1544),
.B2(n_1573),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1581),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1594),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1595),
.B(n_1574),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1579),
.B(n_1552),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1606),
.A2(n_1570),
.B1(n_1565),
.B2(n_1529),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1591),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1596),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1579),
.B(n_1552),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1599),
.Y(n_1638)
);

NOR2xp67_ASAP7_75t_L g1639 ( 
.A(n_1585),
.B(n_1552),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1579),
.B(n_1552),
.Y(n_1640)
);

NOR2xp67_ASAP7_75t_L g1641 ( 
.A(n_1585),
.B(n_1561),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1581),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1581),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1598),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1605),
.B(n_1510),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1563),
.Y(n_1647)
);

INVxp33_ASAP7_75t_L g1648 ( 
.A(n_1599),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1596),
.Y(n_1649)
);

NAND4xp25_ASAP7_75t_L g1650 ( 
.A(n_1583),
.B(n_1548),
.C(n_1469),
.D(n_1467),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1611),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1633),
.B(n_1584),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1611),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1632),
.A2(n_1643),
.B(n_1617),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1627),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1615),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1633),
.B(n_1637),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1627),
.A2(n_1583),
.B(n_1577),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1620),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1618),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1609),
.B(n_1585),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1623),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1623),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1626),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1630),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1631),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1631),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1584),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1609),
.A2(n_1584),
.B(n_1577),
.C(n_1567),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1640),
.B(n_1577),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1630),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1621),
.B(n_1599),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1638),
.B(n_1601),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1614),
.B(n_1561),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1616),
.B(n_1561),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1610),
.B(n_1601),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1646),
.B(n_1604),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1622),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1619),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1685)
);

AOI21xp33_ASAP7_75t_R g1686 ( 
.A1(n_1656),
.A2(n_1641),
.B(n_1639),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1658),
.B(n_1619),
.Y(n_1687)
);

OAI21xp33_ASAP7_75t_SL g1688 ( 
.A1(n_1659),
.A2(n_1650),
.B(n_1610),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1656),
.A2(n_1629),
.B1(n_1648),
.B2(n_1634),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1656),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1651),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1655),
.B(n_1644),
.C(n_1642),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1684),
.B(n_1644),
.C(n_1642),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1662),
.A2(n_1628),
.B(n_1612),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1673),
.A2(n_1606),
.B1(n_1612),
.B2(n_1547),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1651),
.Y(n_1696)
);

OAI32xp33_ASAP7_75t_L g1697 ( 
.A1(n_1683),
.A2(n_1647),
.A3(n_1625),
.B1(n_1585),
.B2(n_1649),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1673),
.A2(n_1649),
.B(n_1544),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1653),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1653),
.Y(n_1700)
);

OAI33xp33_ASAP7_75t_L g1701 ( 
.A1(n_1677),
.A2(n_1645),
.A3(n_1613),
.B1(n_1636),
.B2(n_1635),
.B3(n_1625),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1654),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1654),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1658),
.B(n_1647),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1657),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1657),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1661),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1660),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1660),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1661),
.A2(n_1606),
.B(n_1645),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

OAI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1688),
.A2(n_1663),
.B(n_1664),
.C(n_1665),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1689),
.A2(n_1668),
.B1(n_1676),
.B2(n_1678),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1687),
.B(n_1681),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1690),
.A2(n_1606),
.B1(n_1544),
.B2(n_1676),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1687),
.B(n_1704),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1690),
.B(n_1679),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1704),
.Y(n_1718)
);

OAI31xp33_ASAP7_75t_L g1719 ( 
.A1(n_1698),
.A2(n_1676),
.A3(n_1668),
.B(n_1681),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1692),
.A2(n_1606),
.B1(n_1544),
.B2(n_1668),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1710),
.A2(n_1682),
.B(n_1664),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1710),
.A2(n_1707),
.B1(n_1694),
.B2(n_1680),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1693),
.B(n_1675),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1701),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1696),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1699),
.B(n_1675),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1674),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1718),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1727),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1714),
.B(n_1671),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1717),
.B(n_1695),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1724),
.A2(n_1685),
.B1(n_1708),
.B2(n_1706),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1723),
.B(n_1685),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1728),
.B(n_1674),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1725),
.Y(n_1738)
);

XNOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1722),
.B(n_1702),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1721),
.A2(n_1705),
.B(n_1703),
.C(n_1709),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1735),
.A2(n_1719),
.B1(n_1720),
.B2(n_1726),
.C(n_1713),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1733),
.B(n_1725),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1730),
.A2(n_1721),
.B(n_1712),
.C(n_1729),
.Y(n_1743)
);

AND3x2_ASAP7_75t_L g1744 ( 
.A(n_1738),
.B(n_1711),
.C(n_1672),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1731),
.Y(n_1745)
);

XOR2xp5_ASAP7_75t_L g1746 ( 
.A(n_1739),
.B(n_1715),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1735),
.A2(n_1734),
.B1(n_1740),
.B2(n_1712),
.Y(n_1747)
);

NOR4xp25_ASAP7_75t_L g1748 ( 
.A(n_1732),
.B(n_1663),
.C(n_1665),
.D(n_1666),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1736),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1737),
.B(n_1652),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1741),
.A2(n_1666),
.B1(n_1670),
.B2(n_1669),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1742),
.B(n_1697),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1743),
.A2(n_1669),
.B(n_1667),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1744),
.Y(n_1754)
);

OAI211xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1747),
.A2(n_1686),
.B(n_1670),
.C(n_1667),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1748),
.B(n_1746),
.Y(n_1756)
);

AOI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1754),
.A2(n_1745),
.B(n_1750),
.Y(n_1757)
);

AOI311xp33_ASAP7_75t_L g1758 ( 
.A1(n_1752),
.A2(n_1753),
.A3(n_1749),
.B(n_1751),
.C(n_1603),
.Y(n_1758)
);

AOI211xp5_ASAP7_75t_L g1759 ( 
.A1(n_1755),
.A2(n_1672),
.B(n_1652),
.C(n_1582),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1751),
.A2(n_1593),
.B1(n_1592),
.B2(n_1589),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1754),
.B(n_1582),
.C(n_1472),
.Y(n_1761)
);

XNOR2xp5_ASAP7_75t_L g1762 ( 
.A(n_1757),
.B(n_1471),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1761),
.B(n_1608),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1756),
.A2(n_1582),
.B(n_1592),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1759),
.Y(n_1765)
);

NAND4xp75_ASAP7_75t_L g1766 ( 
.A(n_1758),
.B(n_1589),
.C(n_1587),
.D(n_1588),
.Y(n_1766)
);

OAI322xp33_ASAP7_75t_L g1767 ( 
.A1(n_1765),
.A2(n_1760),
.A3(n_1582),
.B1(n_1545),
.B2(n_1567),
.C1(n_1555),
.C2(n_1553),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1762),
.B(n_1598),
.Y(n_1768)
);

NOR2x1p5_ASAP7_75t_L g1769 ( 
.A(n_1766),
.B(n_1608),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1768),
.Y(n_1770)
);

OAI22x1_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1769),
.B1(n_1763),
.B2(n_1764),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1771),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1771),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1772),
.A2(n_1767),
.B1(n_1600),
.B2(n_1598),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1773),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1775),
.B(n_1545),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1774),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1776),
.Y(n_1778)
);

AOI21xp33_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1777),
.B(n_1545),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1602),
.B1(n_1600),
.B2(n_1567),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_R g1781 ( 
.A1(n_1780),
.A2(n_1541),
.B1(n_1557),
.B2(n_1607),
.C(n_1604),
.Y(n_1781)
);

AOI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1497),
.B(n_1502),
.C(n_1545),
.Y(n_1782)
);


endmodule