module fake_jpeg_27318_n_65 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_38),
.C(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_13),
.B(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_30),
.B1(n_25),
.B2(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_10),
.B1(n_21),
.B2(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_46),
.B1(n_12),
.B2(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_23),
.B1(n_16),
.B2(n_15),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_1),
.B(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_53),
.B1(n_58),
.B2(n_57),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_59),
.B1(n_60),
.B2(n_52),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_44),
.B1(n_50),
.B2(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_44),
.B1(n_62),
.B2(n_9),
.Y(n_64)
);

OAI31xp33_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_65)
);


endmodule