module fake_jpeg_31536_n_55 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_6),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_21),
.B(n_19),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_36),
.C(n_3),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_34),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_24),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_25),
.C(n_19),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.C(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_28),
.B1(n_1),
.B2(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_18),
.B1(n_11),
.B2(n_12),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_38),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_10),
.C(n_15),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_14),
.C(n_17),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_50),
.B(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_47),
.B(n_44),
.C(n_7),
.Y(n_55)
);


endmodule