module fake_ariane_2638_n_107 (n_8, n_3, n_2, n_11, n_7, n_5, n_14, n_1, n_0, n_12, n_6, n_13, n_9, n_4, n_10, n_107);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_6;
input n_13;
input n_9;
input n_4;
input n_10;

output n_107;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_17;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_15;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_16;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVxp67_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_23),
.B(n_26),
.C(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_37),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_28),
.B(n_27),
.C(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_30),
.B(n_3),
.C(n_4),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

OAI21x1_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_47),
.B(n_49),
.Y(n_59)
);

OAI21x1_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_47),
.B(n_41),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_35),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_50),
.B1(n_33),
.B2(n_35),
.Y(n_65)
);

NOR2xp67_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_46),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_61),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_69),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_65),
.Y(n_74)
);

OR2x6_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_72),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_74),
.B1(n_80),
.B2(n_78),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_71),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_39),
.B1(n_57),
.B2(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_60),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_60),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_84),
.B1(n_83),
.B2(n_86),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_83),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_71),
.C(n_39),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_88),
.B1(n_89),
.B2(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_99),
.B1(n_98),
.B2(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_61),
.B1(n_6),
.B2(n_5),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_R g106 ( 
.A1(n_105),
.A2(n_103),
.B1(n_39),
.B2(n_5),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_61),
.B1(n_59),
.B2(n_6),
.Y(n_107)
);


endmodule