module fake_jpeg_8781_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_45),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_23),
.B1(n_26),
.B2(n_20),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_29),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_27),
.B1(n_25),
.B2(n_29),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_27),
.B1(n_25),
.B2(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_63),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_20),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_70),
.A2(n_90),
.B1(n_95),
.B2(n_97),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_52),
.B1(n_27),
.B2(n_46),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_45),
.B1(n_40),
.B2(n_25),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_44),
.B1(n_26),
.B2(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_83),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_44),
.B1(n_28),
.B2(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_86),
.B1(n_65),
.B2(n_32),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_92),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_0),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_34),
.B(n_32),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_44),
.B1(n_16),
.B2(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_31),
.B1(n_21),
.B2(n_24),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_39),
.C(n_42),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_35),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_39),
.B1(n_42),
.B2(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_113),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_118),
.B(n_115),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_115),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_35),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_125),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_93),
.B1(n_84),
.B2(n_118),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_34),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_82),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_35),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_150),
.Y(n_161)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_134),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_130),
.A2(n_21),
.B1(n_34),
.B2(n_30),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_92),
.C(n_77),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_151),
.C(n_106),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_78),
.B1(n_93),
.B2(n_68),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_142),
.B1(n_98),
.B2(n_99),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_90),
.B(n_95),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_138),
.B(n_143),
.Y(n_185)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_140),
.Y(n_190)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_84),
.B1(n_83),
.B2(n_73),
.Y(n_142)
);

BUFx12f_ASAP7_75t_SL g143 ( 
.A(n_108),
.Y(n_143)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_89),
.B1(n_24),
.B2(n_21),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_128),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_85),
.B1(n_87),
.B2(n_82),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_102),
.B1(n_98),
.B2(n_99),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_87),
.C(n_39),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_101),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_66),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_125),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_162),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_116),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_160),
.B(n_168),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_123),
.B1(n_104),
.B2(n_121),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_179),
.B1(n_140),
.B2(n_34),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_102),
.B1(n_107),
.B2(n_111),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_181),
.B1(n_191),
.B2(n_139),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_42),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_174),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_39),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_111),
.B1(n_107),
.B2(n_39),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_39),
.B1(n_32),
.B2(n_34),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_66),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_154),
.C(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_66),
.C(n_89),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_0),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_213),
.B1(n_164),
.B2(n_34),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_196),
.C(n_198),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_145),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_145),
.Y(n_198)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_209),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_144),
.B(n_137),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_216),
.B(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_126),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_183),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_139),
.B1(n_127),
.B2(n_126),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_179),
.B1(n_193),
.B2(n_169),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_217),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_33),
.B(n_30),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_159),
.B(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_9),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_166),
.B(n_158),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_233),
.B(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_226),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_162),
.B1(n_175),
.B2(n_168),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_244),
.Y(n_254)
);

XOR2x2_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_171),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_207),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_238),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_180),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_181),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_189),
.C(n_173),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_212),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_242),
.C(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_33),
.B1(n_9),
.B2(n_10),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_220),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_247),
.A2(n_264),
.B(n_14),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_251),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_192),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_192),
.C(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_195),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_198),
.C(n_197),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_201),
.B(n_208),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_8),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_8),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_227),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_276),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_246),
.B1(n_224),
.B2(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_229),
.B1(n_8),
.B2(n_11),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_275),
.B(n_284),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_15),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_265),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_14),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_267),
.Y(n_290)
);

AOI321xp33_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_11),
.A3(n_12),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_263),
.CI(n_251),
.CON(n_285),
.SN(n_285)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_284),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_286),
.B(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_279),
.C(n_271),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_255),
.C(n_248),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_295),
.C(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_254),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_248),
.C(n_254),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_11),
.C(n_12),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_279),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_300),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_274),
.B1(n_278),
.B2(n_268),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_285),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_1),
.C(n_2),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_309),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_1),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_293),
.C(n_286),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_289),
.B(n_292),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_306),
.B1(n_308),
.B2(n_299),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_291),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_2),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_320),
.A2(n_324),
.B(n_325),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_319),
.C(n_317),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_316),
.B(n_311),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_310),
.B(n_3),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_321),
.B(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_328),
.Y(n_330)
);

NAND4xp25_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_326),
.C(n_318),
.D(n_4),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_2),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_3),
.Y(n_333)
);


endmodule