module fake_aes_7617_n_30 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_SL g11 ( .A(n_3), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
BUFx6f_ASAP7_75t_SL g13 ( .A(n_0), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_0), .B(n_1), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_17), .B(n_2), .Y(n_19) );
OAI22xp5_ASAP7_75t_SL g20 ( .A1(n_14), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_20) );
AO32x2_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_13), .A3(n_17), .B1(n_11), .B2(n_12), .Y(n_21) );
CKINVDCx16_ASAP7_75t_R g22 ( .A(n_19), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
HB1xp67_ASAP7_75t_SL g24 ( .A(n_21), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_13), .B1(n_12), .B2(n_16), .Y(n_25) );
OAI321xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_12), .A3(n_18), .B1(n_24), .B2(n_21), .C(n_4), .Y(n_26) );
XOR2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_24), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_12), .B1(n_7), .B2(n_8), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
OAI222xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_5), .B1(n_7), .B2(n_9), .C1(n_24), .C2(n_28), .Y(n_30) );
endmodule