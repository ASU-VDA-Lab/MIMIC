module fake_jpeg_25981_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_6),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_72),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_56),
.B(n_62),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_54),
.B(n_57),
.C(n_61),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_59),
.C(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_46),
.Y(n_97)
);

NAND2x1_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_63),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_52),
.B1(n_68),
.B2(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_52),
.B1(n_65),
.B2(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_104),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_102),
.B1(n_60),
.B2(n_51),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_105),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_53),
.B1(n_49),
.B2(n_67),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_78),
.Y(n_103)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_1),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_98),
.B1(n_83),
.B2(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_114),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_67),
.A3(n_60),
.B1(n_51),
.B2(n_24),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_106),
.B(n_102),
.C(n_26),
.Y(n_118)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_113),
.B1(n_103),
.B2(n_27),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_126),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_1),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_2),
.B(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_135),
.B(n_130),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_139),
.B1(n_5),
.B2(n_7),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_22),
.B(n_42),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_101),
.B1(n_115),
.B2(n_5),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_3),
.B(n_4),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_21),
.C(n_41),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_127),
.C(n_17),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_143),
.C(n_141),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_151),
.A2(n_152),
.B1(n_150),
.B2(n_147),
.Y(n_153)
);

XNOR2x2_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_153),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_30),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_138),
.C(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_44),
.Y(n_159)
);

AOI321xp33_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_15),
.A3(n_38),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_14),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_29),
.Y(n_162)
);


endmodule