module real_jpeg_2585_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_1),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_26),
.C(n_31),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_2),
.B(n_29),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_42),
.C(n_46),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_2),
.B(n_101),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_54),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_55),
.C(n_57),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_2),
.B(n_48),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_3),
.A2(n_24),
.B1(n_56),
.B2(n_57),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_38),
.B1(n_56),
.B2(n_57),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_6),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_87),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_85),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_71),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_15),
.B(n_71),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_64),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_36),
.C(n_51),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_17),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_17),
.A2(n_73),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_17),
.A2(n_73),
.B1(n_147),
.B2(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_17),
.B(n_147),
.C(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B1(n_29),
.B2(n_34),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_19),
.A2(n_66),
.B(n_68),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_26),
.Y(n_28)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_21),
.B(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_25),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_31),
.B(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_34),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_51),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_48),
.B2(n_49),
.Y(n_36)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_39),
.A2(n_48),
.B1(n_108),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_40),
.A2(n_44),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22x1_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_46),
.B1(n_55),
.B2(n_60),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_46),
.B(n_231),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_48),
.A2(n_83),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_78),
.C(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_51),
.A2(n_77),
.B1(n_80),
.B2(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_63),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_61),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_61),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_53),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_53),
.A2(n_61),
.B1(n_96),
.B2(n_97),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_53),
.A2(n_61),
.B(n_97),
.Y(n_173)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_54),
.A2(n_63),
.B1(n_119),
.B2(n_146),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_54)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_57),
.B(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_66),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.C(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_72),
.A2(n_78),
.B1(n_130),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_72),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_92),
.C(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_78),
.A2(n_130),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_78),
.A2(n_129),
.B1(n_130),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_78),
.A2(n_130),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_79),
.B(n_275),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_80),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_261),
.B(n_278),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_151),
.B(n_260),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_131),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_90),
.B(n_131),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_110),
.C(n_121),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_91),
.B(n_110),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_105),
.B2(n_106),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_94),
.A2(n_95),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_94),
.A2(n_95),
.B1(n_211),
.B2(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_95),
.B(n_206),
.C(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_95),
.B(n_162),
.C(n_238),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_101),
.B1(n_126),
.B2(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_103),
.B(n_125),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_103),
.A2(n_125),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_130),
.C(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_107),
.A2(n_109),
.B1(n_173),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_107),
.A2(n_109),
.B1(n_127),
.B2(n_128),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_107),
.B(n_127),
.C(n_246),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_120),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_120),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_113),
.B(n_126),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_120),
.A2(n_135),
.B(n_142),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_121),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_129),
.C(n_130),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_122),
.A2(n_123),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_127),
.A2(n_128),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_127),
.B(n_232),
.Y(n_240)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_150),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_143),
.B2(n_144),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_134),
.B(n_143),
.C(n_150),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_147),
.B(n_149),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_147),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_181),
.C(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_165),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_149),
.A2(n_265),
.B1(n_266),
.B2(n_270),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_149),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_255),
.B(n_259),
.Y(n_151)
);

OAI211xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_184),
.B(n_198),
.C(n_199),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_174),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_166),
.B2(n_167),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_169),
.C(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_161),
.A2(n_162),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_162),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_226),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_180),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_180),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_182),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_200),
.C(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_188),
.B(n_190),
.C(n_196),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21x1_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_217),
.B(n_254),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_205),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_248),
.B(n_253),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_242),
.B(n_247),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_234),
.B(n_241),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_228),
.B(n_233),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_252),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_273),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_272),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_270),
.C(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_277),
.Y(n_280)
);


endmodule