module real_jpeg_16003_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_9),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_2),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_2),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_3),
.A2(n_184),
.B1(n_370),
.B2(n_373),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_3),
.A2(n_184),
.B1(n_190),
.B2(n_438),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_4),
.Y(n_301)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_5),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_5),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_6),
.A2(n_72),
.B1(n_77),
.B2(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_80),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_6),
.A2(n_243),
.A3(n_246),
.B1(n_247),
.B2(n_252),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_37),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_6),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_6),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_6),
.B(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_7),
.A2(n_27),
.B1(n_279),
.B2(n_283),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_7),
.A2(n_27),
.B1(n_357),
.B2(n_361),
.Y(n_356)
);

OAI22x1_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_51),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_8),
.A2(n_51),
.B1(n_210),
.B2(n_213),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_8),
.A2(n_51),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_13),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_13),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_13),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_13),
.Y(n_360)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

XOR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_463),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AO221x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_345),
.B1(n_456),
.B2(n_461),
.C(n_462),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_237),
.B(n_344),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_173),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_22),
.B(n_173),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_103),
.C(n_129),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_23),
.B(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_64),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_24),
.B(n_65),
.C(n_95),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_46),
.Y(n_24)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_25),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_25),
.A2(n_331),
.B(n_437),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_26),
.B(n_55),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_27),
.A2(n_82),
.B(n_84),
.C(n_89),
.Y(n_81)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_32),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g441 ( 
.A(n_36),
.Y(n_441)
);

NOR2x1p5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_37),
.B(n_47),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g352 ( 
.A(n_37),
.B(n_327),
.Y(n_352)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_37),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_37),
.A2(n_436),
.B(n_442),
.Y(n_435)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_42),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_56)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_46),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_55),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_55),
.Y(n_331)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_60),
.Y(n_330)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_94),
.B2(n_95),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_81),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_67),
.B(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_76),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_84),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_68),
.B(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_68),
.A2(n_180),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_74),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_79),
.Y(n_149)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_79),
.Y(n_251)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_79),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_80),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_80),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_80),
.A2(n_202),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_80),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_81),
.B(n_267),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_81),
.Y(n_381)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_88),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_89),
.A2(n_180),
.B(n_186),
.Y(n_179)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_92),
.Y(n_266)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_96),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_96),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_96),
.Y(n_450)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_96)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_103),
.A2(n_129),
.B1(n_130),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_103),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_124),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_104),
.A2(n_124),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_104),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.A3(n_111),
.B1(n_117),
.B2(n_121),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_106),
.A2(n_189),
.B1(n_193),
.B2(n_202),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_109),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_121),
.B(n_328),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_124),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_124),
.A2(n_333),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_124),
.A2(n_333),
.B1(n_449),
.B2(n_451),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_124),
.B(n_411),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B(n_128),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_125),
.A2(n_128),
.B(n_187),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_128),
.A2(n_264),
.B(n_267),
.Y(n_263)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_154),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_132),
.B(n_321),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_134),
.A2(n_143),
.B(n_155),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_134),
.B(n_155),
.Y(n_261)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_141),
.Y(n_375)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_142),
.Y(n_307)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_143),
.B(n_169),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_143),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_154),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_169),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_155),
.B(n_278),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_155),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_162),
.B2(n_166),
.Y(n_156)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_158),
.Y(n_372)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_205),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_175),
.B(n_178),
.C(n_205),
.Y(n_398)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_179),
.B(n_188),
.Y(n_350)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_186),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_230),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_206),
.B(n_231),
.C(n_234),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_207),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_208),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_209),
.B(n_217),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_209),
.Y(n_420)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_214),
.Y(n_362)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_216),
.B(n_355),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_227),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_217),
.B(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_217),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_224),
.B2(n_226),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_227),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_231),
.A2(n_232),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_235),
.B(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_236),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_338),
.B(n_343),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_315),
.B(n_337),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_290),
.B(n_314),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_262),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_241),
.B(n_262),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_259),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_242),
.B(n_259),
.Y(n_312)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

NAND2xp67_ASAP7_75t_L g379 ( 
.A(n_261),
.B(n_277),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_275),
.Y(n_262)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_268),
.Y(n_303)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_277),
.A2(n_412),
.B(n_413),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_288),
.C(n_336),
.Y(n_335)
);

OAI21x1_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_309),
.B(n_313),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_304),
.B(n_308),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_335),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_335),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_332),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_323),
.C(n_332),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_321),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_325),
.B(n_418),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g384 ( 
.A1(n_326),
.A2(n_331),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_333),
.A2(n_449),
.B(n_453),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_342),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_401),
.C(n_425),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_397),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_347),
.B(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_389),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_348),
.B(n_389),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_364),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_365),
.C(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.C(n_353),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_351),
.A2(n_353),
.B1(n_354),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_363),
.Y(n_354)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_377),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_366),
.A2(n_368),
.B(n_376),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_376),
.Y(n_367)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_382),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_380),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_386),
.B2(n_388),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_406),
.C(n_407),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.C(n_396),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_400),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_396),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_398),
.B(n_399),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_401),
.A2(n_457),
.B(n_458),
.C(n_460),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_404),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_414),
.B1(n_423),
.B2(n_424),
.Y(n_408)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_427),
.C(n_428),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_414),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_431),
.C(n_432),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_421),
.A2(n_422),
.B(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_424),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_425),
.Y(n_461)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_429),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_430),
.B(n_434),
.C(n_479),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_446),
.B1(n_454),
.B2(n_455),
.Y(n_433)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_443),
.B(n_445),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_444),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_445),
.A2(n_468),
.B1(n_469),
.B2(n_476),
.Y(n_467)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_446),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_452),
.B2(n_453),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_449),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_452),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_480),
.Y(n_463)
);

INVxp33_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_478),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_478),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_477),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_474),
.B2(n_475),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_472),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);


endmodule