module fake_jpeg_26780_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_20),
.B(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_6),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_17),
.B1(n_14),
.B2(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_28),
.B(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_46),
.B(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_56),
.B1(n_35),
.B2(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_29),
.B(n_26),
.C(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_69),
.Y(n_72)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_56),
.B1(n_53),
.B2(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_68),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_49),
.C(n_33),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_58),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_62),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_85),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_55),
.B1(n_56),
.B2(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_56),
.B1(n_46),
.B2(n_37),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_45),
.B(n_33),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_45),
.B(n_21),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_51),
.B1(n_43),
.B2(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_68),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_97),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_67),
.A3(n_63),
.B1(n_57),
.B2(n_58),
.C1(n_62),
.C2(n_59),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_19),
.A3(n_15),
.B1(n_16),
.B2(n_12),
.C1(n_29),
.C2(n_26),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_96),
.B1(n_84),
.B2(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_64),
.B1(n_66),
.B2(n_35),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_80),
.B(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_106),
.B1(n_98),
.B2(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_76),
.B1(n_74),
.B2(n_83),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_86),
.C(n_97),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_107),
.C(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_83),
.B1(n_22),
.B2(n_20),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_5),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_22),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_125),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_65),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_111),
.C(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_124),
.C(n_26),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_98),
.C(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_83),
.B1(n_64),
.B2(n_51),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_70),
.B1(n_59),
.B2(n_34),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.C(n_65),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_15),
.B(n_16),
.C(n_12),
.D(n_24),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_37),
.B1(n_42),
.B2(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_16),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_115),
.B1(n_116),
.B2(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_137),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_65),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_29),
.C(n_24),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_116),
.C(n_42),
.Y(n_142)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_65),
.B1(n_15),
.B2(n_12),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_31),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_128),
.C(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_148),
.Y(n_157)
);

NAND4xp25_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_65),
.C(n_7),
.D(n_8),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_136),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_15),
.C(n_5),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_156),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_133),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_4),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_7),
.B(n_9),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_11),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_8),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_175),
.B(n_170),
.C(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_162),
.A3(n_11),
.B1(n_2),
.B2(n_3),
.C1(n_1),
.C2(n_0),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_3),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_0),
.C(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_3),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_3),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_184),
.Y(n_186)
);


endmodule