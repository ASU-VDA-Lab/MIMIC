module real_aes_15974_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g103 ( .A(n_0), .B(n_104), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_1), .A2(n_4), .B1(n_274), .B2(n_275), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_2), .A2(n_43), .B1(n_175), .B2(n_223), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_3), .A2(n_24), .B1(n_223), .B2(n_257), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_5), .A2(n_16), .B1(n_523), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_6), .A2(n_61), .B1(n_160), .B2(n_161), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_7), .A2(n_17), .B1(n_175), .B2(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g104 ( .A(n_8), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_9), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_10), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_11), .A2(n_18), .B1(n_524), .B2(n_568), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_12), .A2(n_65), .B1(n_133), .B2(n_134), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
OR2x2_ASAP7_75t_L g110 ( .A(n_13), .B(n_38), .Y(n_110) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_14), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_15), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_19), .A2(n_99), .B1(n_275), .B2(n_523), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_20), .A2(n_39), .B1(n_153), .B2(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_21), .B(n_151), .Y(n_584) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_22), .A2(n_59), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_23), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_25), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_26), .B(n_148), .Y(n_215) );
INVx4_ASAP7_75t_R g199 ( .A(n_27), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_28), .A2(n_47), .B1(n_179), .B2(n_272), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_29), .A2(n_54), .B1(n_179), .B2(n_523), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_30), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_31), .B(n_548), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_32), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_33), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g279 ( .A(n_34), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_SL g254 ( .A1(n_35), .A2(n_147), .B(n_175), .C(n_255), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_36), .A2(n_55), .B1(n_175), .B2(n_179), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_37), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_40), .A2(n_87), .B1(n_175), .B2(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g817 ( .A1(n_41), .A2(n_53), .B1(n_818), .B2(n_819), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_41), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_42), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_44), .A2(n_46), .B1(n_175), .B2(n_176), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_45), .A2(n_60), .B1(n_523), .B2(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g219 ( .A(n_48), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_49), .B(n_175), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_50), .Y(n_233) );
INVx2_ASAP7_75t_L g128 ( .A(n_51), .Y(n_128) );
BUFx3_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g122 ( .A(n_52), .Y(n_122) );
INVx1_ASAP7_75t_L g818 ( .A(n_53), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_56), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_57), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_58), .A2(n_88), .B1(n_175), .B2(n_179), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_62), .A2(n_75), .B1(n_272), .B2(n_540), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_63), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_64), .A2(n_79), .B1(n_175), .B2(n_176), .Y(n_525) );
INVx1_ASAP7_75t_L g134 ( .A(n_65), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_66), .A2(n_98), .B1(n_523), .B2(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g166 ( .A(n_67), .Y(n_166) );
AND2x4_ASAP7_75t_L g169 ( .A(n_68), .B(n_170), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_69), .A2(n_90), .B1(n_179), .B2(n_272), .Y(n_271) );
AO22x1_ASAP7_75t_L g149 ( .A1(n_70), .A2(n_76), .B1(n_150), .B2(n_153), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_71), .Y(n_170) );
AND2x2_ASAP7_75t_L g258 ( .A(n_72), .B(n_211), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_73), .B(n_160), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_74), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_77), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_78), .B(n_223), .Y(n_234) );
INVx2_ASAP7_75t_L g148 ( .A(n_80), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_81), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_82), .B(n_211), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_83), .A2(n_97), .B1(n_160), .B2(n_179), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_84), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_85), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_86), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_89), .B(n_211), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_91), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_92), .B(n_211), .Y(n_230) );
INVx1_ASAP7_75t_L g107 ( .A(n_93), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_93), .B(n_121), .Y(n_120) );
NAND2xp33_ASAP7_75t_L g587 ( .A(n_94), .B(n_151), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_95), .A2(n_160), .B(n_181), .C(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g204 ( .A(n_96), .B(n_205), .Y(n_204) );
NAND2xp33_ASAP7_75t_L g238 ( .A(n_100), .B(n_200), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_111), .B(n_820), .Y(n_101) );
BUFx8_ASAP7_75t_L g822 ( .A(n_102), .Y(n_822) );
AND2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
INVx1_ASAP7_75t_L g805 ( .A(n_105), .Y(n_805) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_106), .Y(n_495) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g130 ( .A(n_109), .Y(n_130) );
INVx1_ASAP7_75t_L g123 ( .A(n_110), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_806), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_124), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_114), .A2(n_812), .B(n_814), .Y(n_811) );
NOR2x1_ASAP7_75t_R g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g813 ( .A(n_117), .Y(n_813) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
CKINVDCx8_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_123), .B(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_131), .B(n_800), .Y(n_124) );
BUFx12f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_128), .B(n_805), .Y(n_804) );
INVx3_ASAP7_75t_L g810 ( .A(n_128), .Y(n_810) );
OAI22xp33_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_135), .B1(n_136), .B2(n_799), .Y(n_131) );
INVx1_ASAP7_75t_L g799 ( .A(n_132), .Y(n_799) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI22x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_494), .B1(n_496), .B2(n_798), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_404), .Y(n_138) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_333), .C(n_375), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_307), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_206), .B1(n_282), .B2(n_293), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_187), .Y(n_143) );
AOI21xp33_ASAP7_75t_L g326 ( .A1(n_144), .A2(n_327), .B(n_329), .Y(n_326) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_144), .A2(n_400), .B(n_401), .Y(n_399) );
OR2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_171), .Y(n_144) );
INVx2_ASAP7_75t_L g319 ( .A(n_145), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_145), .B(n_172), .Y(n_349) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_155), .C(n_167), .Y(n_146) );
INVx6_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_147), .A2(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_147), .B(n_149), .Y(n_291) );
O2A1O1Ixp5_ASAP7_75t_L g582 ( .A1(n_147), .A2(n_176), .B(n_583), .C(n_584), .Y(n_582) );
BUFx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
INVx1_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
INVx1_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
INVxp67_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g523 ( .A(n_151), .Y(n_523) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g154 ( .A(n_152), .Y(n_154) );
INVx1_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx3_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_152), .Y(n_223) );
INVx1_ASAP7_75t_L g251 ( .A(n_152), .Y(n_251) );
INVx2_ASAP7_75t_L g257 ( .A(n_152), .Y(n_257) );
OAI21xp33_ASAP7_75t_SL g214 ( .A1(n_153), .A2(n_215), .B(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g290 ( .A(n_155), .Y(n_290) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_163), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_156), .A2(n_221), .B(n_222), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_156), .A2(n_177), .B1(n_262), .B2(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g506 ( .A(n_157), .Y(n_506) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
INVx1_ASAP7_75t_L g568 ( .A(n_161), .Y(n_568) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_162), .B(n_196), .Y(n_195) );
OAI21xp33_ASAP7_75t_L g167 ( .A1(n_163), .A2(n_164), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g182 ( .A(n_164), .Y(n_182) );
INVx2_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
INVx2_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
INVx1_ASAP7_75t_L g292 ( .A(n_167), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_168), .A2(n_247), .B(n_254), .Y(n_246) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx10_ASAP7_75t_L g183 ( .A(n_169), .Y(n_183) );
BUFx10_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
INVx1_ASAP7_75t_L g277 ( .A(n_169), .Y(n_277) );
AND2x2_ASAP7_75t_L g389 ( .A(n_171), .B(n_228), .Y(n_389) );
INVx1_ASAP7_75t_L g422 ( .A(n_171), .Y(n_422) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g284 ( .A(n_172), .B(n_229), .Y(n_284) );
AND2x2_ASAP7_75t_L g315 ( .A(n_172), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g324 ( .A(n_172), .Y(n_324) );
OR2x2_ASAP7_75t_L g343 ( .A(n_172), .B(n_189), .Y(n_343) );
AND2x2_ASAP7_75t_L g358 ( .A(n_172), .B(n_189), .Y(n_358) );
AO31x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_182), .A3(n_183), .B(n_184), .Y(n_172) );
OAI22x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B1(n_178), .B2(n_180), .Y(n_173) );
INVx4_ASAP7_75t_L g176 ( .A(n_175), .Y(n_176) );
INVx1_ASAP7_75t_L g524 ( .A(n_175), .Y(n_524) );
INVx1_ASAP7_75t_L g540 ( .A(n_175), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_176), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_177), .A2(n_180), .B1(n_271), .B2(n_273), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_177), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_177), .A2(n_180), .B1(n_514), .B2(n_516), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_177), .A2(n_522), .B1(n_525), .B2(n_526), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_177), .A2(n_506), .B1(n_538), .B2(n_539), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_177), .A2(n_506), .B1(n_547), .B2(n_549), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_177), .A2(n_506), .B1(n_557), .B2(n_558), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_177), .A2(n_526), .B1(n_567), .B2(n_569), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_177), .A2(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_179), .B(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_180), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_SL g526 ( .A(n_181), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_182), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_182), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g203 ( .A(n_183), .Y(n_203) );
AO31x2_ASAP7_75t_L g503 ( .A1(n_183), .A2(n_264), .A3(n_504), .B(n_508), .Y(n_503) );
AO31x2_ASAP7_75t_L g545 ( .A1(n_183), .A2(n_512), .A3(n_546), .B(n_551), .Y(n_545) );
AO31x2_ASAP7_75t_L g565 ( .A1(n_183), .A2(n_245), .A3(n_566), .B(n_570), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx2_ASAP7_75t_L g205 ( .A(n_186), .Y(n_205) );
BUFx2_ASAP7_75t_L g245 ( .A(n_186), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_186), .B(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_186), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_188), .B(n_357), .Y(n_400) );
OR2x2_ASAP7_75t_L g488 ( .A(n_188), .B(n_349), .Y(n_488) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g316 ( .A(n_189), .Y(n_316) );
AND2x2_ASAP7_75t_L g325 ( .A(n_189), .B(n_288), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_189), .B(n_229), .Y(n_328) );
AND2x2_ASAP7_75t_L g347 ( .A(n_189), .B(n_228), .Y(n_347) );
AND2x4_ASAP7_75t_L g366 ( .A(n_189), .B(n_289), .Y(n_366) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_193), .B(n_204), .Y(n_189) );
AO31x2_ASAP7_75t_L g536 ( .A1(n_190), .A2(n_527), .A3(n_537), .B(n_541), .Y(n_536) );
AO31x2_ASAP7_75t_L g555 ( .A1(n_190), .A2(n_276), .A3(n_556), .B(n_559), .Y(n_555) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_192), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_SL g570 ( .A(n_192), .B(n_571), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_197), .B(n_203), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g272 ( .A(n_200), .Y(n_272) );
INVx1_ASAP7_75t_L g548 ( .A(n_200), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_201), .Y(n_550) );
INVx1_ASAP7_75t_L g527 ( .A(n_203), .Y(n_527) );
OAI21xp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_226), .B(n_267), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_207), .B(n_361), .Y(n_464) );
CKINVDCx14_ASAP7_75t_R g207 ( .A(n_208), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_209), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g297 ( .A(n_209), .Y(n_297) );
OR2x2_ASAP7_75t_L g305 ( .A(n_209), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_209), .B(n_298), .Y(n_330) );
AND2x2_ASAP7_75t_L g355 ( .A(n_209), .B(n_269), .Y(n_355) );
AND2x2_ASAP7_75t_L g373 ( .A(n_209), .B(n_303), .Y(n_373) );
INVx1_ASAP7_75t_L g412 ( .A(n_209), .Y(n_412) );
AND2x2_ASAP7_75t_L g414 ( .A(n_209), .B(n_415), .Y(n_414) );
NAND2x1p5_ASAP7_75t_SL g433 ( .A(n_209), .B(n_354), .Y(n_433) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_213), .Y(n_209) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_211), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g264 ( .A(n_211), .Y(n_264) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g224 ( .A(n_212), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_212), .B(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g512 ( .A(n_212), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_212), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_212), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g580 ( .A(n_212), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_224), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
BUFx4f_ASAP7_75t_L g253 ( .A(n_218), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_223), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g241 ( .A(n_225), .Y(n_241) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_225), .A2(n_261), .A3(n_264), .B(n_265), .Y(n_260) );
OAI32xp33_ASAP7_75t_L g317 ( .A1(n_226), .A2(n_309), .A3(n_318), .B1(n_320), .B2(n_322), .Y(n_317) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_242), .Y(n_226) );
INVx1_ASAP7_75t_L g357 ( .A(n_227), .Y(n_357) );
AND2x2_ASAP7_75t_L g365 ( .A(n_227), .B(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g364 ( .A(n_228), .B(n_288), .Y(n_364) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx3_ASAP7_75t_L g314 ( .A(n_229), .Y(n_314) );
AND2x2_ASAP7_75t_L g323 ( .A(n_229), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g429 ( .A(n_229), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_237), .B(n_240), .Y(n_231) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g299 ( .A(n_242), .Y(n_299) );
OR2x2_ASAP7_75t_L g309 ( .A(n_242), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g431 ( .A(n_242), .Y(n_431) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_259), .Y(n_242) );
AND2x2_ASAP7_75t_L g332 ( .A(n_243), .B(n_260), .Y(n_332) );
INVx2_ASAP7_75t_L g354 ( .A(n_243), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_243), .B(n_269), .Y(n_374) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g281 ( .A(n_244), .Y(n_281) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_258), .Y(n_244) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_270), .A3(n_276), .B(n_278), .Y(n_269) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_245), .A2(n_521), .A3(n_527), .B(n_528), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B(n_253), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g275 ( .A(n_251), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_SL g515 ( .A(n_257), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_259), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g363 ( .A(n_259), .Y(n_363) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
OR2x2_ASAP7_75t_L g369 ( .A(n_260), .B(n_269), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_260), .B(n_269), .Y(n_402) );
INVx2_ASAP7_75t_L g350 ( .A(n_267), .Y(n_350) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_280), .Y(n_267) );
OR2x2_ASAP7_75t_L g337 ( .A(n_268), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g415 ( .A(n_268), .Y(n_415) );
INVx1_ASAP7_75t_L g298 ( .A(n_269), .Y(n_298) );
INVx1_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
INVx1_ASAP7_75t_L g321 ( .A(n_269), .Y(n_321) );
AO31x2_ASAP7_75t_L g511 ( .A1(n_276), .A2(n_512), .A3(n_513), .B(n_517), .Y(n_511) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_SL g588 ( .A(n_277), .Y(n_588) );
OR2x2_ASAP7_75t_L g425 ( .A(n_280), .B(n_402), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_281), .B(n_297), .Y(n_338) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
OR2x2_ASAP7_75t_L g439 ( .A(n_281), .B(n_363), .Y(n_439) );
INVxp67_ASAP7_75t_L g463 ( .A(n_281), .Y(n_463) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
NAND2x1_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_284), .B(n_325), .Y(n_392) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g341 ( .A(n_286), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g454 ( .A(n_287), .Y(n_454) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g483 ( .A(n_288), .B(n_316), .Y(n_483) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g409 ( .A(n_289), .B(n_316), .Y(n_409) );
AOI21x1_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_292), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_300), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_296), .B(n_332), .Y(n_446) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g310 ( .A(n_297), .Y(n_310) );
AND2x2_ASAP7_75t_L g360 ( .A(n_297), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_297), .B(n_354), .Y(n_403) );
OR2x2_ASAP7_75t_L g475 ( .A(n_297), .B(n_362), .Y(n_475) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g395 ( .A(n_301), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx2_ASAP7_75t_L g386 ( .A(n_302), .Y(n_386) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g376 ( .A(n_305), .B(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_305), .Y(n_387) );
OR2x2_ASAP7_75t_L g438 ( .A(n_305), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g493 ( .A(n_305), .Y(n_493) );
AOI211xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B(n_317), .C(n_326), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g382 ( .A(n_310), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_310), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g455 ( .A(n_310), .B(n_332), .Y(n_455) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_313), .B(n_358), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_313), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g465 ( .A(n_313), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g408 ( .A(n_314), .Y(n_408) );
AND2x2_ASAP7_75t_L g436 ( .A(n_315), .B(n_364), .Y(n_436) );
INVx2_ASAP7_75t_L g459 ( .A(n_315), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_315), .B(n_357), .Y(n_491) );
AND2x4_ASAP7_75t_SL g445 ( .A(n_318), .B(n_323), .Y(n_445) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g398 ( .A(n_319), .B(n_324), .Y(n_398) );
OR2x2_ASAP7_75t_L g450 ( .A(n_319), .B(n_343), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_320), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_320), .B(n_332), .Y(n_486) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g434 ( .A(n_321), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g417 ( .A(n_323), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_323), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g467 ( .A(n_324), .Y(n_467) );
BUFx2_ASAP7_75t_L g335 ( .A(n_325), .Y(n_335) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g453 ( .A(n_328), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_332), .Y(n_394) );
NAND3xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_344), .C(n_359), .Y(n_333) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_336), .B1(n_339), .B2(n_341), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_341), .A2(n_367), .B1(n_448), .B2(n_451), .C1(n_453), .C2(n_455), .Y(n_447) );
AND2x2_ASAP7_75t_L g479 ( .A(n_342), .B(n_428), .Y(n_479) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g427 ( .A(n_343), .B(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_350), .B1(n_351), .B2(n_356), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_SL g423 ( .A(n_347), .Y(n_423) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
AND2x2_ASAP7_75t_L g410 ( .A(n_352), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g368 ( .A(n_353), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g362 ( .A(n_354), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g477 ( .A(n_355), .Y(n_477) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_358), .B(n_454), .Y(n_473) );
INVx1_ASAP7_75t_L g490 ( .A(n_358), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B1(n_365), .B2(n_367), .C1(n_370), .C2(n_371), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_366), .Y(n_370) );
AND2x2_ASAP7_75t_L g388 ( .A(n_366), .B(n_389), .Y(n_388) );
INVx3_ASAP7_75t_L g419 ( .A(n_366), .Y(n_419) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g383 ( .A(n_369), .Y(n_383) );
OR2x2_ASAP7_75t_L g452 ( .A(n_369), .B(n_433), .Y(n_452) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_381), .C(n_390), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_388), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_382), .A2(n_420), .B1(n_469), .B2(n_472), .C(n_474), .Y(n_468) );
AND2x4_ASAP7_75t_L g411 ( .A(n_383), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g442 ( .A(n_389), .Y(n_442) );
AOI211x1_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_395), .C(n_399), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_401), .B(n_449), .C(n_450), .Y(n_448) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g484 ( .A(n_402), .Y(n_484) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_456), .Y(n_404) );
NAND4xp25_ASAP7_75t_L g405 ( .A(n_406), .B(n_413), .C(n_435), .D(n_447), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_410), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
AND2x2_ASAP7_75t_L g466 ( .A(n_409), .B(n_467), .Y(n_466) );
AOI221x1_ASAP7_75t_L g435 ( .A1(n_411), .A2(n_436), .B1(n_437), .B2(n_440), .C(n_443), .Y(n_435) );
AND2x2_ASAP7_75t_L g461 ( .A(n_411), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g471 ( .A(n_412), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_420), .B2(n_424), .C(n_426), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_418), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_423), .A2(n_427), .B1(n_430), .B2(n_432), .Y(n_426) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_427), .A2(n_444), .B(n_446), .Y(n_443) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g449 ( .A(n_429), .Y(n_449) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g470 ( .A(n_439), .Y(n_470) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_452), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .C(n_480), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B1(n_464), .B2(n_465), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g476 ( .A(n_463), .B(n_477), .Y(n_476) );
NAND2x1_ASAP7_75t_L g492 ( .A(n_463), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_478), .Y(n_474) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B1(n_485), .B2(n_487), .C(n_489), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g798 ( .A(n_494), .Y(n_798) );
BUFx12f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
XNOR2xp5_ASAP7_75t_L g816 ( .A(n_496), .B(n_817), .Y(n_816) );
NOR2x1p5_ASAP7_75t_L g496 ( .A(n_497), .B(n_708), .Y(n_496) );
NAND4xp75_ASAP7_75t_L g497 ( .A(n_498), .B(n_653), .C(n_673), .D(n_689), .Y(n_497) );
NOR2x1p5_ASAP7_75t_SL g498 ( .A(n_499), .B(n_623), .Y(n_498) );
NAND4xp75_ASAP7_75t_L g499 ( .A(n_500), .B(n_561), .C(n_600), .D(n_609), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_530), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
AND2x4_ASAP7_75t_L g733 ( .A(n_502), .B(n_660), .Y(n_733) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_503), .Y(n_576) );
INVx2_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
AND2x2_ASAP7_75t_L g617 ( .A(n_503), .B(n_579), .Y(n_617) );
OR2x2_ASAP7_75t_L g672 ( .A(n_503), .B(n_511), .Y(n_672) );
AND2x2_ASAP7_75t_L g590 ( .A(n_510), .B(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g740 ( .A(n_510), .B(n_617), .Y(n_740) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
OR2x2_ASAP7_75t_L g577 ( .A(n_511), .B(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g608 ( .A(n_511), .Y(n_608) );
AND2x2_ASAP7_75t_L g614 ( .A(n_511), .B(n_520), .Y(n_614) );
INVx1_ASAP7_75t_L g632 ( .A(n_511), .Y(n_632) );
INVx2_ASAP7_75t_L g661 ( .A(n_511), .Y(n_661) );
INVx3_ASAP7_75t_L g637 ( .A(n_519), .Y(n_637) );
INVx2_ASAP7_75t_L g642 ( .A(n_519), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_519), .B(n_593), .Y(n_647) );
AND2x2_ASAP7_75t_L g670 ( .A(n_519), .B(n_649), .Y(n_670) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_519), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_519), .B(n_725), .Y(n_724) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g659 ( .A(n_520), .Y(n_659) );
AND2x2_ASAP7_75t_L g707 ( .A(n_520), .B(n_661), .Y(n_707) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_543), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_532), .B(n_651), .Y(n_698) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_533), .B(n_651), .Y(n_695) );
INVx1_ASAP7_75t_L g796 ( .A(n_533), .Y(n_796) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g746 ( .A(n_534), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g599 ( .A(n_535), .Y(n_599) );
OR2x2_ASAP7_75t_L g680 ( .A(n_535), .B(n_554), .Y(n_680) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g622 ( .A(n_536), .Y(n_622) );
AND2x4_ASAP7_75t_L g628 ( .A(n_536), .B(n_629), .Y(n_628) );
AOI32xp33_ASAP7_75t_L g766 ( .A1(n_543), .A2(n_669), .A3(n_767), .B1(n_769), .B2(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g715 ( .A(n_544), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_545), .Y(n_563) );
OR2x2_ASAP7_75t_L g597 ( .A(n_545), .B(n_555), .Y(n_597) );
INVx1_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
AND2x2_ASAP7_75t_L g621 ( .A(n_545), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g627 ( .A(n_545), .Y(n_627) );
INVx2_ASAP7_75t_L g652 ( .A(n_545), .Y(n_652) );
AND2x2_ASAP7_75t_L g771 ( .A(n_545), .B(n_565), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_553), .B(n_604), .Y(n_691) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g564 ( .A(n_555), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
INVx2_ASAP7_75t_L g629 ( .A(n_555), .Y(n_629) );
AND2x4_ASAP7_75t_L g651 ( .A(n_555), .B(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_555), .Y(n_743) );
AOI22x1_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_572), .B1(n_590), .B2(n_595), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_564), .B(n_721), .C(n_722), .D(n_723), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_564), .B(n_621), .Y(n_751) );
INVx4_ASAP7_75t_SL g604 ( .A(n_565), .Y(n_604) );
BUFx2_ASAP7_75t_L g667 ( .A(n_565), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_565), .B(n_612), .Y(n_730) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g692 ( .A(n_574), .B(n_641), .Y(n_692) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g615 ( .A(n_578), .B(n_593), .Y(n_615) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_579), .B(n_594), .Y(n_639) );
OAI21x1_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_589), .Y(n_579) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_580), .A2(n_581), .B(n_589), .Y(n_634) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_588), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_591), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g657 ( .A(n_591), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g696 ( .A(n_592), .B(n_614), .Y(n_696) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g739 ( .A(n_594), .B(n_649), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_595), .A2(n_712), .B1(n_714), .B2(n_717), .C(n_719), .Y(n_711) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_L g605 ( .A(n_597), .Y(n_605) );
OR2x2_ASAP7_75t_L g705 ( .A(n_597), .B(n_644), .Y(n_705) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_606), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_601), .A2(n_727), .B1(n_731), .B2(n_734), .Y(n_726) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
AND2x4_ASAP7_75t_L g650 ( .A(n_602), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g762 ( .A(n_602), .B(n_680), .Y(n_762) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g610 ( .A(n_604), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g626 ( .A(n_604), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g685 ( .A(n_604), .B(n_622), .Y(n_685) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_604), .Y(n_702) );
INVx1_ASAP7_75t_L g716 ( .A(n_604), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_604), .B(n_629), .Y(n_759) );
AND2x4_ASAP7_75t_L g666 ( .A(n_605), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g664 ( .A(n_607), .Y(n_664) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_608), .B(n_649), .Y(n_648) );
NAND2x1_ASAP7_75t_L g768 ( .A(n_608), .B(n_670), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_613), .B1(n_616), .B2(n_618), .Y(n_609) );
AND2x2_ASAP7_75t_L g635 ( .A(n_610), .B(n_628), .Y(n_635) );
INVx1_ASAP7_75t_L g676 ( .A(n_610), .Y(n_676) );
AND2x2_ASAP7_75t_L g783 ( .A(n_610), .B(n_644), .Y(n_783) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_SL g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g616 ( .A(n_614), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g756 ( .A(n_614), .Y(n_756) );
AND2x2_ASAP7_75t_L g773 ( .A(n_614), .B(n_633), .Y(n_773) );
AND2x2_ASAP7_75t_L g789 ( .A(n_614), .B(n_739), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_615), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g712 ( .A(n_615), .B(n_713), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_615), .A2(n_705), .B1(n_720), .B2(n_724), .Y(n_719) );
INVx1_ASAP7_75t_L g675 ( .A(n_617), .Y(n_675) );
AND2x2_ASAP7_75t_L g706 ( .A(n_617), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_617), .B(n_713), .Y(n_735) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g741 ( .A(n_621), .B(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_621), .A2(n_645), .B1(n_750), .B2(n_752), .Y(n_749) );
INVx3_ASAP7_75t_L g644 ( .A(n_622), .Y(n_644) );
AND2x2_ASAP7_75t_L g776 ( .A(n_622), .B(n_629), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_640), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_630), .A3(n_633), .B1(n_635), .B2(n_636), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_627), .Y(n_722) );
INVx1_ASAP7_75t_L g747 ( .A(n_627), .Y(n_747) );
INVx3_ASAP7_75t_L g703 ( .A(n_628), .Y(n_703) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_631), .A2(n_779), .B1(n_780), .B2(n_781), .C(n_782), .Y(n_778) );
BUFx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g755 ( .A(n_633), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g791 ( .A(n_633), .B(n_752), .Y(n_791) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g649 ( .A(n_634), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_636), .B(n_664), .Y(n_663) );
AO22x1_ASAP7_75t_L g693 ( .A1(n_636), .A2(n_694), .B1(n_696), .B2(n_697), .Y(n_693) );
NAND2x1p5_ASAP7_75t_L g797 ( .A(n_636), .B(n_664), .Y(n_797) );
AND2x4_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx2_ASAP7_75t_L g713 ( .A(n_637), .Y(n_713) );
INVx1_ASAP7_75t_L g723 ( .A(n_637), .Y(n_723) );
AND2x2_ASAP7_75t_L g643 ( .A(n_638), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_639), .Y(n_725) );
INVx1_ASAP7_75t_L g765 ( .A(n_639), .Y(n_765) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_645), .C(n_650), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR2x1p5_ASAP7_75t_L g752 ( .A(n_642), .B(n_672), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_643), .B(n_702), .Y(n_779) );
AOI31xp33_ASAP7_75t_L g662 ( .A1(n_644), .A2(n_663), .A3(n_665), .B(n_668), .Y(n_662) );
INVx4_ASAP7_75t_L g721 ( .A(n_644), .Y(n_721) );
OR2x2_ASAP7_75t_L g758 ( .A(n_644), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x4_ASAP7_75t_L g660 ( .A(n_649), .B(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_651), .Y(n_656) );
AND2x2_ASAP7_75t_L g687 ( .A(n_651), .B(n_685), .Y(n_687) );
NOR2xp67_ASAP7_75t_L g653 ( .A(n_654), .B(n_662), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g780 ( .A(n_657), .Y(n_780) );
INVx1_ASAP7_75t_L g688 ( .A(n_658), .Y(n_688) );
AND2x4_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g718 ( .A(n_659), .Y(n_718) );
AND2x2_ASAP7_75t_L g717 ( .A(n_660), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .A3(n_677), .B1(n_681), .B2(n_684), .C1(n_686), .C2(n_688), .Y(n_674) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI211x1_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B(n_693), .C(n_699), .Y(n_689) );
INVx1_ASAP7_75t_L g794 ( .A(n_690), .Y(n_794) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g748 ( .A(n_692), .Y(n_748) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OA21x2_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B(n_706), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx2_ASAP7_75t_L g769 ( .A(n_703), .Y(n_769) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp33_ASAP7_75t_L g764 ( .A(n_707), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_777), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_744), .C(n_760), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_726), .C(n_736), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_713), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_717), .A2(n_773), .B(n_774), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_721), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_721), .B(n_771), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_722), .B(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_723), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_733), .A2(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_740), .B(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_749), .C(n_753), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_SL g763 ( .A(n_755), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_759), .Y(n_781) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B(n_766), .C(n_772), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_771), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g792 ( .A(n_771), .Y(n_792) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g788 ( .A(n_776), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_786), .C(n_793), .Y(n_777) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI21xp33_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_790), .B(n_792), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI21xp33_ASAP7_75t_R g793 ( .A1(n_794), .A2(n_795), .B(n_797), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx6_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
BUFx10_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .Y(n_806) );
INVxp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
endmodule