module fake_netlist_5_2125_n_81 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_81);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_81;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

INVx4_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_1),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_20),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AO21x2_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_22),
.B(n_29),
.Y(n_44)
);

OAI21x1_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_24),
.B(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_35),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_41),
.B1(n_21),
.B2(n_31),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_31),
.Y(n_53)
);

OAI221xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_30),
.B1(n_32),
.B2(n_27),
.C(n_25),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

XNOR2x1_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_48),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_49),
.B(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_49),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_32),
.B(n_27),
.Y(n_67)
);

OAI221xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_54),
.B1(n_51),
.B2(n_23),
.C(n_11),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_51),
.B1(n_23),
.B2(n_9),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_65),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_63),
.C(n_8),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_7),
.C(n_13),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_69),
.B1(n_67),
.B2(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_69),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_76),
.B1(n_23),
.B2(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_67),
.B1(n_75),
.B2(n_79),
.Y(n_81)
);


endmodule