module real_jpeg_15221_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_404),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_0),
.B(n_405),
.Y(n_404)
);

NAND2x1p5_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_24),
.Y(n_23)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_1),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AND2x4_ASAP7_75t_SL g123 ( 
.A(n_1),
.B(n_124),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_1),
.B(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_3),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_3),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_4),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_4),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_4),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_4),
.B(n_318),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_5),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_5),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_5),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_6),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_6),
.B(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_7),
.Y(n_170)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_8),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_9),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_9),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_9),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_9),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_9),
.B(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

BUFx4f_ASAP7_75t_L g304 ( 
.A(n_12),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_148),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

CKINVDCx11_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2x1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_19),
.B(n_128),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_95),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_20),
.B(n_70),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_46),
.B1(n_47),
.B2(n_69),
.Y(n_20)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_33),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_35),
.C(n_41),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.C(n_27),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_23),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_122),
.C(n_125),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_23),
.A2(n_72),
.B1(n_73),
.B2(n_120),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_23),
.B(n_52),
.C(n_66),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_23),
.A2(n_120),
.B1(n_125),
.B2(n_144),
.Y(n_357)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_24),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_104),
.C(n_107),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_25),
.A2(n_65),
.B1(n_66),
.B2(n_119),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_25),
.A2(n_66),
.B(n_167),
.C(n_211),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g347 ( 
.A1(n_25),
.A2(n_107),
.B1(n_108),
.B2(n_119),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_26),
.Y(n_163)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_41),
.B2(n_45),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_65),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_41),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_41),
.A2(n_270),
.B(n_276),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_41),
.B(n_270),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_42),
.B(n_106),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_42),
.B(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_60),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_48),
.B(n_60),
.C(n_69),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_49),
.B(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_49),
.A2(n_123),
.B(n_206),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_62),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_51),
.A2(n_52),
.B1(n_179),
.B2(n_183),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_51),
.A2(n_52),
.B1(n_142),
.B2(n_143),
.Y(n_290)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_63),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_65),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_52),
.B(n_56),
.C(n_138),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_52),
.A2(n_179),
.B(n_205),
.C(n_211),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_52),
.B(n_179),
.Y(n_211)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_56),
.B(n_105),
.C(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_56),
.A2(n_57),
.B1(n_104),
.B2(n_105),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_56),
.A2(n_57),
.B1(n_260),
.B2(n_264),
.Y(n_332)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_57),
.B(n_62),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_57),
.B(n_86),
.C(n_260),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_57),
.A2(n_61),
.B(n_68),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B(n_68),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_65),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_65),
.B(n_218),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.C(n_79),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_71),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_74),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_75),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_75),
.A2(n_123),
.B(n_182),
.Y(n_181)
);

NAND2x1p5_ASAP7_75t_L g182 ( 
.A(n_75),
.B(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_75),
.A2(n_102),
.B1(n_194),
.B2(n_195),
.Y(n_247)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_78),
.Y(n_208)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.C(n_89),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_82),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_81),
.A2(n_82),
.B1(n_232),
.B2(n_236),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_81),
.A2(n_82),
.B1(n_181),
.B2(n_184),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_102),
.C(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_82),
.B(n_182),
.C(n_232),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_86),
.A2(n_115),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_86),
.B(n_125),
.C(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_96),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_116),
.C(n_121),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_98),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_112),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_99),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2x1_ASAP7_75t_R g173 ( 
.A(n_102),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_103),
.B(n_112),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_104),
.A2(n_105),
.B1(n_232),
.B2(n_236),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_104),
.B(n_236),
.C(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_105),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_115),
.B(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_116),
.B(n_121),
.Y(n_392)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_122),
.B(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_123),
.A2(n_190),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_123),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_123),
.B(n_206),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_123),
.A2(n_200),
.B1(n_206),
.B2(n_209),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_125),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_125),
.B(n_316),
.C(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_125),
.B(n_296),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_125),
.A2(n_144),
.B1(n_317),
.B2(n_340),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_146),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_145),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_144),
.B(n_296),
.C(n_320),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_396),
.B(n_401),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_384),
.Y(n_149)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_310),
.A3(n_371),
.B1(n_377),
.B2(n_382),
.C(n_383),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_280),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_249),
.B(n_279),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_226),
.B(n_248),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_202),
.B(n_225),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_185),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_156),
.B(n_185),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_171),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_165),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_165),
.C(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_162),
.A2(n_245),
.B1(n_259),
.B2(n_265),
.Y(n_258)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_167),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_166),
.A2(n_167),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_217),
.B(n_219),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_173),
.A2(n_179),
.B(n_184),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_198),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_198),
.B1(n_199),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_190),
.B(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_194),
.A2(n_195),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_195),
.B(n_297),
.C(n_301),
.Y(n_316)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_215),
.B(n_224),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_206),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_206),
.A2(n_209),
.B1(n_260),
.B2(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_206),
.B(n_245),
.C(n_260),
.Y(n_307)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_220),
.B(n_223),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

XOR2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_238),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_237),
.C(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_243),
.C(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_278),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_278),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_266),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_253),
.C(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_258),
.C(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_257),
.B(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_277),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_269),
.C(n_277),
.Y(n_309)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_276),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_281),
.B(n_282),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_293),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_283),
.B(n_294),
.C(n_309),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_289),
.B2(n_290),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_367)
);

XNOR2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_309),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_305),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_307),
.C(n_308),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_359),
.Y(n_310)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_348),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_312),
.B(n_348),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_333),
.C(n_341),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_313),
.B(n_341),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_319),
.B1(n_324),
.B2(n_325),
.Y(n_314)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_325),
.C(n_326),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_327),
.A2(n_328),
.B1(n_330),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.C(n_337),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_344),
.C(n_346),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_353),
.C(n_387),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_356),
.C(n_358),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

AOI31xp67_ASAP7_75t_SL g377 ( 
.A1(n_359),
.A2(n_372),
.A3(n_378),
.B(n_381),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_362),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.C(n_368),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_363),
.A2(n_364),
.B1(n_368),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_376),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_388),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_391),
.C(n_393),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_400),
.Y(n_403)
);


endmodule