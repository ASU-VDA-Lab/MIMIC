module fake_ariane_186_n_57 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_57);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_57;

wire n_56;
wire n_24;
wire n_22;
wire n_43;
wire n_49;
wire n_27;
wire n_20;
wire n_48;
wire n_29;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_47;
wire n_32;
wire n_18;
wire n_28;
wire n_37;
wire n_51;
wire n_45;
wire n_34;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_33;
wire n_44;
wire n_19;
wire n_30;
wire n_39;
wire n_40;
wire n_31;
wire n_42;
wire n_53;
wire n_21;
wire n_23;
wire n_35;
wire n_54;
wire n_25;

AND2x6_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_14),
.Y(n_18)
);

AND2x6_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_6),
.B1(n_11),
.B2(n_7),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_13),
.B1(n_3),
.B2(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

OAI22x1_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_4),
.B1(n_15),
.B2(n_3),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_21),
.Y(n_32)
);

NOR2x1p5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_28),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_18),
.B(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_35),
.B1(n_30),
.B2(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_40),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_50),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_29),
.C(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_18),
.B1(n_29),
.B2(n_19),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_48),
.Y(n_57)
);


endmodule