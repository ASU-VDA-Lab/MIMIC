module fake_jpeg_22261_n_241 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_48),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_29),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_35),
.Y(n_74)
);

NAND2x1_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_28),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_56),
.A2(n_75),
.B1(n_81),
.B2(n_42),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_23),
.B1(n_17),
.B2(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_31),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_63),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_25),
.B1(n_19),
.B2(n_27),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_58),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_19),
.B1(n_38),
.B2(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_36),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_74),
.B(n_1),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_35),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_34),
.C(n_33),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_5),
.B(n_6),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_32),
.B1(n_26),
.B2(n_18),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_32),
.B1(n_26),
.B2(n_18),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_89),
.B1(n_93),
.B2(n_105),
.Y(n_116)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_96),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_44),
.B1(n_23),
.B2(n_17),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_46),
.B1(n_42),
.B2(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_23),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_46),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_55),
.Y(n_127)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_78),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_46),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_105),
.B1(n_102),
.B2(n_86),
.Y(n_122)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_115),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_121),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_74),
.B(n_70),
.C(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_131),
.B1(n_109),
.B2(n_73),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_67),
.B(n_65),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_129),
.B(n_130),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_68),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_67),
.B(n_70),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_70),
.B(n_55),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_73),
.B1(n_82),
.B2(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_68),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_138),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_54),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_151),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_107),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_126),
.B(n_114),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_159),
.C(n_119),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_154),
.B1(n_158),
.B2(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_120),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_114),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_157),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_54),
.B1(n_100),
.B2(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_108),
.B1(n_96),
.B2(n_84),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_76),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_76),
.B1(n_97),
.B2(n_95),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_84),
.B1(n_97),
.B2(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_142),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_171),
.C(n_180),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_124),
.C(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_172),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_132),
.B(n_115),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_174),
.B1(n_175),
.B2(n_147),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_117),
.C(n_113),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_162),
.B1(n_147),
.B2(n_140),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_126),
.B(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_131),
.C(n_123),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_123),
.C(n_92),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_145),
.C(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_190),
.C(n_193),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_189),
.B1(n_195),
.B2(n_165),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_175),
.C(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_197),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_149),
.C(n_158),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_153),
.B1(n_150),
.B2(n_163),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_154),
.C(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_198),
.C(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_152),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_180),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_205),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_176),
.A3(n_168),
.B1(n_179),
.B2(n_181),
.C1(n_172),
.C2(n_177),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_210),
.B(n_202),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_176),
.B(n_165),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_206),
.B(n_207),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_194),
.B(n_184),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_205),
.B(n_203),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_188),
.C(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_7),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_207),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_202),
.C(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_7),
.C(n_8),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_218),
.B(n_216),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_12),
.B1(n_219),
.B2(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_219),
.C(n_11),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_224),
.Y(n_227)
);

BUFx12f_ASAP7_75t_SL g223 ( 
.A(n_211),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_10),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_221),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_230),
.C(n_227),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.C(n_233),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_234),
.C(n_12),
.Y(n_240)
);


endmodule