module fake_jpeg_31825_n_542 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_56),
.B(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g158 ( 
.A(n_70),
.Y(n_158)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_28),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_71),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_22),
.A2(n_16),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_72),
.B(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_22),
.B(n_0),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_28),
.Y(n_84)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_23),
.B(n_3),
.Y(n_100)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_29),
.B(n_4),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_30),
.B1(n_34),
.B2(n_44),
.Y(n_124)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_37),
.B1(n_21),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_111),
.A2(n_118),
.B1(n_130),
.B2(n_143),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_37),
.B1(n_21),
.B2(n_32),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_49),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_57),
.A2(n_32),
.B1(n_40),
.B2(n_50),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_159),
.B1(n_53),
.B2(n_41),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_34),
.B1(n_30),
.B2(n_40),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_58),
.A2(n_34),
.B1(n_30),
.B2(n_45),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_27),
.B1(n_46),
.B2(n_45),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_144),
.A2(n_148),
.B1(n_151),
.B2(n_59),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_24),
.B1(n_46),
.B2(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_48),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_87),
.A2(n_24),
.B1(n_36),
.B2(n_33),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_62),
.A2(n_53),
.B1(n_33),
.B2(n_27),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_60),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_159)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_173),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_109),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_178),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_125),
.B1(n_139),
.B2(n_137),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_106),
.B1(n_105),
.B2(n_64),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_179),
.B1(n_183),
.B2(n_209),
.Y(n_225)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_110),
.B(n_29),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_108),
.A2(n_86),
.B1(n_98),
.B2(n_65),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_182),
.A2(n_215),
.B1(n_220),
.B2(n_221),
.Y(n_236)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_188),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_43),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_191),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_107),
.B(n_90),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_48),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_101),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_195),
.B(n_200),
.Y(n_257)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_199),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_95),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_97),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_201),
.Y(n_248)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_162),
.B(n_59),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_203),
.B(n_213),
.Y(n_235)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_134),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_66),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_208),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_164),
.B1(n_156),
.B2(n_163),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_96),
.C(n_63),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_212),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_74),
.Y(n_214)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx3_ASAP7_75t_SL g218 ( 
.A(n_119),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_151),
.A2(n_70),
.A3(n_89),
.B1(n_80),
.B2(n_78),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_219),
.A2(n_130),
.B(n_112),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_224),
.A2(n_218),
.B(n_222),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_161),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_216),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_161),
.B1(n_149),
.B2(n_142),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_239),
.A2(n_241),
.B1(n_253),
.B2(n_208),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_176),
.A2(n_149),
.B1(n_129),
.B2(n_142),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_265),
.B1(n_243),
.B2(n_249),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_179),
.B1(n_136),
.B2(n_117),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_143),
.B(n_5),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_256),
.A2(n_5),
.B(n_6),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_209),
.A2(n_118),
.B1(n_111),
.B2(n_92),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_260),
.A2(n_264),
.B1(n_61),
.B2(n_194),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_207),
.A2(n_67),
.B1(n_125),
.B2(n_129),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_221),
.A2(n_139),
.B1(n_137),
.B2(n_136),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_292),
.B(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_270),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_171),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_196),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_274),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_192),
.C(n_181),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_273),
.B(n_275),
.C(n_255),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_229),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_233),
.B(n_169),
.C(n_205),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_231),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_278),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_227),
.B(n_204),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_281),
.Y(n_318)
);

AO22x1_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_197),
.B1(n_187),
.B2(n_173),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_293),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_206),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_224),
.A2(n_210),
.B(n_177),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_282),
.A2(n_295),
.B(n_296),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_206),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_286),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_285),
.B1(n_294),
.B2(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_231),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_297),
.Y(n_333)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_246),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_291),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_172),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_236),
.A2(n_224),
.B(n_231),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_172),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_51),
.B1(n_6),
.B2(n_7),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_238),
.A2(n_51),
.B(n_6),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_264),
.B1(n_262),
.B2(n_249),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_245),
.A2(n_51),
.B(n_8),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_248),
.B(n_243),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_230),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_225),
.A2(n_51),
.B1(n_8),
.B2(n_10),
.Y(n_301)
);

OA22x2_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_51),
.B1(n_8),
.B2(n_10),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_226),
.Y(n_326)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_303),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_234),
.A2(n_7),
.B(n_8),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_252),
.B(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_274),
.B(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_309),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_307),
.A2(n_316),
.B(n_282),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_271),
.B(n_251),
.Y(n_309)
);

NAND2x1_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_265),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_310),
.A2(n_313),
.B(n_304),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_315),
.B1(n_339),
.B2(n_285),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_280),
.A2(n_267),
.B1(n_248),
.B2(n_226),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_251),
.B1(n_249),
.B2(n_259),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_234),
.B(n_255),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_279),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_319),
.B(n_281),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_326),
.A2(n_298),
.B1(n_269),
.B2(n_302),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_327),
.B(n_283),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_240),
.C(n_252),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_334),
.C(n_327),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_286),
.B(n_240),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_331),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_226),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_261),
.C(n_254),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_261),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_302),
.Y(n_362)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_338),
.B(n_291),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_259),
.B1(n_232),
.B2(n_250),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_268),
.B(n_293),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_340),
.A2(n_369),
.B(n_333),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_321),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_341),
.B(n_346),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_293),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_342),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_326),
.A2(n_296),
.B1(n_298),
.B2(n_282),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_365),
.B1(n_367),
.B2(n_322),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_321),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_361),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_349),
.A2(n_354),
.B1(n_356),
.B2(n_317),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_272),
.Y(n_350)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_351),
.A2(n_360),
.B(n_340),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_352),
.B(n_358),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_311),
.A2(n_339),
.B1(n_308),
.B2(n_323),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_275),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_371),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_315),
.B1(n_296),
.B2(n_294),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_357),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_337),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_359),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_323),
.A2(n_293),
.B(n_288),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_362),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_366),
.C(n_328),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_275),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_364),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_317),
.A2(n_284),
.B1(n_301),
.B2(n_302),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_370),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_300),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_303),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_320),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_325),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_376),
.C(n_379),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_374),
.A2(n_349),
.B1(n_365),
.B2(n_367),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_351),
.A2(n_316),
.B(n_314),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_375),
.A2(n_389),
.B(n_393),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_334),
.C(n_306),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_399),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_334),
.C(n_312),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_356),
.A2(n_322),
.B1(n_305),
.B2(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_335),
.C(n_314),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_391),
.C(n_394),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_318),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_387),
.B(n_404),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_333),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_348),
.A2(n_324),
.B(n_338),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_392),
.B(n_369),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_320),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_345),
.B(n_324),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_398),
.C(n_341),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_330),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_352),
.Y(n_407)
);

AO22x1_ASAP7_75t_L g402 ( 
.A1(n_343),
.A2(n_310),
.B1(n_307),
.B2(n_302),
.Y(n_402)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_402),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_332),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_420),
.Y(n_435)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_396),
.Y(n_408)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_390),
.Y(n_410)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_402),
.Y(n_413)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_406),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_346),
.Y(n_417)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_417),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_418),
.B(n_431),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_347),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_383),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_381),
.B(n_347),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_426),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_388),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_354),
.C(n_342),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_382),
.C(n_376),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_428),
.A2(n_429),
.B1(n_377),
.B2(n_402),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_374),
.A2(n_342),
.B1(n_310),
.B2(n_368),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_430),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_295),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_397),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_237),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_433),
.B(n_400),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_382),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_437),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_439),
.B(n_452),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_441),
.A2(n_443),
.B1(n_419),
.B2(n_423),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_403),
.B1(n_404),
.B2(n_391),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_420),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_451),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_SL g450 ( 
.A(n_411),
.B(n_392),
.Y(n_450)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_411),
.B(n_389),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_379),
.C(n_387),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_456),
.C(n_457),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_412),
.B(n_416),
.C(n_418),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_393),
.C(n_378),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_430),
.C(n_432),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_468),
.C(n_469),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_457),
.A2(n_438),
.B(n_456),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_463),
.A2(n_424),
.B(n_421),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_415),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_474),
.Y(n_493)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_435),
.Y(n_466)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_449),
.A2(n_405),
.B1(n_425),
.B2(n_413),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_467),
.A2(n_449),
.B1(n_469),
.B2(n_447),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_406),
.C(n_415),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_405),
.C(n_429),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_470),
.B(n_299),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_442),
.B(n_408),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_473),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_417),
.C(n_409),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_474),
.C(n_440),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_441),
.A2(n_410),
.B1(n_426),
.B2(n_422),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_436),
.C(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_476),
.B(n_447),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_479),
.B(n_480),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_461),
.A2(n_446),
.B1(n_452),
.B2(n_419),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_486),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_448),
.C(n_453),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_494),
.C(n_465),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_459),
.B(n_453),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_483),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_487),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_485),
.A2(n_492),
.B(n_287),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_419),
.B(n_431),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_468),
.A2(n_310),
.B1(n_344),
.B2(n_361),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_490),
.A2(n_237),
.B1(n_250),
.B2(n_254),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_458),
.B(n_460),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_493),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_462),
.A2(n_344),
.B1(n_325),
.B2(n_329),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_325),
.C(n_332),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_493),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_497),
.B(n_509),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_488),
.A2(n_464),
.B1(n_472),
.B2(n_284),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_503),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_465),
.C(n_289),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_501),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_228),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_301),
.B1(n_259),
.B2(n_302),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_479),
.C(n_482),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_242),
.C(n_12),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_266),
.C(n_232),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_506),
.Y(n_519)
);

INVx11_ASAP7_75t_L g509 ( 
.A(n_490),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_496),
.A2(n_481),
.B(n_477),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_510),
.A2(n_511),
.B(n_501),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_486),
.B(n_489),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_508),
.A2(n_487),
.B1(n_242),
.B2(n_228),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_520),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_495),
.A2(n_228),
.B(n_242),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_514),
.B(n_520),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_242),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_521),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_11),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_507),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_508),
.B1(n_500),
.B2(n_509),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_523),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_515),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_527),
.C(n_528),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_525),
.A2(n_516),
.B(n_517),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_526),
.C(n_518),
.Y(n_533)
);

OAI21x1_ASAP7_75t_SL g531 ( 
.A1(n_525),
.A2(n_513),
.B(n_519),
.Y(n_531)
);

O2A1O1Ixp33_ASAP7_75t_SL g535 ( 
.A1(n_531),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_533),
.A2(n_534),
.B(n_16),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_532),
.C(n_13),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_11),
.B(n_14),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_536),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_537),
.B(n_14),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_15),
.C(n_537),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_15),
.Y(n_542)
);


endmodule