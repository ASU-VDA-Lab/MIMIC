module fake_jpeg_23405_n_322 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_26),
.B(n_37),
.C(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_33),
.B1(n_28),
.B2(n_18),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_52),
.B1(n_55),
.B2(n_68),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_28),
.B1(n_29),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_33),
.B1(n_25),
.B2(n_30),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_56),
.A2(n_17),
.B(n_16),
.Y(n_114)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_33),
.B1(n_20),
.B2(n_27),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_59),
.B1(n_72),
.B2(n_81),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_38),
.B1(n_37),
.B2(n_24),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_83),
.B1(n_68),
.B2(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_82),
.B1(n_87),
.B2(n_0),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_85),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_26),
.B1(n_35),
.B2(n_34),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_35),
.B1(n_34),
.B2(n_22),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_86),
.B1(n_0),
.B2(n_1),
.Y(n_98)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_41),
.A2(n_19),
.B1(n_36),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_39),
.A2(n_36),
.B1(n_23),
.B2(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_10),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_39),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_104),
.Y(n_137)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_97),
.B(n_100),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_153)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_99),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_102),
.B(n_103),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_112),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_50),
.B1(n_69),
.B2(n_54),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_109),
.B(n_120),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_52),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_121),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_15),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_52),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_65),
.B(n_13),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_124),
.B(n_130),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_52),
.B1(n_87),
.B2(n_51),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_142),
.B1(n_151),
.B2(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_127),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_191)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_138),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_12),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_143),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_50),
.B1(n_69),
.B2(n_75),
.Y(n_136)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_107),
.B1(n_113),
.B2(n_93),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_105),
.B1(n_112),
.B2(n_91),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_77),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_76),
.B(n_119),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_57),
.B1(n_75),
.B2(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_63),
.C(n_64),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_78),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_1),
.Y(n_146)
);

XOR2x2_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_2),
.Y(n_187)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_78),
.B1(n_76),
.B2(n_79),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_158),
.B(n_159),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx24_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_164),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_108),
.B(n_117),
.C(n_114),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_163),
.A2(n_177),
.B(n_181),
.Y(n_219)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_111),
.B1(n_122),
.B2(n_118),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_137),
.B1(n_125),
.B2(n_151),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_89),
.B(n_104),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_184),
.B(n_187),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_157),
.C(n_143),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_126),
.B1(n_150),
.B2(n_125),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_130),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_200),
.C(n_201),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_126),
.B1(n_125),
.B2(n_150),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_199),
.B1(n_187),
.B2(n_182),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_134),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_151),
.B(n_124),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_158),
.B(n_189),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_151),
.B1(n_147),
.B2(n_106),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_215),
.B1(n_220),
.B2(n_164),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_129),
.C(n_89),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_217),
.C(n_146),
.Y(n_242)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_162),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_106),
.B1(n_96),
.B2(n_133),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_146),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_106),
.B1(n_96),
.B2(n_133),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_236),
.C(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_171),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_230),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_241),
.B1(n_195),
.B2(n_198),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_167),
.C(n_212),
.Y(n_229)
);

OAI322xp33_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_239),
.A3(n_209),
.B1(n_193),
.B2(n_202),
.C1(n_206),
.C2(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_169),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_192),
.CI(n_219),
.CON(n_247),
.SN(n_247)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_233),
.B(n_234),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_215),
.B1(n_213),
.B2(n_206),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_179),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_204),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_238),
.B(n_240),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_192),
.B(n_123),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_165),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_244),
.B(n_216),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_186),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_258),
.B1(n_222),
.B2(n_227),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_262),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_200),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_254),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_239),
.B(n_234),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_199),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_256),
.C(n_225),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_211),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_195),
.B1(n_213),
.B2(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_210),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_230),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_231),
.A2(n_220),
.B1(n_214),
.B2(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_238),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_264),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_242),
.A3(n_237),
.B1(n_232),
.B2(n_240),
.C1(n_228),
.C2(n_223),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_279),
.B(n_257),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_274),
.C(n_277),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_226),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_258),
.B1(n_252),
.B2(n_246),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_243),
.C(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_160),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_160),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_129),
.C(n_123),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_138),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_180),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_276),
.B(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_247),
.B1(n_277),
.B2(n_178),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_245),
.C(n_252),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_293),
.B(n_274),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_245),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_278),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_262),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_280),
.B1(n_264),
.B2(n_247),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_254),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_297),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_299),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_271),
.B1(n_259),
.B2(n_263),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_298),
.B(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_281),
.B(n_3),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_178),
.B(n_116),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_284),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_295),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_308),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_291),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_283),
.B(n_284),
.Y(n_314)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_288),
.B(n_293),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_289),
.A3(n_116),
.B1(n_95),
.B2(n_8),
.C1(n_7),
.C2(n_6),
.Y(n_317)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_290),
.B(n_283),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

OAI31xp33_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_304),
.A3(n_306),
.B(n_308),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_317),
.A3(n_312),
.B1(n_95),
.B2(n_7),
.C1(n_8),
.C2(n_6),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_319),
.C(n_95),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_5),
.B1(n_8),
.B2(n_304),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_5),
.Y(n_322)
);


endmodule