module real_jpeg_32921_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_653;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_531;
wire n_172;
wire n_285;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_686;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g192 ( 
.A(n_0),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_0),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_0),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_1),
.A2(n_54),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_1),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_1),
.A2(n_238),
.B1(n_358),
.B2(n_363),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g530 ( 
.A1(n_1),
.A2(n_238),
.B1(n_531),
.B2(n_534),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_1),
.A2(n_238),
.B1(n_571),
.B2(n_577),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_2),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_4),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_4),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_4),
.A2(n_117),
.B1(n_256),
.B2(n_312),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_4),
.A2(n_256),
.B1(n_404),
.B2(n_510),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_4),
.A2(n_256),
.B1(n_552),
.B2(n_557),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_R g25 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_5),
.A2(n_34),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_34),
.B1(n_148),
.B2(n_153),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_5),
.A2(n_34),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_6),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_6),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_6),
.A2(n_248),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_6),
.A2(n_248),
.B1(n_342),
.B2(n_344),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_6),
.A2(n_248),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_7),
.B(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_7),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_7),
.B(n_36),
.Y(n_388)
);

OAI32xp33_ASAP7_75t_L g483 ( 
.A1(n_7),
.A2(n_484),
.A3(n_486),
.B1(n_490),
.B2(n_496),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g528 ( 
.A1(n_7),
.A2(n_484),
.A3(n_486),
.B1(n_490),
.B2(n_496),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_7),
.A2(n_354),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

OAI21xp33_ASAP7_75t_L g616 ( 
.A1(n_7),
.A2(n_280),
.B(n_562),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_8),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_8),
.A2(n_286),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_8),
.A2(n_286),
.B1(n_379),
.B2(n_383),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_8),
.A2(n_286),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_9),
.A2(n_27),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_9),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_115),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_9),
.A2(n_115),
.B1(n_293),
.B2(n_298),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_9),
.A2(n_115),
.B1(n_262),
.B2(n_433),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_12),
.Y(n_576)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_20),
.B(n_685),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_14),
.B(n_686),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_15),
.A2(n_52),
.B1(n_153),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_15),
.A2(n_52),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_15),
.A2(n_52),
.B1(n_404),
.B2(n_408),
.Y(n_403)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_16),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_16),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_16),
.Y(n_407)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_17),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_17),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_18),
.A2(n_55),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_18),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_18),
.A2(n_124),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_18),
.A2(n_124),
.B1(n_326),
.B2(n_329),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_18),
.A2(n_124),
.B1(n_426),
.B2(n_429),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_177),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_176),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_70),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_24),
.B(n_70),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_35),
.B1(n_51),
.B2(n_59),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_29),
.Y(n_225)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_33),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_33),
.Y(n_418)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_35),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_35),
.A2(n_51),
.B1(n_59),
.B2(n_170),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g648 ( 
.A1(n_35),
.A2(n_59),
.B1(n_114),
.B2(n_414),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_36),
.B(n_237),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g310 ( 
.A1(n_36),
.A2(n_60),
.B1(n_237),
.B2(n_311),
.Y(n_310)
);

NAND2x1_ASAP7_75t_SL g348 ( 
.A(n_36),
.B(n_243),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_36),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_41),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_41),
.Y(n_431)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_42),
.Y(n_221)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_44),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_45),
.A2(n_157),
.B1(n_160),
.B2(n_163),
.Y(n_156)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_45),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_46),
.Y(n_259)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_58),
.Y(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_58),
.Y(n_250)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_60),
.B(n_243),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_60),
.A2(n_226),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_60),
.B(n_311),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_63),
.Y(n_313)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_169),
.C(n_171),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_71),
.B(n_642),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_110),
.C(n_130),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_72),
.A2(n_73),
.B1(n_652),
.B2(n_653),
.Y(n_663)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_73),
.B(n_131),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_73),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_90),
.B(n_105),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_74),
.A2(n_90),
.B1(n_341),
.B2(n_346),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_74),
.A2(n_90),
.B1(n_105),
.B2(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_74),
.B(n_341),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_74),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_75),
.Y(n_301)
);

OAI22x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_83),
.B2(n_87),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_82),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_82),
.Y(n_279)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_82),
.Y(n_382)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_83),
.Y(n_595)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_86),
.Y(n_321)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_86),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_88),
.Y(n_587)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_89),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_90),
.B(n_606),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_91),
.A2(n_283),
.B1(n_292),
.B2(n_301),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_91),
.A2(n_292),
.B1(n_301),
.B2(n_325),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_91),
.A2(n_301),
.B1(n_325),
.B2(n_403),
.Y(n_402)
);

OAI21xp33_ASAP7_75t_SL g508 ( 
.A1(n_91),
.A2(n_509),
.B(n_513),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_91),
.A2(n_301),
.B1(n_509),
.B2(n_530),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_91),
.A2(n_530),
.B1(n_546),
.B2(n_547),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_100),
.B2(n_102),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_95),
.Y(n_501)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_102),
.Y(n_343)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_104),
.Y(n_285)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_104),
.Y(n_297)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_109),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_111),
.B(n_647),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_123),
.B2(n_129),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_122),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g415 ( 
.A(n_128),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_147),
.B1(n_155),
.B2(n_166),
.Y(n_131)
);

AOI22x1_ASAP7_75t_L g355 ( 
.A1(n_132),
.A2(n_356),
.B1(n_357),
.B2(n_366),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_132),
.A2(n_155),
.B1(n_425),
.B2(n_432),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_132),
.A2(n_166),
.B1(n_356),
.B2(n_425),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_133),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_133),
.A2(n_155),
.B1(n_306),
.B2(n_432),
.Y(n_445)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_141),
.B2(n_145),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_139),
.Y(n_300)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_140),
.Y(n_489)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_144),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_155),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_151),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_152),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_152),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_155),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_155),
.B(n_261),
.Y(n_376)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_159),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_168),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_643),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_169),
.Y(n_643)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g374 ( 
.A1(n_174),
.A2(n_375),
.B(n_376),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g303 ( 
.A1(n_175),
.A2(n_252),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_175),
.B(n_354),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_637),
.B(n_674),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_473),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_393),
.B(n_467),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_332),
.C(n_367),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_182),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_266),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_183),
.B(n_267),
.C(n_314),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_235),
.C(n_251),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_185),
.B(n_335),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_216),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_186),
.B(n_216),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_193),
.B1(n_203),
.B2(n_209),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_187),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_187),
.B(n_504),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_187),
.A2(n_569),
.B1(n_580),
.B2(n_582),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_190),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_192),
.Y(n_318)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_194),
.A2(n_280),
.B1(n_378),
.B2(n_384),
.Y(n_377)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_198),
.Y(n_275)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_198),
.Y(n_556)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_201),
.Y(n_383)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_203),
.B(n_504),
.Y(n_562)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_208),
.Y(n_386)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_211),
.Y(n_506)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_214),
.Y(n_505)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_221),
.A3(n_222),
.B1(n_226),
.B2(n_228),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_219),
.Y(n_231)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_220),
.Y(n_436)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_231),
.Y(n_491)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_235),
.B(n_251),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_242),
.B(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B(n_260),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_252),
.A2(n_260),
.B(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_253),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_314),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_302),
.Y(n_267)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_268),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_282),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_282),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_273),
.B1(n_280),
.B2(n_281),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_273),
.A2(n_280),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_279),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_280),
.A2(n_319),
.B(n_400),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_280),
.A2(n_551),
.B(n_562),
.Y(n_550)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_285),
.Y(n_409)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_291),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_291),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_291),
.Y(n_600)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_297),
.Y(n_593)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_303),
.Y(n_459)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_310),
.Y(n_458)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_316),
.B(n_324),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_332),
.Y(n_476)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.C(n_338),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_333),
.A2(n_334),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_339),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_347),
.C(n_355),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_341),
.Y(n_547)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NAND2x1_ASAP7_75t_SL g440 ( 
.A(n_348),
.B(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_354),
.B(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_354),
.B(n_590),
.Y(n_589)
);

OAI21xp33_ASAP7_75t_SL g606 ( 
.A1(n_354),
.A2(n_589),
.B(n_607),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_354),
.B(n_546),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_354),
.B(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_389),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_368),
.B(n_389),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.C(n_372),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_369),
.B(n_519),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_371),
.B(n_373),
.Y(n_519)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.C(n_387),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_374),
.B(n_516),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_377),
.A2(n_387),
.B1(n_388),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_377),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_378),
.A2(n_400),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx12f_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_394),
.B(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_395),
.A2(n_447),
.B(n_462),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_395),
.B(n_447),
.Y(n_472)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_396),
.B(n_448),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_420),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_397),
.B(n_669),
.C(n_670),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_410),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_398),
.A2(n_412),
.B(n_419),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_399),
.A2(n_411),
.B1(n_412),
.B2(n_419),
.Y(n_410)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_399),
.A2(n_402),
.B1(n_419),
.B2(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_400),
.A2(n_503),
.B(n_570),
.Y(n_614)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_403),
.Y(n_423)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_406),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_438),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_421),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_424),
.B(n_437),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_424),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_437),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_437),
.Y(n_673)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_438),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.C(n_446),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_440),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_445),
.Y(n_454)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_443),
.A2(n_452),
.B(n_454),
.Y(n_451)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_446),
.Y(n_455)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_456),
.C(n_460),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_465),
.Y(n_464)
);

XNOR2x1_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_455),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.C(n_459),
.Y(n_456)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_460),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_463),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_466),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_471),
.B(n_472),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_478),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_520),
.B(n_635),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_518),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_481),
.B(n_636),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_507),
.C(n_514),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_482),
.A2(n_507),
.B1(n_508),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_502),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_500),
.Y(n_609)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_502),
.B(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_511),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_513),
.B(n_605),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_518),
.Y(n_636)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_563),
.B(n_634),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_541),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_523),
.B(n_526),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_529),
.C(n_535),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_527),
.B(n_543),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_535),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_532),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_542),
.B(n_544),
.Y(n_541)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_542),
.Y(n_632)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_548),
.C(n_550),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_545),
.B(n_549),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_550),
.B(n_627),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_551),
.Y(n_582)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_556),
.Y(n_561)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_630),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_625),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_566),
.A2(n_610),
.B(n_624),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_583),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_568),
.B(n_583),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_581),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_604),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_584),
.B(n_604),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_585),
.A2(n_588),
.B1(n_594),
.B2(n_596),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_587),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_601),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_612),
.A2(n_615),
.B(n_623),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_614),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_613),
.B(n_614),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_616),
.B(n_617),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_618),
.B(n_620),
.Y(n_617)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_626),
.B(n_628),
.Y(n_625)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_626),
.Y(n_633)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_629),
.A2(n_631),
.B1(n_632),
.B2(n_633),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_638),
.B(n_655),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_638),
.A2(n_675),
.B(n_683),
.Y(n_674)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_640),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_644),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_641),
.B(n_644),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_645),
.B(n_648),
.C(n_649),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_646),
.B(n_654),
.Y(n_659)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_648),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_663),
.Y(n_662)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g658 ( 
.A(n_650),
.B(n_659),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_652),
.C(n_654),
.Y(n_650)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_657),
.B(n_667),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_657),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_658),
.B(n_660),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_658),
.B(n_681),
.C(n_682),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_661),
.B(n_665),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_661),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_664),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_662),
.A2(n_664),
.B(n_666),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_SL g671 ( 
.A(n_662),
.B(n_672),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_665),
.Y(n_681)
);

XOR2xp5_ASAP7_75t_L g672 ( 
.A(n_666),
.B(n_673),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_668),
.B(n_671),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_668),
.B(n_671),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_676),
.A2(n_677),
.B(n_679),
.Y(n_675)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_678),
.Y(n_677)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_680),
.Y(n_679)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_684),
.Y(n_683)
);


endmodule