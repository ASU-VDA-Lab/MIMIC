module real_aes_8809_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_148;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g163 ( .A1(n_0), .A2(n_164), .B(n_167), .C(n_171), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_1), .B(n_155), .Y(n_174) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_3), .B(n_165), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_4), .A2(n_124), .B(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_129), .B(n_132), .C(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_6), .A2(n_124), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_7), .B(n_155), .Y(n_473) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_8), .A2(n_157), .B(n_232), .Y(n_231) );
AND2x6_ASAP7_75t_L g129 ( .A(n_9), .B(n_130), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_10), .A2(n_129), .B(n_132), .C(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g507 ( .A(n_11), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_12), .B(n_42), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_13), .B(n_170), .Y(n_496) );
INVx1_ASAP7_75t_L g150 ( .A(n_14), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_15), .B(n_165), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_16), .A2(n_166), .B(n_527), .C(n_529), .Y(n_526) );
AOI222xp33_ASAP7_75t_SL g102 ( .A1(n_17), .A2(n_103), .B1(n_104), .B2(n_107), .C1(n_691), .C2(n_695), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_18), .B(n_155), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_19), .B(n_144), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_20), .A2(n_132), .B(n_135), .C(n_143), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_21), .A2(n_169), .B(n_225), .C(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_22), .B(n_170), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_23), .A2(n_41), .B1(n_105), .B2(n_106), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_23), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_24), .B(n_170), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_25), .Y(n_441) );
INVx1_ASAP7_75t_L g480 ( .A(n_26), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_27), .A2(n_132), .B(n_143), .C(n_235), .Y(n_234) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_28), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_29), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_30), .A2(n_101), .B1(n_700), .B2(n_709), .C1(n_721), .C2(n_727), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_30), .A2(n_77), .B1(n_713), .B2(n_714), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_30), .Y(n_714) );
INVx1_ASAP7_75t_L g458 ( .A(n_31), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_32), .A2(n_124), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g127 ( .A(n_33), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_34), .A2(n_183), .B(n_184), .C(n_188), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_35), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_36), .A2(n_169), .B(n_470), .C(n_472), .Y(n_469) );
INVxp67_ASAP7_75t_L g459 ( .A(n_37), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_38), .B(n_237), .Y(n_236) );
CKINVDCx14_ASAP7_75t_R g468 ( .A(n_39), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_40), .A2(n_132), .B(n_143), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_41), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_43), .A2(n_171), .B(n_505), .C(n_506), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_44), .B(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_45), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_46), .B(n_165), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_47), .B(n_124), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_48), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_49), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_50), .A2(n_183), .B(n_188), .C(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g168 ( .A(n_51), .Y(n_168) );
INVx1_ASAP7_75t_L g211 ( .A(n_52), .Y(n_211) );
INVx1_ASAP7_75t_L g513 ( .A(n_53), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_54), .B(n_124), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_55), .Y(n_152) );
CKINVDCx14_ASAP7_75t_R g503 ( .A(n_56), .Y(n_503) );
INVx1_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_58), .B(n_124), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_59), .B(n_155), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_60), .A2(n_142), .B(n_198), .C(n_200), .Y(n_197) );
INVx1_ASAP7_75t_L g149 ( .A(n_61), .Y(n_149) );
INVx1_ASAP7_75t_SL g471 ( .A(n_62), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_63), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_64), .B(n_165), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_65), .B(n_155), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_66), .B(n_166), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_67), .Y(n_719) );
INVx1_ASAP7_75t_L g444 ( .A(n_68), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_69), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_70), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_71), .A2(n_132), .B(n_188), .C(n_251), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_72), .Y(n_196) );
INVx1_ASAP7_75t_L g704 ( .A(n_73), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_74), .A2(n_124), .B(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_75), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_76), .A2(n_124), .B(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_77), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_78), .A2(n_123), .B(n_454), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_79), .Y(n_477) );
INVx1_ASAP7_75t_L g525 ( .A(n_80), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_81), .B(n_140), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_82), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_83), .A2(n_124), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g528 ( .A(n_84), .Y(n_528) );
INVx2_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
INVx1_ASAP7_75t_L g495 ( .A(n_86), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_87), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_88), .B(n_170), .Y(n_223) );
OR2x2_ASAP7_75t_L g110 ( .A(n_89), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g429 ( .A(n_89), .Y(n_429) );
OR2x2_ASAP7_75t_L g708 ( .A(n_89), .B(n_694), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_90), .A2(n_132), .B(n_188), .C(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_91), .B(n_124), .Y(n_181) );
INVx1_ASAP7_75t_L g185 ( .A(n_92), .Y(n_185) );
INVxp67_ASAP7_75t_L g201 ( .A(n_93), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_94), .B(n_157), .Y(n_508) );
INVx1_ASAP7_75t_L g218 ( .A(n_95), .Y(n_218) );
INVx1_ASAP7_75t_L g252 ( .A(n_96), .Y(n_252) );
INVx2_ASAP7_75t_L g516 ( .A(n_97), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_98), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g213 ( .A(n_99), .B(n_146), .Y(n_213) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_114), .B1(n_428), .B2(n_430), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g696 ( .A(n_109), .Y(n_696) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g428 ( .A(n_111), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g694 ( .A(n_111), .Y(n_694) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_114), .A2(n_712), .B1(n_715), .B2(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_114), .Y(n_715) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g695 ( .A1(n_115), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
AND2x2_ASAP7_75t_SL g115 ( .A(n_116), .B(n_364), .Y(n_115) );
NOR5xp2_ASAP7_75t_L g116 ( .A(n_117), .B(n_295), .C(n_324), .D(n_344), .E(n_351), .Y(n_116) );
OAI211xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_175), .B(n_239), .C(n_282), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_119), .A2(n_367), .B1(n_369), .B2(n_370), .Y(n_366) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_154), .Y(n_119) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_120), .Y(n_242) );
AND2x4_ASAP7_75t_L g275 ( .A(n_120), .B(n_276), .Y(n_275) );
INVx5_ASAP7_75t_L g293 ( .A(n_120), .Y(n_293) );
AND2x2_ASAP7_75t_L g302 ( .A(n_120), .B(n_294), .Y(n_302) );
AND2x2_ASAP7_75t_L g314 ( .A(n_120), .B(n_179), .Y(n_314) );
AND2x2_ASAP7_75t_L g410 ( .A(n_120), .B(n_278), .Y(n_410) );
OR2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_151), .Y(n_120) );
AOI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_131), .B(n_144), .Y(n_121) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_125), .B(n_129), .Y(n_219) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g142 ( .A(n_126), .Y(n_142) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
INVx1_ASAP7_75t_L g226 ( .A(n_127), .Y(n_226) );
INVx1_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_128), .Y(n_138) );
INVx3_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
INVx1_ASAP7_75t_L g237 ( .A(n_128), .Y(n_237) );
BUFx3_ASAP7_75t_L g143 ( .A(n_129), .Y(n_143) );
INVx4_ASAP7_75t_SL g173 ( .A(n_129), .Y(n_173) );
INVx5_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx3_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_133), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B(n_141), .Y(n_135) );
INVx2_ASAP7_75t_L g140 ( .A(n_137), .Y(n_140) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_140), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_140), .A2(n_187), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_140), .A2(n_444), .B(n_445), .C(n_446), .Y(n_443) );
O2A1O1Ixp5_ASAP7_75t_L g494 ( .A1(n_140), .A2(n_446), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_141), .A2(n_165), .B(n_480), .C(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_142), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_145), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g153 ( .A(n_146), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_146), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_146), .A2(n_208), .B(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_146), .A2(n_219), .B(n_477), .C(n_478), .Y(n_476) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_146), .A2(n_501), .B(n_508), .Y(n_500) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x2_ASAP7_75t_L g158 ( .A(n_147), .B(n_148), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_153), .A2(n_491), .B(n_497), .Y(n_490) );
INVx2_ASAP7_75t_L g276 ( .A(n_154), .Y(n_276) );
AND2x2_ASAP7_75t_L g294 ( .A(n_154), .B(n_248), .Y(n_294) );
AND2x2_ASAP7_75t_L g313 ( .A(n_154), .B(n_247), .Y(n_313) );
AND2x2_ASAP7_75t_L g353 ( .A(n_154), .B(n_293), .Y(n_353) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_159), .B(n_174), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_156), .B(n_190), .Y(n_189) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_156), .A2(n_217), .B(n_227), .Y(n_216) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_156), .A2(n_249), .B(n_257), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_156), .B(n_258), .Y(n_257) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_156), .A2(n_440), .B(n_447), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_156), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_156), .B(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_233), .B(n_234), .Y(n_232) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_SL g160 ( .A1(n_161), .A2(n_162), .B(n_163), .C(n_173), .Y(n_160) );
INVx2_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_162), .A2(n_173), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_162), .A2(n_173), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_162), .A2(n_173), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_162), .A2(n_173), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g512 ( .A1(n_162), .A2(n_173), .B(n_513), .C(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_162), .A2(n_173), .B(n_525), .C(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_165), .B(n_201), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_165), .A2(n_199), .B1(n_458), .B2(n_459), .Y(n_457) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_166), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_169), .B(n_471), .Y(n_470) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g505 ( .A(n_170), .Y(n_505) );
INVx2_ASAP7_75t_L g446 ( .A(n_171), .Y(n_446) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
INVx1_ASAP7_75t_L g529 ( .A(n_172), .Y(n_529) );
INVx1_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
INVxp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_203), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI322xp5_ASAP7_75t_L g412 ( .A1(n_178), .A2(n_214), .A3(n_267), .B1(n_275), .B2(n_329), .C1(n_413), .C2(n_416), .Y(n_412) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
INVx5_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
AND2x2_ASAP7_75t_L g261 ( .A(n_179), .B(n_246), .Y(n_261) );
BUFx2_ASAP7_75t_L g339 ( .A(n_179), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_179), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g416 ( .A(n_179), .B(n_323), .Y(n_416) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_189), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_191), .B(n_205), .Y(n_270) );
INVx1_ASAP7_75t_L g297 ( .A(n_191), .Y(n_297) );
AND2x2_ASAP7_75t_L g310 ( .A(n_191), .B(n_230), .Y(n_310) );
AND2x2_ASAP7_75t_L g411 ( .A(n_191), .B(n_329), .Y(n_411) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g265 ( .A(n_192), .B(n_205), .Y(n_265) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_192), .Y(n_273) );
OR2x2_ASAP7_75t_L g280 ( .A(n_192), .B(n_230), .Y(n_280) );
AND2x2_ASAP7_75t_L g290 ( .A(n_192), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_192), .B(n_216), .Y(n_319) );
INVxp67_ASAP7_75t_L g343 ( .A(n_192), .Y(n_343) );
AND2x2_ASAP7_75t_L g350 ( .A(n_192), .B(n_214), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_192), .B(n_230), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_192), .B(n_215), .Y(n_376) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_202), .Y(n_192) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_193), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_193), .A2(n_511), .B(n_517), .Y(n_510) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_193), .A2(n_523), .B(n_530), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_198), .A2(n_252), .B(n_253), .C(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_199), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_199), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_214), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_205), .B(n_231), .Y(n_320) );
OR2x2_ASAP7_75t_L g342 ( .A(n_205), .B(n_215), .Y(n_342) );
AND2x2_ASAP7_75t_L g355 ( .A(n_205), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_205), .B(n_310), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_205), .A2(n_366), .B(n_371), .C(n_380), .Y(n_365) );
AND2x2_ASAP7_75t_L g426 ( .A(n_205), .B(n_230), .Y(n_426) );
INVx5_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g279 ( .A(n_206), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_206), .B(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_206), .B(n_274), .Y(n_286) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
OR2x2_ASAP7_75t_L g299 ( .A(n_206), .B(n_215), .Y(n_299) );
AND2x2_ASAP7_75t_SL g304 ( .A(n_206), .B(n_290), .Y(n_304) );
AND2x2_ASAP7_75t_L g329 ( .A(n_206), .B(n_215), .Y(n_329) );
AND2x2_ASAP7_75t_L g349 ( .A(n_206), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g387 ( .A(n_206), .B(n_214), .Y(n_387) );
OR2x2_ASAP7_75t_L g390 ( .A(n_206), .B(n_376), .Y(n_390) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_213), .Y(n_206) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_230), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_215), .A2(n_334), .B(n_337), .C(n_343), .Y(n_333) );
INVx5_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_216), .B(n_230), .Y(n_264) );
AND2x2_ASAP7_75t_L g268 ( .A(n_216), .B(n_231), .Y(n_268) );
OR2x2_ASAP7_75t_L g274 ( .A(n_216), .B(n_230), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_219), .A2(n_441), .B(n_442), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_219), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_224), .A2(n_236), .B(n_238), .Y(n_235) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g451 ( .A(n_229), .Y(n_451) );
INVx1_ASAP7_75t_SL g291 ( .A(n_230), .Y(n_291) );
OR2x2_ASAP7_75t_L g419 ( .A(n_230), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_259), .B(n_262), .C(n_271), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AOI31xp33_ASAP7_75t_L g344 ( .A1(n_241), .A2(n_345), .A3(n_347), .B(n_348), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_242), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_243), .B(n_275), .Y(n_281) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_244), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g301 ( .A(n_244), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g306 ( .A(n_244), .B(n_276), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_244), .B(n_275), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_244), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g336 ( .A(n_244), .B(n_293), .Y(n_336) );
AND2x2_ASAP7_75t_L g341 ( .A(n_244), .B(n_313), .Y(n_341) );
OR2x2_ASAP7_75t_L g360 ( .A(n_244), .B(n_246), .Y(n_360) );
OR2x2_ASAP7_75t_L g362 ( .A(n_244), .B(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_244), .Y(n_409) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g309 ( .A(n_246), .B(n_276), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_246), .B(n_293), .Y(n_332) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g278 ( .A(n_248), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_256), .Y(n_249) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g472 ( .A(n_255), .Y(n_472) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g369 ( .A(n_261), .B(n_293), .Y(n_369) );
AOI322xp5_ASAP7_75t_L g371 ( .A1(n_261), .A2(n_275), .A3(n_313), .B1(n_372), .B2(n_373), .C1(n_374), .C2(n_377), .Y(n_371) );
INVx1_ASAP7_75t_L g379 ( .A(n_261), .Y(n_379) );
NAND2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_SL g373 ( .A(n_263), .Y(n_373) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
OR2x2_ASAP7_75t_L g325 ( .A(n_264), .B(n_270), .Y(n_325) );
INVx1_ASAP7_75t_L g356 ( .A(n_264), .Y(n_356) );
INVx2_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI32xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_275), .A3(n_277), .B1(n_279), .B2(n_281), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AOI21xp33_ASAP7_75t_SL g311 ( .A1(n_274), .A2(n_289), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g326 ( .A(n_275), .Y(n_326) );
AND2x4_ASAP7_75t_L g323 ( .A(n_276), .B(n_293), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_276), .B(n_359), .Y(n_358) );
AOI322xp5_ASAP7_75t_L g388 ( .A1(n_277), .A2(n_304), .A3(n_323), .B1(n_356), .B2(n_389), .C1(n_391), .C2(n_392), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_277), .A2(n_354), .B1(n_418), .B2(n_419), .C(n_421), .Y(n_417) );
AND2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g285 ( .A(n_280), .Y(n_285) );
OR2x2_ASAP7_75t_L g357 ( .A(n_280), .B(n_342), .Y(n_357) );
OAI31xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_286), .A3(n_287), .B(n_292), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_316), .B1(n_317), .B2(n_321), .Y(n_315) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_287), .A2(n_328), .B1(n_381), .B2(n_384), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g370 ( .A(n_290), .B(n_339), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_290), .B(n_329), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_291), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g404 ( .A(n_291), .B(n_342), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_292), .A2(n_387), .B1(n_400), .B2(n_403), .Y(n_399) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g308 ( .A(n_293), .Y(n_308) );
AND2x2_ASAP7_75t_L g391 ( .A(n_293), .B(n_313), .Y(n_391) );
OR2x2_ASAP7_75t_L g393 ( .A(n_293), .B(n_360), .Y(n_393) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_293), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_294), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_294), .B(n_339), .Y(n_347) );
OAI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B(n_303), .C(n_315), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_307), .B2(n_310), .C(n_311), .Y(n_303) );
INVxp67_ASAP7_75t_L g415 ( .A(n_306), .Y(n_415) );
INVx1_ASAP7_75t_L g382 ( .A(n_307), .Y(n_382) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g346 ( .A(n_308), .B(n_313), .Y(n_346) );
INVx1_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_309), .B(n_336), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g378 ( .A(n_313), .Y(n_378) );
AND2x2_ASAP7_75t_L g384 ( .A(n_313), .B(n_339), .Y(n_384) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_SL g372 ( .A(n_320), .Y(n_372) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_323), .B(n_359), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_327), .B2(n_330), .C(n_333), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g420 ( .A(n_329), .Y(n_420) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g338 ( .A(n_332), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_336), .B(n_395), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_342), .Y(n_337) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_340), .A2(n_386), .B(n_388), .C(n_394), .Y(n_385) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g397 ( .A(n_342), .Y(n_397) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI222xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B1(n_357), .B2(n_358), .C1(n_361), .C2(n_362), .Y(n_351) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g427 ( .A(n_358), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_359), .B(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_359), .A2(n_406), .B1(n_408), .B2(n_411), .Y(n_405) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NOR4xp25_ASAP7_75t_L g364 ( .A(n_365), .B(n_385), .C(n_398), .D(n_417), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_367), .B(n_397), .Y(n_407) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g374 ( .A(n_372), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_375), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_405), .C(n_412), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx2_ASAP7_75t_L g414 ( .A(n_410), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_424), .B(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g699 ( .A(n_428), .Y(n_699) );
NOR2x2_ASAP7_75t_L g693 ( .A(n_429), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g697 ( .A(n_430), .Y(n_697) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_625), .Y(n_430) );
NAND5xp2_ASAP7_75t_L g431 ( .A(n_432), .B(n_554), .C(n_584), .D(n_605), .E(n_611), .Y(n_431) );
AOI221xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_487), .B1(n_518), .B2(n_520), .C(n_531), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_484), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_462), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_SL g605 ( .A1(n_437), .A2(n_474), .B(n_606), .C(n_609), .Y(n_605) );
AND2x2_ASAP7_75t_L g675 ( .A(n_437), .B(n_475), .Y(n_675) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_449), .Y(n_437) );
AND2x2_ASAP7_75t_L g533 ( .A(n_438), .B(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g537 ( .A(n_438), .B(n_534), .Y(n_537) );
OR2x2_ASAP7_75t_L g563 ( .A(n_438), .B(n_475), .Y(n_563) );
AND2x2_ASAP7_75t_L g565 ( .A(n_438), .B(n_465), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_438), .B(n_464), .Y(n_583) );
INVx1_ASAP7_75t_L g616 ( .A(n_438), .Y(n_616) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
AND2x2_ASAP7_75t_L g519 ( .A(n_439), .B(n_465), .Y(n_519) );
AND2x2_ASAP7_75t_L g672 ( .A(n_439), .B(n_475), .Y(n_672) );
AND2x2_ASAP7_75t_L g553 ( .A(n_449), .B(n_463), .Y(n_553) );
OR2x2_ASAP7_75t_L g557 ( .A(n_449), .B(n_475), .Y(n_557) );
AND2x2_ASAP7_75t_L g582 ( .A(n_449), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g629 ( .A(n_449), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_449), .B(n_591), .Y(n_677) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B(n_460), .Y(n_449) );
INVx1_ASAP7_75t_L g535 ( .A(n_450), .Y(n_535) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_453), .A2(n_461), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI322xp33_ASAP7_75t_L g678 ( .A1(n_462), .A2(n_614), .A3(n_637), .B1(n_658), .B2(n_679), .C1(n_681), .C2(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_463), .B(n_534), .Y(n_681) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
AND2x2_ASAP7_75t_L g485 ( .A(n_464), .B(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g550 ( .A(n_464), .B(n_475), .Y(n_550) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g591 ( .A(n_465), .B(n_475), .Y(n_591) );
AND2x2_ASAP7_75t_L g635 ( .A(n_465), .B(n_474), .Y(n_635) );
AND2x2_ASAP7_75t_L g518 ( .A(n_474), .B(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g536 ( .A(n_474), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_474), .B(n_565), .Y(n_689) );
INVx3_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g484 ( .A(n_475), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_475), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g603 ( .A(n_475), .B(n_534), .Y(n_603) );
AND2x2_ASAP7_75t_L g630 ( .A(n_475), .B(n_565), .Y(n_630) );
OR2x2_ASAP7_75t_L g686 ( .A(n_475), .B(n_537), .Y(n_686) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
INVx1_ASAP7_75t_SL g572 ( .A(n_484), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_485), .B(n_603), .Y(n_604) );
AND2x2_ASAP7_75t_L g638 ( .A(n_485), .B(n_628), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_485), .B(n_561), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_485), .B(n_683), .Y(n_682) );
OAI31xp33_ASAP7_75t_L g656 ( .A1(n_487), .A2(n_518), .A3(n_657), .B(n_659), .Y(n_656) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_499), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_488), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g639 ( .A(n_488), .B(n_574), .Y(n_639) );
OR2x2_ASAP7_75t_L g646 ( .A(n_488), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g658 ( .A(n_488), .B(n_547), .Y(n_658) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g592 ( .A(n_489), .B(n_593), .Y(n_592) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g520 ( .A(n_490), .B(n_521), .Y(n_520) );
INVx4_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
AND2x2_ASAP7_75t_L g578 ( .A(n_490), .B(n_522), .Y(n_578) );
AND2x2_ASAP7_75t_L g577 ( .A(n_499), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g647 ( .A(n_499), .Y(n_647) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_500), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g547 ( .A(n_500), .B(n_510), .Y(n_547) );
INVx2_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
AND2x2_ASAP7_75t_L g581 ( .A(n_500), .B(n_510), .Y(n_581) );
AND2x2_ASAP7_75t_L g588 ( .A(n_500), .B(n_544), .Y(n_588) );
BUFx3_ASAP7_75t_L g598 ( .A(n_500), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_500), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g543 ( .A(n_509), .Y(n_543) );
AND2x2_ASAP7_75t_L g551 ( .A(n_509), .B(n_541), .Y(n_551) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g521 ( .A(n_510), .B(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_510), .Y(n_575) );
INVx2_ASAP7_75t_SL g558 ( .A(n_519), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_519), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_519), .B(n_628), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_520), .B(n_598), .Y(n_651) );
INVx1_ASAP7_75t_SL g685 ( .A(n_520), .Y(n_685) );
INVx1_ASAP7_75t_SL g593 ( .A(n_521), .Y(n_593) );
INVx1_ASAP7_75t_SL g544 ( .A(n_522), .Y(n_544) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_522), .Y(n_555) );
OR2x2_ASAP7_75t_L g566 ( .A(n_522), .B(n_541), .Y(n_566) );
AND2x2_ASAP7_75t_L g580 ( .A(n_522), .B(n_541), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_522), .B(n_570), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_536), .B(n_538), .C(n_549), .Y(n_531) );
AOI31xp33_ASAP7_75t_L g648 ( .A1(n_532), .A2(n_649), .A3(n_650), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g621 ( .A(n_533), .B(n_550), .Y(n_621) );
BUFx3_ASAP7_75t_L g561 ( .A(n_534), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_534), .B(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g597 ( .A(n_534), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_534), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g552 ( .A(n_537), .Y(n_552) );
OAI222xp33_ASAP7_75t_L g661 ( .A1(n_537), .A2(n_662), .B1(n_665), .B2(n_666), .C1(n_667), .C2(n_668), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
INVx1_ASAP7_75t_L g667 ( .A(n_539), .Y(n_667) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_541), .B(n_544), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_541), .B(n_567), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_541), .B(n_542), .Y(n_637) );
INVx1_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_542), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g690 ( .A(n_542), .Y(n_690) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g570 ( .A(n_543), .Y(n_570) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
AOI32xp33_ASAP7_75t_L g549 ( .A1(n_545), .A2(n_550), .A3(n_551), .B1(n_552), .B2(n_553), .Y(n_549) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_547), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g624 ( .A(n_547), .Y(n_624) );
OR2x2_ASAP7_75t_L g665 ( .A(n_547), .B(n_566), .Y(n_665) );
INVx1_ASAP7_75t_L g601 ( .A(n_548), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_550), .B(n_561), .Y(n_586) );
INVx3_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g611 ( .A1(n_550), .A2(n_595), .A3(n_612), .B1(n_614), .B2(n_617), .C1(n_621), .C2(n_622), .Y(n_611) );
AND2x2_ASAP7_75t_L g587 ( .A(n_551), .B(n_588), .Y(n_587) );
INVxp67_ASAP7_75t_L g664 ( .A(n_551), .Y(n_664) );
A2O1A1O1Ixp25_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_559), .C(n_567), .D(n_568), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_555), .B(n_598), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_557), .A2(n_569), .B1(n_572), .B2(n_573), .C(n_576), .Y(n_568) );
INVx1_ASAP7_75t_SL g683 ( .A(n_557), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B(n_566), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_561), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_563), .A2(n_647), .B1(n_654), .B2(n_655), .C(n_656), .Y(n_653) );
OAI222xp33_ASAP7_75t_L g684 ( .A1(n_564), .A2(n_685), .B1(n_686), .B2(n_687), .C1(n_689), .C2(n_690), .Y(n_684) );
AND2x2_ASAP7_75t_L g642 ( .A(n_565), .B(n_628), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_565), .A2(n_580), .B(n_627), .Y(n_654) );
INVx1_ASAP7_75t_L g668 ( .A(n_565), .Y(n_668) );
INVx2_ASAP7_75t_SL g571 ( .A(n_566), .Y(n_571) );
AND2x2_ASAP7_75t_L g574 ( .A(n_567), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_SL g608 ( .A(n_570), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_570), .B(n_580), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_571), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_571), .B(n_581), .Y(n_610) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_579), .B(n_582), .Y(n_576) );
INVx1_ASAP7_75t_SL g594 ( .A(n_578), .Y(n_594) );
AND2x2_ASAP7_75t_L g641 ( .A(n_578), .B(n_624), .Y(n_641) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AND2x2_ASAP7_75t_L g680 ( .A(n_580), .B(n_598), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_581), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g666 ( .A(n_582), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B1(n_589), .B2(n_596), .C(n_599), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B1(n_594), .B2(n_595), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_593), .A2(n_600), .B1(n_602), .B2(n_604), .Y(n_599) );
OR2x2_ASAP7_75t_L g670 ( .A(n_594), .B(n_598), .Y(n_670) );
OR2x2_ASAP7_75t_L g673 ( .A(n_594), .B(n_608), .Y(n_673) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_615), .A2(n_670), .B1(n_671), .B2(n_673), .C(n_674), .Y(n_669) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_640), .C(n_652), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_631), .B1(n_633), .B2(n_636), .C1(n_638), .C2(n_639), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_628), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g650 ( .A(n_630), .Y(n_650) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_645), .C(n_648), .Y(n_640) );
INVx1_ASAP7_75t_L g655 ( .A(n_641), .Y(n_655) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR5xp2_ASAP7_75t_L g652 ( .A(n_653), .B(n_661), .C(n_669), .D(n_678), .E(n_684), .Y(n_652) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .Y(n_701) );
NOR2xp33_ASAP7_75t_SL g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_SL g726 ( .A(n_703), .Y(n_726) );
INVx1_ASAP7_75t_L g725 ( .A(n_705), .Y(n_725) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_705), .A2(n_726), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_708), .Y(n_717) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_708), .Y(n_720) );
BUFx2_ASAP7_75t_L g729 ( .A(n_708), .Y(n_729) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_717), .B(n_718), .Y(n_710) );
INVx1_ASAP7_75t_L g716 ( .A(n_712), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
endmodule