module fake_ariane_1757_n_1170 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1170);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1170;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_183;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_1154;
wire n_1166;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_162;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_154;
wire n_883;
wire n_338;
wire n_142;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_145;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_731;
wire n_779;
wire n_903;
wire n_871;
wire n_315;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_167;
wire n_422;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_158;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_143;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_1107;
wire n_173;
wire n_989;
wire n_242;
wire n_645;
wire n_858;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_1134;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_600;
wire n_433;
wire n_721;
wire n_840;
wire n_481;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_1099;
wire n_271;
wire n_1153;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_1074;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_163;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_977;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1144;
wire n_149;
wire n_838;
wire n_623;
wire n_383;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_616;
wire n_658;
wire n_705;
wire n_630;
wire n_617;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_1135;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_673;
wire n_452;
wire n_1114;
wire n_676;
wire n_178;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_171;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_697;
wire n_274;
wire n_437;
wire n_622;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_156;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1148;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_159;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_608;
wire n_959;
wire n_494;
wire n_892;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_165;
wire n_1037;
wire n_144;
wire n_981;
wire n_1010;
wire n_1110;
wire n_990;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_815;
wire n_542;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVxp33_ASAP7_75t_SL g142 ( 
.A(n_65),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_53),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_28),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_82),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_37),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_15),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_110),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_80),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_18),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_109),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_41),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_50),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_62),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_34),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_104),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_79),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_57),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_14),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_95),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_125),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_44),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_40),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_27),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_108),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_32),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_134),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_151),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_173),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_160),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_175),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_169),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_202),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_208),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_199),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_224),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_197),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_202),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_202),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_202),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_202),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_209),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g275 ( 
.A(n_231),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_231),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_250),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_226),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_232),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_251),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_250),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_229),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_248),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_235),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_244),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_241),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_253),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_260),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_306),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_278),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_277),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_308),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_277),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_285),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_313),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_285),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_315),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_R g345 ( 
.A(n_317),
.B(n_262),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_315),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_263),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_317),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_283),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_294),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_283),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_287),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_287),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_303),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_292),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_297),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_275),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_327),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_321),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_362),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_345),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_324),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_310),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_335),
.A2(n_312),
.B1(n_311),
.B2(n_305),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_328),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_331),
.B(n_164),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_320),
.Y(n_379)
);

XNOR2x2_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_249),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_333),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

NOR2x1_ASAP7_75t_L g386 ( 
.A(n_322),
.B(n_257),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_351),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

BUFx8_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_264),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_301),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_350),
.B(n_275),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_267),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_297),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_314),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_300),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_329),
.B(n_300),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_329),
.B(n_269),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

BUFx8_ASAP7_75t_SL g409 ( 
.A(n_343),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_346),
.A2(n_309),
.B(n_167),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_316),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_259),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_330),
.B(n_307),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_349),
.B(n_247),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_359),
.B(n_164),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_345),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_345),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_321),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_326),
.B(n_246),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_347),
.B(n_248),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_246),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_330),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_325),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_322),
.B(n_165),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_325),
.A2(n_156),
.B(n_153),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_345),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_347),
.B(n_248),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_325),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_325),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_325),
.A2(n_176),
.B(n_159),
.Y(n_437)
);

BUFx8_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_349),
.A2(n_249),
.B1(n_142),
.B2(n_172),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_432),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_365),
.B(n_274),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_142),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_367),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_172),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_370),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_366),
.B(n_191),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_366),
.B(n_389),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_382),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_384),
.B(n_191),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

BUFx8_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_417),
.B(n_174),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_428),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_420),
.B(n_427),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_420),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_427),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_389),
.B(n_192),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_435),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_192),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_379),
.B(n_195),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_419),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_379),
.B(n_181),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_375),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_379),
.B(n_181),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_483),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_461),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_461),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_461),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_448),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_457),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_479),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_466),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_457),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_465),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_465),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_442),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_462),
.Y(n_501)
);

HB1xp67_ASAP7_75t_SL g502 ( 
.A(n_480),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_475),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_R g504 ( 
.A(n_446),
.B(n_371),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_441),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_446),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_463),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_441),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_449),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_458),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_460),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_482),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_467),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_R g516 ( 
.A(n_450),
.B(n_371),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_467),
.B(n_368),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_444),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_463),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_463),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_388),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_495),
.A2(n_378),
.B1(n_380),
.B2(n_410),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_506),
.A2(n_404),
.B1(n_439),
.B2(n_364),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_502),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_490),
.B(n_441),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_487),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_447),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_523),
.A2(n_392),
.B1(n_399),
.B2(n_405),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_513),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_406),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_517),
.Y(n_535)
);

AND3x2_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_484),
.C(n_482),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_447),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_519),
.Y(n_539)
);

INVxp33_ASAP7_75t_SL g540 ( 
.A(n_486),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_518),
.B(n_441),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_515),
.B(n_459),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_499),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_521),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_503),
.B(n_406),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_493),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_496),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_497),
.B(n_484),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_508),
.B(n_445),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_502),
.B(n_408),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_510),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_505),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_L g556 ( 
.A(n_508),
.B(n_416),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_505),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_504),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_487),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_512),
.B(n_445),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_505),
.B(n_459),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_522),
.B(n_456),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_512),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_512),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_512),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_520),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_514),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_488),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_489),
.B(n_456),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_491),
.B(n_408),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_516),
.Y(n_573)
);

AO21x2_ASAP7_75t_L g574 ( 
.A1(n_519),
.A2(n_468),
.B(n_464),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_490),
.B(n_445),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_519),
.A2(n_468),
.B(n_464),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_500),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_486),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_496),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_490),
.B(n_424),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_500),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_500),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_496),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_500),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_500),
.Y(n_587)
);

OAI21xp33_ASAP7_75t_SL g588 ( 
.A1(n_490),
.A2(n_477),
.B(n_459),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_490),
.B(n_445),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_496),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_500),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_490),
.B(n_445),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_490),
.B(n_434),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_485),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_504),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_486),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_485),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_490),
.B(n_469),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_515),
.B(n_378),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_490),
.B(n_397),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_490),
.B(n_469),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_487),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_485),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_490),
.B(n_451),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_600),
.A2(n_400),
.B1(n_398),
.B2(n_396),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_573),
.B(n_393),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_574),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_601),
.B(n_388),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_376),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_558),
.B(n_418),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_574),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_576),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_537),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_527),
.B(n_484),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_596),
.B(n_368),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_545),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_527),
.B(n_548),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_595),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_582),
.B(n_470),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_582),
.B(n_470),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_529),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_581),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_543),
.B(n_477),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_533),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_543),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_598),
.Y(n_630)
);

INVx3_ASAP7_75t_R g631 ( 
.A(n_569),
.Y(n_631)
);

NOR2x1p5_ASAP7_75t_L g632 ( 
.A(n_580),
.B(n_407),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_581),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_524),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_594),
.B(n_472),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_604),
.Y(n_636)
);

NAND3x1_ASAP7_75t_L g637 ( 
.A(n_553),
.B(n_407),
.C(n_402),
.Y(n_637)
);

NOR2x1p5_ASAP7_75t_L g638 ( 
.A(n_580),
.B(n_403),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_543),
.B(n_477),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_600),
.B(n_410),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_585),
.B(n_393),
.Y(n_642)
);

NOR2x1p5_ASAP7_75t_L g643 ( 
.A(n_570),
.B(n_403),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_541),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_544),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_597),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_553),
.B(n_401),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_594),
.B(n_472),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_597),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_576),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_531),
.B(n_401),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_599),
.B(n_602),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_532),
.B(n_376),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_549),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_577),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_526),
.A2(n_418),
.B1(n_433),
.B2(n_421),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_534),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_549),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_590),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_540),
.B(n_422),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_393),
.Y(n_664)
);

AND2x6_ASAP7_75t_SL g665 ( 
.A(n_572),
.B(n_546),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_538),
.B(n_476),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_545),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

BUFx6f_ASAP7_75t_SL g670 ( 
.A(n_568),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_534),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_583),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_565),
.B(n_451),
.Y(n_673)
);

AND2x4_ASAP7_75t_SL g674 ( 
.A(n_561),
.B(n_422),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_R g675 ( 
.A(n_536),
.B(n_421),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_584),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_588),
.B(n_525),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_586),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_587),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_549),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_591),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_578),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_578),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_571),
.B(n_454),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_578),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_606),
.Y(n_686)
);

INVxp67_ASAP7_75t_SL g687 ( 
.A(n_528),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_563),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_542),
.B(n_369),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_550),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_554),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_689),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_659),
.B(n_546),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_611),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_616),
.B(n_528),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_619),
.B(n_536),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_655),
.B(n_671),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_645),
.Y(n_698)
);

NAND2x1p5_ASAP7_75t_L g699 ( 
.A(n_638),
.B(n_530),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_669),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_612),
.B(n_610),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_675),
.A2(n_525),
.B1(n_572),
.B2(n_556),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_625),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_647),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_633),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_632),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_618),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_622),
.B(n_575),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_642),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_663),
.B(n_369),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_624),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_658),
.B(n_381),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_669),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_623),
.B(n_575),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_635),
.B(n_650),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_688),
.B(n_589),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_634),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_646),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_654),
.B(n_589),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_653),
.B(n_565),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_634),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_631),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_620),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_621),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_630),
.B(n_593),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_634),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_636),
.B(n_593),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_639),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_677),
.A2(n_547),
.B1(n_605),
.B2(n_559),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_644),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_642),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_609),
.Y(n_733)
);

AND2x6_ASAP7_75t_L g734 ( 
.A(n_626),
.B(n_530),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_626),
.B(n_579),
.Y(n_735)
);

OAI221xp5_ASAP7_75t_L g736 ( 
.A1(n_607),
.A2(n_430),
.B1(n_395),
.B2(n_386),
.C(n_411),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_657),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_672),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_609),
.A2(n_547),
.B1(n_605),
.B2(n_557),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_667),
.B(n_555),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_687),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_613),
.B(n_381),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_639),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_620),
.B(n_578),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_608),
.B(n_179),
.C(n_178),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_676),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_614),
.A2(n_542),
.B1(n_566),
.B2(n_425),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_661),
.B(n_372),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_639),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_681),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_684),
.B(n_564),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_651),
.B(n_395),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_637),
.A2(n_556),
.B1(n_410),
.B2(n_425),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_656),
.B(n_579),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_691),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_614),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_656),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_678),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_629),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_656),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_668),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_615),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_670),
.B(n_433),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_683),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_698),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_698),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_724),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_715),
.B(n_679),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_648),
.B(n_641),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_755),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_719),
.B(n_686),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_701),
.A2(n_689),
.B1(n_643),
.B2(n_664),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_708),
.B(n_666),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_692),
.B(n_683),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_714),
.B(n_665),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_692),
.B(n_683),
.Y(n_776)
);

AND2x2_ASAP7_75t_SL g777 ( 
.A(n_696),
.B(n_674),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_763),
.B(n_670),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_704),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_707),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_693),
.B(n_627),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_724),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_736),
.B(n_680),
.C(n_627),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_705),
.B(n_409),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_700),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_713),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_705),
.Y(n_787)
);

AO22x1_ASAP7_75t_L g788 ( 
.A1(n_692),
.A2(n_390),
.B1(n_617),
.B2(n_438),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_703),
.B(n_409),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_SL g790 ( 
.A(n_722),
.B(n_649),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_759),
.B(n_680),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_706),
.B(n_640),
.Y(n_792)
);

NOR3x1_ASAP7_75t_L g793 ( 
.A(n_741),
.B(n_474),
.C(n_390),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_718),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_695),
.B(n_741),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_738),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_716),
.B(n_685),
.Y(n_797)
);

XNOR2xp5_ASAP7_75t_L g798 ( 
.A(n_720),
.B(n_423),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_740),
.B(n_615),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_725),
.B(n_685),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_727),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_730),
.A2(n_560),
.B(n_552),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_751),
.B(n_640),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_746),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_761),
.B(n_673),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_758),
.B(n_652),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_696),
.B(n_664),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_752),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_723),
.B(n_649),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_744),
.B(n_673),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_694),
.B(n_673),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_709),
.B(n_673),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_706),
.B(n_660),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_733),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_733),
.B(n_652),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_711),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_732),
.B(n_660),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_710),
.B(n_748),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_756),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_742),
.B(n_712),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_707),
.B(n_699),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_734),
.B(n_662),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_734),
.B(n_662),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_734),
.B(n_682),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_735),
.B(n_682),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_754),
.B(n_592),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_717),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_756),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_735),
.B(n_564),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_730),
.A2(n_560),
.B(n_552),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_747),
.B(n_690),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_762),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_762),
.B(n_592),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_717),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_721),
.B(n_561),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_728),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_721),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_739),
.A2(n_561),
.B(n_603),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_731),
.B(n_603),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_737),
.B(n_454),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_818),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_787),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_801),
.B(n_739),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_795),
.B(n_726),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_787),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_815),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_779),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_814),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_781),
.B(n_726),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_820),
.B(n_729),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_775),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_777),
.Y(n_853)
);

INVx8_ASAP7_75t_L g854 ( 
.A(n_780),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_819),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_828),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_827),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_803),
.B(n_729),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_832),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_765),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_799),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_780),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_806),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_766),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_790),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_780),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_838),
.Y(n_867)
);

AND2x2_ASAP7_75t_SL g868 ( 
.A(n_793),
.B(n_702),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_767),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_835),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_782),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_802),
.A2(n_753),
.B(n_745),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_830),
.A2(n_750),
.B(n_437),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_791),
.B(n_743),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_831),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_785),
.Y(n_876)
);

NAND2x1p5_ASAP7_75t_L g877 ( 
.A(n_774),
.B(n_743),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_789),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_838),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_786),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_807),
.B(n_822),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_797),
.B(n_749),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_794),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_770),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_773),
.B(n_749),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_796),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_808),
.B(n_804),
.Y(n_888)
);

INVxp33_ASAP7_75t_L g889 ( 
.A(n_778),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_784),
.Y(n_890)
);

AND2x2_ASAP7_75t_SL g891 ( 
.A(n_793),
.B(n_783),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_836),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_834),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_837),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_836),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_811),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_823),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_891),
.A2(n_839),
.B(n_813),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_861),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_889),
.B(n_772),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_848),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_891),
.A2(n_792),
.B(n_824),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_891),
.A2(n_868),
.B(n_872),
.C(n_852),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_868),
.A2(n_805),
.B1(n_769),
.B2(n_807),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_888),
.B(n_768),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_846),
.B(n_821),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_856),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_888),
.B(n_800),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_857),
.B(n_809),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_893),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_868),
.A2(n_833),
.B1(n_825),
.B2(n_826),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_860),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_844),
.A2(n_840),
.B(n_771),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_848),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_856),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_865),
.A2(n_776),
.B(n_788),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_875),
.A2(n_841),
.B(n_817),
.C(n_170),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_848),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_846),
.B(n_810),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_843),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_842),
.A2(n_798),
.B(n_812),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_853),
.B(n_757),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_851),
.A2(n_760),
.B(n_757),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_860),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_L g925 ( 
.A1(n_875),
.A2(n_871),
.B(n_869),
.C(n_849),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_854),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_897),
.A2(n_764),
.B(n_760),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_846),
.B(n_764),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_883),
.B(n_816),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_897),
.A2(n_471),
.B(n_423),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_883),
.B(n_180),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_886),
.B(n_184),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_853),
.A2(n_454),
.B1(n_481),
.B2(n_452),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_886),
.B(n_876),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_846),
.B(n_0),
.Y(n_935)
);

OAI321xp33_ASAP7_75t_L g936 ( 
.A1(n_877),
.A2(n_143),
.A3(n_170),
.B1(n_193),
.B2(n_196),
.C(n_154),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_881),
.A2(n_473),
.B(n_481),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_843),
.B(n_0),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_881),
.A2(n_481),
.B(n_452),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_881),
.A2(n_854),
.B(n_896),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_864),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_878),
.Y(n_942)
);

BUFx8_ASAP7_75t_L g943 ( 
.A(n_843),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_L g944 ( 
.A(n_887),
.B(n_1),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_853),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_876),
.B(n_1),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_881),
.A2(n_452),
.B(n_451),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_873),
.A2(n_195),
.B(n_150),
.C(n_177),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_862),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_869),
.A2(n_871),
.B(n_849),
.C(n_887),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_870),
.A2(n_431),
.B(n_394),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_864),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_887),
.B(n_2),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_869),
.A2(n_374),
.B(n_373),
.C(n_394),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_856),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_862),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_869),
.A2(n_871),
.B(n_849),
.C(n_885),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_854),
.A2(n_452),
.B(n_451),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_880),
.B(n_2),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_857),
.A2(n_394),
.B(n_416),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_900),
.Y(n_961)
);

OA22x2_ASAP7_75t_L g962 ( 
.A1(n_911),
.A2(n_890),
.B1(n_887),
.B2(n_847),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_903),
.A2(n_854),
.B(n_880),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_945),
.B(n_866),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_898),
.A2(n_854),
.B(n_847),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_943),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_901),
.B(n_862),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_905),
.A2(n_877),
.B1(n_866),
.B2(n_862),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_942),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_909),
.B(n_845),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_901),
.B(n_862),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_899),
.B(n_871),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_920),
.B(n_866),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_934),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_936),
.A2(n_847),
.B(n_855),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_914),
.B(n_879),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_944),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_902),
.A2(n_855),
.B(n_849),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_977),
.A2(n_962),
.B1(n_904),
.B2(n_961),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_963),
.A2(n_940),
.B1(n_916),
.B2(n_908),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_969),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_965),
.A2(n_975),
.B(n_953),
.C(n_978),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_966),
.B(n_918),
.Y(n_983)
);

AO32x1_ASAP7_75t_L g984 ( 
.A1(n_968),
.A2(n_867),
.A3(n_933),
.B1(n_941),
.B2(n_952),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_976),
.A2(n_932),
.B(n_931),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_970),
.A2(n_913),
.B1(n_921),
.B2(n_960),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_967),
.A2(n_917),
.B(n_948),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_974),
.A2(n_925),
.B(n_930),
.C(n_938),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_976),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_972),
.B(n_946),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_971),
.A2(n_959),
.B(n_957),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_973),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_964),
.A2(n_950),
.B(n_935),
.C(n_954),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_973),
.B(n_918),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_964),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_966),
.B(n_943),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_961),
.B(n_912),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_962),
.A2(n_915),
.B1(n_955),
.B2(n_907),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_977),
.A2(n_919),
.B(n_922),
.C(n_906),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_976),
.B(n_922),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_961),
.A2(n_951),
.B(n_910),
.C(n_937),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_966),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_961),
.A2(n_926),
.B(n_929),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_1002),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_981),
.B(n_956),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_981),
.Y(n_1006)
);

AND3x1_ASAP7_75t_SL g1007 ( 
.A(n_992),
.B(n_924),
.C(n_928),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_989),
.B(n_956),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_996),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_989),
.B(n_988),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1010),
.A2(n_982),
.B(n_984),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1004),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_1008),
.A2(n_987),
.B(n_979),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1011),
.A2(n_993),
.B1(n_998),
.B2(n_999),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_1012),
.B(n_1006),
.Y(n_1015)
);

BUFx10_ASAP7_75t_L g1016 ( 
.A(n_1013),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_1014),
.A2(n_1001),
.B(n_1005),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_1015),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_1018),
.A2(n_985),
.B(n_994),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1017),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1020),
.B(n_1016),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_1019),
.B(n_983),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1021),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_1022),
.A2(n_1009),
.B(n_991),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1024),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1025),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1025),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1027),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1027),
.B(n_1026),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1031),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_1030),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_1029),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1034),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1035),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1036),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_1037),
.B(n_1038),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1038),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1039),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1040),
.B(n_989),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_1041),
.B(n_438),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1042),
.B(n_995),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1043),
.B(n_997),
.Y(n_1045)
);

INVxp33_ASAP7_75t_L g1046 ( 
.A(n_1044),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1046),
.B(n_1000),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1045),
.Y(n_1048)
);

XNOR2xp5_ASAP7_75t_L g1049 ( 
.A(n_1046),
.B(n_3),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1049),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1047),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1048),
.B(n_990),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_1051),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_1050),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1053),
.B(n_1052),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1054),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1056),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1055),
.Y(n_1058)
);

OAI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1057),
.A2(n_980),
.B1(n_1003),
.B2(n_1007),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_186),
.B(n_183),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1060),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1059),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_1062),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1061),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1063),
.A2(n_154),
.B1(n_188),
.B2(n_187),
.Y(n_1065)
);

OAI31xp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1063),
.A2(n_189),
.B1(n_190),
.B2(n_154),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1067),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1066),
.B(n_1065),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1067),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1068),
.B(n_956),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1070),
.B(n_949),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_1071),
.B(n_1069),
.Y(n_1073)
);

OAI211xp5_ASAP7_75t_SL g1074 ( 
.A1(n_1072),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1073),
.B(n_154),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_862),
.B1(n_986),
.B2(n_949),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1076),
.A2(n_387),
.B1(n_383),
.B2(n_416),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_6),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1078),
.A2(n_984),
.B(n_7),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_1079),
.B(n_7),
.C(n_8),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1080),
.B(n_8),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_867),
.C(n_9),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_1081),
.A2(n_867),
.B(n_927),
.C(n_11),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_1082),
.B(n_867),
.C(n_9),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1083),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_879),
.Y(n_1087)
);

AOI211xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1084),
.A2(n_923),
.B(n_11),
.C(n_12),
.Y(n_1088)
);

AOI221xp5_ASAP7_75t_L g1089 ( 
.A1(n_1086),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_1089)
);

OAI211xp5_ASAP7_75t_SL g1090 ( 
.A1(n_1087),
.A2(n_10),
.B(n_13),
.C(n_15),
.Y(n_1090)
);

NOR2x1p5_ASAP7_75t_L g1091 ( 
.A(n_1090),
.B(n_1088),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_1089),
.B(n_16),
.C(n_17),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1091),
.Y(n_1093)
);

NOR2x1p5_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_17),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_SL g1095 ( 
.A(n_1093),
.B(n_18),
.C(n_19),
.Y(n_1095)
);

OA211x2_ASAP7_75t_L g1096 ( 
.A1(n_1094),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_20),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_21),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1097),
.B(n_22),
.Y(n_1099)
);

AO22x2_ASAP7_75t_L g1100 ( 
.A1(n_1098),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1100),
.B(n_23),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_1099),
.B(n_895),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_1102),
.B(n_1103),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1101),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1101),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1104),
.A2(n_895),
.B1(n_892),
.B2(n_24),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1105),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1108),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1107),
.A2(n_1106),
.B1(n_895),
.B2(n_892),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_SL g1111 ( 
.A1(n_1109),
.A2(n_895),
.B1(n_892),
.B2(n_879),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1110),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_895),
.B1(n_845),
.B2(n_877),
.Y(n_1113)
);

AOI22x1_ASAP7_75t_L g1114 ( 
.A1(n_1111),
.A2(n_895),
.B1(n_874),
.B2(n_850),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1113),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_1115)
);

XOR2xp5_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_31),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_1116),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1115),
.Y(n_1118)
);

AO21x2_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_874),
.Y(n_1119)
);

OA21x2_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_850),
.B(n_858),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1117),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1117),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_858),
.B(n_882),
.Y(n_1123)
);

AO22x1_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_882),
.B1(n_35),
.B2(n_36),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1119),
.A2(n_947),
.B(n_33),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1120),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1123),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1124),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_SL g1129 ( 
.A(n_1125),
.B(n_1126),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1129),
.B(n_43),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1127),
.A2(n_45),
.B(n_46),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1128),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1129),
.A2(n_51),
.B(n_52),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1129),
.A2(n_54),
.B(n_55),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1129),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1129),
.A2(n_56),
.B(n_58),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1129),
.A2(n_59),
.B(n_60),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1129),
.A2(n_61),
.B(n_63),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1129),
.B(n_64),
.Y(n_1139)
);

XNOR2xp5_ASAP7_75t_L g1140 ( 
.A(n_1129),
.B(n_67),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1129),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1135),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1140),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1131),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_1130),
.B(n_72),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1139),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1141),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1132),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1133),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_1149)
);

BUFx2_ASAP7_75t_SL g1150 ( 
.A(n_1134),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1142),
.A2(n_1138),
.B1(n_1136),
.B2(n_1137),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1143),
.A2(n_939),
.B(n_958),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_R g1153 ( 
.A1(n_1150),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1147),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1146),
.B(n_91),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1144),
.A2(n_863),
.B(n_93),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1145),
.A2(n_92),
.B(n_94),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1151),
.A2(n_1152),
.B(n_1154),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1155),
.A2(n_1148),
.B(n_1149),
.Y(n_1159)
);

AOI221xp5_ASAP7_75t_L g1160 ( 
.A1(n_1153),
.A2(n_859),
.B1(n_863),
.B2(n_98),
.C(n_99),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1156),
.B(n_96),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1159),
.A2(n_1157),
.B1(n_100),
.B2(n_101),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1158),
.A2(n_859),
.B1(n_102),
.B2(n_103),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1162),
.Y(n_1164)
);

AOI22x1_ASAP7_75t_L g1165 ( 
.A1(n_1164),
.A2(n_1163),
.B1(n_1160),
.B2(n_1161),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_859),
.B1(n_106),
.B2(n_107),
.Y(n_1166)
);

AO22x1_ASAP7_75t_L g1167 ( 
.A1(n_1166),
.A2(n_97),
.B1(n_111),
.B2(n_112),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1167),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_1168)
);

AOI211xp5_ASAP7_75t_L g1169 ( 
.A1(n_1168),
.A2(n_894),
.B(n_119),
.C(n_120),
.Y(n_1169)
);

AOI211xp5_ASAP7_75t_L g1170 ( 
.A1(n_1169),
.A2(n_894),
.B(n_884),
.C(n_123),
.Y(n_1170)
);


endmodule