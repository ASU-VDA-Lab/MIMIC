module real_jpeg_1290_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_0),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_0),
.B(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_66),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_44),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_41),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_1),
.B(n_30),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_1),
.B(n_66),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_4),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_4),
.B(n_41),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_9),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_60),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_9),
.B(n_38),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_44),
.Y(n_165)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_10),
.B(n_44),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_10),
.B(n_38),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_10),
.B(n_41),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_11),
.B(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_12),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_12),
.B(n_34),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_14),
.B(n_44),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_14),
.B(n_38),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_142),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_20),
.B(n_105),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_56),
.C(n_71),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_21),
.A2(n_22),
.B1(n_56),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_48),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_23),
.A2(n_24),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_31),
.C(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_29),
.B(n_101),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_32),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_32),
.B(n_82),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_39),
.B(n_48),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.C(n_54),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_51),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_53),
.B(n_101),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_54),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_55),
.B(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_56),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_69),
.C(n_70),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_64),
.C(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_71),
.B(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_94),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_92),
.B2(n_93),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_92),
.C(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_88),
.C(n_90),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_78),
.A2(n_79),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_81),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_87),
.B(n_101),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_99),
.C(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_121),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_133),
.B2(n_134),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_132),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_219),
.B(n_224),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_207),
.B(n_218),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_193),
.B(n_206),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_174),
.B(n_192),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_147),
.B(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.C(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_149),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_150),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_164),
.C(n_168),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_161),
.C(n_162),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_173),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_170),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_183),
.B(n_191),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_179),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.C(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);


endmodule