module fake_jpeg_17127_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_54),
.Y(n_68)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_62),
.B1(n_65),
.B2(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_45),
.B1(n_40),
.B2(n_43),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_49),
.C(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_39),
.B1(n_46),
.B2(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_18),
.B1(n_33),
.B2(n_31),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_59),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_81),
.B(n_12),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_15),
.C(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_88),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_90),
.CI(n_13),
.CON(n_94),
.SN(n_94)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_78),
.B1(n_91),
.B2(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_86),
.C(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_101),
.C(n_97),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_98),
.B(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_95),
.C(n_94),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_14),
.B1(n_20),
.B2(n_23),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_24),
.B(n_25),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_92),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_26),
.Y(n_110)
);


endmodule