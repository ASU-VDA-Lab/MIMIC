module fake_jpeg_7116_n_18 (n_3, n_2, n_1, n_0, n_4, n_5, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_18;

wire n_13;
wire n_11;
wire n_14;
wire n_17;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_7;

AOI22xp5_ASAP7_75t_SL g6 ( 
.A1(n_1),
.A2(n_4),
.B1(n_5),
.B2(n_0),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_6),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

XNOR2x1_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_13),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_3),
.C(n_8),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_15),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_7),
.B(n_15),
.C(n_12),
.Y(n_18)
);


endmodule