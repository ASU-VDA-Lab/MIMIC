module real_jpeg_21476_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_0),
.A2(n_26),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_0),
.A2(n_68),
.B(n_70),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_0),
.B(n_68),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_71),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_0),
.A2(n_10),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_0),
.B(n_141),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_0),
.A2(n_52),
.B(n_55),
.C(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_68),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_3),
.B(n_31),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_179),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_81),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_81),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_81),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_9),
.A2(n_32),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_9),
.A2(n_32),
.B1(n_68),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_35),
.B(n_38),
.C(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_10),
.B(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_122),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_104),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_16),
.B(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.C(n_91),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_17),
.A2(n_18),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.C(n_63),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_19),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_20),
.B(n_33),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_21),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_22),
.B(n_28),
.Y(n_169)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_23),
.A2(n_29),
.B(n_30),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_24),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_26),
.A2(n_36),
.B(n_39),
.C(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_26),
.B(n_34),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_26),
.B(n_30),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_26),
.A2(n_38),
.B(n_57),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_27),
.A2(n_30),
.B(n_131),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_27),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_28),
.B(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_29),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_43),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_34),
.A2(n_96),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_35),
.B(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_35),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_37),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_43),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_45),
.B(n_85),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_45),
.B(n_187),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_50),
.A2(n_60),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_50),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_54),
.B(n_55),
.C(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_52),
.B(n_73),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_53),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_54),
.A2(n_61),
.B(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_58),
.B(n_140),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_59),
.B(n_141),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_59),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_61),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_72),
.B(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_76),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_72),
.B(n_77),
.C(n_78),
.Y(n_76)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_80),
.Y(n_137)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_76),
.B(n_110),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_82),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_90),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_84),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_140),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_105),
.CI(n_121),
.CON(n_104),
.SN(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_94),
.A2(n_99),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_94),
.B(n_214),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_95),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_97),
.B(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_101),
.B(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_104),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_136),
.C(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_116),
.B1(n_138),
.B2(n_139),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_276),
.B(n_282),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_264),
.B(n_275),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_170),
.B(n_246),
.C(n_263),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_159),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_127),
.B(n_159),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_143),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_129),
.B(n_135),
.C(n_143),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_130),
.B(n_133),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_137),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_144),
.Y(n_261)
);

FAx1_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.CI(n_151),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_243),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_162),
.Y(n_243)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_165),
.B(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_166),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_245),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_239),
.B(n_244),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_225),
.B(n_238),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_210),
.B(n_224),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_199),
.B(n_209),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_188),
.B(n_198),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_184),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_193),
.B(n_197),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_201),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_206),
.C(n_208),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_223),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_213),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_227),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_234),
.C(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_234),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_261),
.B2(n_262),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.C(n_262),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_274),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_272),
.C(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);


endmodule