module fake_jpeg_24707_n_60 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_30),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_30),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_7),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_40),
.B(n_41),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_51),
.B1(n_15),
.B2(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_17),
.C(n_18),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_57),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_19),
.C(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_60)
);


endmodule