module fake_jpeg_11810_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_41),
.B(n_51),
.Y(n_97)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_28),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_62),
.Y(n_65)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_0),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_67),
.A2(n_74),
.B1(n_81),
.B2(n_88),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_SL g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_25),
.B1(n_17),
.B2(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_31),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_38),
.B1(n_20),
.B2(n_19),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_39),
.A2(n_38),
.B1(n_20),
.B2(n_19),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_93),
.B1(n_36),
.B2(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_18),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_36),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_33),
.B1(n_37),
.B2(n_30),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_29),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_26),
.B1(n_21),
.B2(n_36),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_61),
.B1(n_52),
.B2(n_49),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_45),
.B1(n_57),
.B2(n_56),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_118),
.B1(n_124),
.B2(n_125),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_60),
.B1(n_21),
.B2(n_26),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_102),
.B1(n_117),
.B2(n_126),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_82),
.B1(n_76),
.B2(n_89),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_14),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_64),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_0),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_36),
.B1(n_48),
.B2(n_3),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_127),
.C(n_71),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_76),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_8),
.B1(n_90),
.B2(n_66),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_116),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_115),
.B1(n_113),
.B2(n_108),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_138),
.B1(n_142),
.B2(n_144),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_108),
.B1(n_107),
.B2(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_127),
.B1(n_99),
.B2(n_91),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_92),
.B1(n_72),
.B2(n_66),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_95),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_73),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_105),
.B1(n_121),
.B2(n_111),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_154),
.B1(n_153),
.B2(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_105),
.Y(n_172)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_128),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_126),
.B1(n_125),
.B2(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_175),
.B1(n_177),
.B2(n_143),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_173),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_91),
.B1(n_112),
.B2(n_119),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_164),
.B1(n_152),
.B2(n_135),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_91),
.B1(n_95),
.B2(n_79),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_170),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_130),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_71),
.B(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_142),
.B1(n_131),
.B2(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_135),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_131),
.B1(n_139),
.B2(n_144),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_130),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_193),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_173),
.C(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_151),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_195),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_155),
.B1(n_159),
.B2(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_178),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_181),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_204),
.B(n_206),
.Y(n_211)
);

AOI22x1_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_161),
.B1(n_164),
.B2(n_157),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_158),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_209),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_174),
.B(n_168),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_212),
.B(n_214),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_196),
.Y(n_224)
);

AOI321xp33_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_193),
.A3(n_192),
.B1(n_189),
.B2(n_182),
.C(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_184),
.C(n_191),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_223),
.C(n_187),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_215),
.B(n_216),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_186),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_225),
.B1(n_202),
.B2(n_214),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_196),
.B(n_204),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_227),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_198),
.B1(n_202),
.B2(n_211),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_204),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_226),
.B(n_186),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_187),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_232),
.A2(n_221),
.B1(n_225),
.B2(n_227),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_231),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_220),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_231),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_237),
.B(n_234),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_183),
.B(n_169),
.C(n_176),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_242),
.C(n_183),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_151),
.Y(n_247)
);


endmodule