module fake_jpeg_11611_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_30),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_0),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_43),
.B(n_50),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_1),
.B(n_2),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_51),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_46),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_43),
.C(n_36),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_45),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_76),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_79),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_20),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_3),
.B(n_4),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_5),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_7),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_8),
.B(n_9),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_10),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_12),
.C(n_13),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_22),
.CI(n_27),
.CON(n_102),
.SN(n_102)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_15),
.B(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_21),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_111),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_95),
.B(n_91),
.C(n_88),
.D(n_98),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_107),
.C(n_93),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_113),
.B1(n_104),
.B2(n_110),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_108),
.C(n_106),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_105),
.Y(n_119)
);


endmodule