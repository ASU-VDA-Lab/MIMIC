module real_aes_6402_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp5_ASAP7_75t_SL g377 ( .A1(n_0), .A2(n_236), .B1(n_333), .B2(n_378), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_1), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_2), .A2(n_230), .B1(n_527), .B2(n_594), .Y(n_700) );
INVx1_ASAP7_75t_L g287 ( .A(n_3), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_4), .A2(n_112), .B1(n_386), .B2(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_5), .A2(n_16), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_6), .A2(n_62), .B1(n_390), .B2(n_422), .Y(n_653) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_7), .A2(n_17), .B1(n_389), .B2(n_476), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_8), .A2(n_124), .B1(n_637), .B2(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_9), .A2(n_35), .B1(n_504), .B2(n_836), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_10), .A2(n_148), .B1(n_432), .B2(n_526), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_11), .A2(n_121), .B1(n_430), .B2(n_594), .Y(n_752) );
AOI222xp33_ASAP7_75t_L g506 ( .A1(n_12), .A2(n_123), .B1(n_218), .B2(n_386), .C1(n_507), .C2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_13), .A2(n_53), .B1(n_457), .B2(n_468), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_14), .A2(n_59), .B1(n_472), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_15), .A2(n_139), .B1(n_504), .B2(n_670), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_18), .Y(n_383) );
AOI222xp33_ASAP7_75t_L g475 ( .A1(n_19), .A2(n_84), .B1(n_138), .B2(n_407), .C1(n_476), .C2(n_477), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_20), .A2(n_165), .B1(n_434), .B2(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_21), .B(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_22), .A2(n_122), .B1(n_435), .B2(n_704), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_23), .Y(n_368) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_24), .A2(n_87), .B1(n_295), .B2(n_300), .Y(n_303) );
INVx1_ASAP7_75t_L g779 ( .A(n_24), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_25), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_26), .A2(n_197), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_27), .A2(n_268), .B1(n_330), .B2(n_333), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_28), .A2(n_209), .B1(n_365), .B2(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_29), .A2(n_145), .B1(n_597), .B2(n_600), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_30), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_31), .A2(n_269), .B1(n_325), .B2(n_526), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_32), .Y(n_812) );
INVx1_ASAP7_75t_L g615 ( .A(n_33), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_34), .A2(n_249), .B1(n_306), .B2(n_660), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_36), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g712 ( .A1(n_37), .A2(n_194), .B1(n_245), .B2(n_352), .C1(n_508), .C2(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_38), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_39), .B(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_40), .A2(n_187), .B1(n_416), .B2(n_523), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_41), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_42), .A2(n_258), .B1(n_320), .B2(n_599), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_43), .Y(n_423) );
INVx1_ASAP7_75t_L g655 ( .A(n_44), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_45), .A2(n_172), .B1(n_390), .B2(n_523), .Y(n_522) );
AO22x2_ASAP7_75t_L g305 ( .A1(n_46), .A2(n_90), .B1(n_295), .B2(n_296), .Y(n_305) );
INVx1_ASAP7_75t_L g780 ( .A(n_46), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_47), .Y(n_443) );
INVx1_ASAP7_75t_L g578 ( .A(n_48), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_49), .A2(n_144), .B1(n_792), .B2(n_793), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_50), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_51), .A2(n_255), .B1(n_394), .B2(n_519), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_52), .A2(n_161), .B1(n_291), .B2(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_54), .A2(n_208), .B1(n_357), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_55), .A2(n_83), .B1(n_467), .B2(n_468), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_56), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_57), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_58), .Y(n_805) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_60), .A2(n_63), .B1(n_556), .B2(n_557), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_61), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_64), .A2(n_73), .B1(n_330), .B2(n_639), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_65), .Y(n_760) );
AOI22xp5_ASAP7_75t_SL g373 ( .A1(n_66), .A2(n_156), .B1(n_374), .B2(n_375), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_67), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_68), .A2(n_134), .B1(n_635), .B2(n_699), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_69), .A2(n_150), .B1(n_356), .B2(n_389), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_70), .A2(n_193), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_71), .A2(n_198), .B1(n_526), .B2(n_527), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_72), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_74), .A2(n_191), .B1(n_417), .B2(n_710), .Y(n_807) );
AOI22xp5_ASAP7_75t_SL g371 ( .A1(n_75), .A2(n_137), .B1(n_306), .B2(n_372), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_76), .A2(n_224), .B1(n_394), .B2(n_397), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_77), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_78), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g406 ( .A1(n_79), .A2(n_407), .B(n_408), .C(n_419), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_80), .A2(n_107), .B1(n_500), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_81), .A2(n_226), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp5_ASAP7_75t_SL g290 ( .A1(n_82), .A2(n_147), .B1(n_291), .B2(n_306), .Y(n_290) );
INVx1_ASAP7_75t_L g664 ( .A(n_85), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_86), .A2(n_149), .B1(n_325), .B2(n_497), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_88), .A2(n_135), .B1(n_476), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_89), .A2(n_259), .B1(n_374), .B2(n_597), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_91), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_92), .A2(n_203), .B1(n_331), .B2(n_464), .Y(n_730) );
XOR2xp5_ASAP7_75t_L g782 ( .A(n_93), .B(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_94), .Y(n_790) );
AND2x2_ASAP7_75t_L g277 ( .A(n_95), .B(n_278), .Y(n_277) );
AOI22xp5_ASAP7_75t_SL g608 ( .A1(n_96), .A2(n_609), .B1(n_644), .B2(n_645), .Y(n_608) );
INVx1_ASAP7_75t_L g645 ( .A(n_96), .Y(n_645) );
INVx1_ASAP7_75t_L g684 ( .A(n_97), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_98), .A2(n_252), .B1(n_704), .B2(n_706), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_99), .A2(n_132), .B1(n_430), .B2(n_432), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_100), .A2(n_202), .B1(n_490), .B2(n_526), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_101), .Y(n_788) );
AOI22xp5_ASAP7_75t_SL g319 ( .A1(n_102), .A2(n_239), .B1(n_320), .B2(n_325), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_103), .A2(n_183), .B1(n_352), .B2(n_356), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_104), .A2(n_204), .B1(n_430), .B2(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g274 ( .A(n_105), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_106), .A2(n_146), .B1(n_353), .B2(n_365), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_108), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_109), .A2(n_166), .B1(n_493), .B2(n_496), .Y(n_729) );
XOR2x2_ASAP7_75t_L g692 ( .A(n_110), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_111), .B(n_519), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_113), .A2(n_241), .B1(n_499), .B2(n_500), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_114), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g560 ( .A1(n_115), .A2(n_561), .B(n_562), .C(n_568), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_116), .A2(n_219), .B1(n_365), .B2(n_389), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_117), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_118), .A2(n_167), .B1(n_311), .B2(n_317), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_119), .B(n_504), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_120), .A2(n_177), .B1(n_497), .B2(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g674 ( .A(n_125), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_126), .A2(n_234), .B1(n_464), .B2(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_127), .A2(n_240), .B1(n_356), .B2(n_710), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_128), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_129), .A2(n_262), .B1(n_490), .B2(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_130), .A2(n_180), .B1(n_357), .B2(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_131), .A2(n_213), .B1(n_416), .B2(n_417), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_133), .A2(n_261), .B1(n_463), .B2(n_704), .Y(n_753) );
AOI22xp5_ASAP7_75t_SL g736 ( .A1(n_136), .A2(n_737), .B1(n_763), .B2(n_764), .Y(n_736) );
INVx1_ASAP7_75t_L g764 ( .A(n_136), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_140), .A2(n_222), .B1(n_642), .B2(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_141), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_142), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g278 ( .A(n_143), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_151), .Y(n_543) );
INVx1_ASAP7_75t_L g586 ( .A(n_152), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_153), .A2(n_232), .B1(n_357), .B2(n_416), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_154), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_155), .Y(n_740) );
AND2x6_ASAP7_75t_L g273 ( .A(n_157), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_157), .Y(n_773) );
AO22x2_ASAP7_75t_L g294 ( .A1(n_158), .A2(n_231), .B1(n_295), .B2(n_296), .Y(n_294) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_159), .Y(n_404) );
INVx1_ASAP7_75t_L g587 ( .A(n_160), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_162), .A2(n_248), .B1(n_311), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_163), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_164), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_168), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_169), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_170), .A2(n_250), .B1(n_291), .B2(n_490), .Y(n_662) );
OA22x2_ASAP7_75t_L g572 ( .A1(n_171), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_171), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_173), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_174), .A2(n_266), .B1(n_527), .B2(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_175), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_176), .A2(n_184), .B1(n_545), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_178), .A2(n_200), .B1(n_493), .B2(n_556), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_179), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_181), .A2(n_217), .B1(n_633), .B2(n_635), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_182), .A2(n_246), .B1(n_325), .B2(n_497), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_185), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_186), .A2(n_220), .B1(n_352), .B2(n_356), .Y(n_584) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_188), .A2(n_244), .B1(n_295), .B2(n_300), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_189), .A2(n_223), .B1(n_561), .B2(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_190), .A2(n_257), .B1(n_386), .B2(n_523), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_192), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_195), .A2(n_221), .B1(n_591), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g447 ( .A(n_196), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_199), .A2(n_215), .B1(n_461), .B2(n_463), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_201), .A2(n_214), .B1(n_620), .B2(n_831), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_205), .A2(n_264), .B1(n_621), .B2(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g612 ( .A(n_206), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_207), .A2(n_260), .B1(n_306), .B2(n_435), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_210), .B(n_504), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_211), .A2(n_271), .B(n_279), .C(n_781), .Y(n_270) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_212), .A2(n_247), .B1(n_372), .B2(n_375), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_216), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_225), .Y(n_824) );
OA22x2_ASAP7_75t_L g825 ( .A1(n_225), .A2(n_824), .B1(n_826), .B2(n_846), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_227), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_228), .A2(n_237), .B1(n_499), .B2(n_639), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_229), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_231), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_233), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g582 ( .A(n_235), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_238), .Y(n_755) );
INVx1_ASAP7_75t_L g579 ( .A(n_242), .Y(n_579) );
XNOR2xp5_ASAP7_75t_L g539 ( .A(n_243), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g776 ( .A(n_244), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_251), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_253), .A2(n_256), .B1(n_696), .B2(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
OA22x2_ASAP7_75t_L g452 ( .A1(n_263), .A2(n_453), .B1(n_454), .B2(n_478), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_263), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_265), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_267), .Y(n_718) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_274), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_275), .A2(n_771), .B(n_823), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_604), .B1(n_766), .B2(n_767), .C(n_768), .Y(n_279) );
INVx1_ASAP7_75t_L g766 ( .A(n_280), .Y(n_766) );
OAI22xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_282), .B1(n_482), .B2(n_483), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_400), .B1(n_480), .B2(n_481), .Y(n_282) );
INVx1_ASAP7_75t_L g480 ( .A(n_283), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_369), .B2(n_399), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
XNOR2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND3x1_ASAP7_75t_SL g288 ( .A(n_289), .B(n_318), .C(n_335), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_310), .Y(n_289) );
INVx1_ASAP7_75t_L g459 ( .A(n_291), .Y(n_459) );
BUFx2_ASAP7_75t_L g557 ( .A(n_291), .Y(n_557) );
BUFx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g497 ( .A(n_292), .Y(n_497) );
BUFx3_ASAP7_75t_L g592 ( .A(n_292), .Y(n_592) );
BUFx3_ASAP7_75t_L g699 ( .A(n_292), .Y(n_699) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_301), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_293), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_293), .B(n_301), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_293), .B(n_309), .Y(n_564) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
INVx2_ASAP7_75t_L g315 ( .A(n_294), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_294), .B(n_299), .Y(n_328) );
AND2x2_ASAP7_75t_L g344 ( .A(n_294), .B(n_303), .Y(n_344) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_297), .Y(n_300) );
INVx1_ASAP7_75t_L g358 ( .A(n_298), .Y(n_358) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
AND2x2_ASAP7_75t_L g332 ( .A(n_299), .B(n_315), .Y(n_332) );
INVx1_ASAP7_75t_L g355 ( .A(n_299), .Y(n_355) );
AND2x2_ASAP7_75t_L g313 ( .A(n_301), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g326 ( .A(n_301), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g331 ( .A(n_301), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
AND2x2_ASAP7_75t_L g309 ( .A(n_302), .B(n_305), .Y(n_309) );
OR2x2_ASAP7_75t_L g324 ( .A(n_302), .B(n_305), .Y(n_324) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g359 ( .A(n_303), .B(n_305), .Y(n_359) );
INVx1_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
AND2x2_ASAP7_75t_L g367 ( .A(n_304), .B(n_355), .Y(n_367) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g392 ( .A(n_305), .Y(n_392) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g434 ( .A(n_307), .Y(n_434) );
INVx4_ASAP7_75t_L g462 ( .A(n_307), .Y(n_462) );
INVx5_ASAP7_75t_L g493 ( .A(n_307), .Y(n_493) );
INVx2_ASAP7_75t_L g600 ( .A(n_307), .Y(n_600) );
BUFx3_ASAP7_75t_L g638 ( .A(n_307), .Y(n_638) );
INVx8_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g317 ( .A(n_309), .B(n_314), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_309), .B(n_332), .Y(n_339) );
AND2x6_ASAP7_75t_L g397 ( .A(n_309), .B(n_332), .Y(n_397) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx3_ASAP7_75t_L g526 ( .A(n_312), .Y(n_526) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_SL g374 ( .A(n_313), .Y(n_374) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_313), .Y(n_446) );
BUFx2_ASAP7_75t_SL g561 ( .A(n_313), .Y(n_561) );
AND2x6_ASAP7_75t_L g322 ( .A(n_314), .B(n_323), .Y(n_322) );
AND2x6_ASAP7_75t_L g362 ( .A(n_314), .B(n_359), .Y(n_362) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
BUFx3_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
INVx6_ASAP7_75t_L g441 ( .A(n_317), .Y(n_441) );
BUFx3_ASAP7_75t_L g556 ( .A(n_317), .Y(n_556) );
BUFx3_ASAP7_75t_L g599 ( .A(n_317), .Y(n_599) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_329), .Y(n_318) );
INVx1_ASAP7_75t_L g570 ( .A(n_320), .Y(n_570) );
INVx4_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx3_ASAP7_75t_L g372 ( .A(n_321), .Y(n_372) );
INVx2_ASAP7_75t_SL g468 ( .A(n_321), .Y(n_468) );
INVx4_ASAP7_75t_L g696 ( .A(n_321), .Y(n_696) );
INVx11_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx11_ASAP7_75t_L g491 ( .A(n_322), .Y(n_491) );
AND2x4_ASAP7_75t_L g396 ( .A(n_323), .B(n_332), .Y(n_396) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g348 ( .A(n_324), .B(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
BUFx2_ASAP7_75t_L g432 ( .A(n_326), .Y(n_432) );
BUFx3_ASAP7_75t_L g500 ( .A(n_326), .Y(n_500) );
BUFx3_ASAP7_75t_L g594 ( .A(n_326), .Y(n_594) );
BUFx2_ASAP7_75t_SL g635 ( .A(n_326), .Y(n_635) );
BUFx2_ASAP7_75t_SL g800 ( .A(n_326), .Y(n_800) );
AND2x2_ASAP7_75t_L g333 ( .A(n_327), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x6_ASAP7_75t_L g436 ( .A(n_328), .B(n_392), .Y(n_436) );
INVx4_ASAP7_75t_L g431 ( .A(n_330), .Y(n_431) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g380 ( .A(n_331), .Y(n_380) );
BUFx3_ASAP7_75t_L g499 ( .A(n_331), .Y(n_499) );
BUFx3_ASAP7_75t_L g527 ( .A(n_331), .Y(n_527) );
INVx2_ASAP7_75t_L g634 ( .A(n_331), .Y(n_634) );
INVx1_ASAP7_75t_L g349 ( .A(n_332), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_334), .B(n_344), .Y(n_343) );
NOR3xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_346), .C(n_360), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_340), .B1(n_341), .B2(n_345), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g412 ( .A(n_339), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_341), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
INVx3_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_343), .A2(n_421), .B1(n_586), .B2(n_587), .Y(n_585) );
BUFx3_ASAP7_75t_L g624 ( .A(n_343), .Y(n_624) );
AND2x4_ASAP7_75t_L g353 ( .A(n_344), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g366 ( .A(n_344), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g390 ( .A(n_344), .B(n_391), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_350), .B(n_351), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_347), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_577) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g614 ( .A(n_348), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_348), .A2(n_412), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g547 ( .A(n_352), .Y(n_547) );
BUFx4f_ASAP7_75t_L g745 ( .A(n_352), .Y(n_745) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_353), .Y(n_386) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_353), .Y(n_621) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g418 ( .A(n_356), .Y(n_418) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g523 ( .A(n_357), .Y(n_523) );
BUFx2_ASAP7_75t_SL g657 ( .A(n_357), .Y(n_657) );
BUFx2_ASAP7_75t_SL g720 ( .A(n_357), .Y(n_720) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g630 ( .A(n_358), .Y(n_630) );
INVx1_ASAP7_75t_L g629 ( .A(n_359), .Y(n_629) );
OAI22xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_363), .B1(n_364), .B2(n_368), .Y(n_360) );
INVx4_ASAP7_75t_L g713 ( .A(n_361), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_361), .A2(n_743), .B(n_744), .Y(n_742) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
BUFx3_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_362), .Y(n_507) );
INVx2_ASAP7_75t_L g514 ( .A(n_362), .Y(n_514) );
INVx2_ASAP7_75t_SL g811 ( .A(n_362), .Y(n_811) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
BUFx4f_ASAP7_75t_SL g476 ( .A(n_366), .Y(n_476) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_366), .Y(n_508) );
BUFx2_ASAP7_75t_L g831 ( .A(n_366), .Y(n_831) );
INVx2_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
XOR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_398), .Y(n_369) );
NAND4xp75_ASAP7_75t_SL g370 ( .A(n_371), .B(n_373), .C(n_376), .D(n_381), .Y(n_370) );
INVx1_ASAP7_75t_L g439 ( .A(n_372), .Y(n_439) );
INVx1_ASAP7_75t_L g789 ( .A(n_375), .Y(n_789) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_380), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_387), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_385), .Y(n_382) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_384), .A2(n_543), .B1(n_544), .B2(n_546), .C1(n_547), .C2(n_548), .Y(n_542) );
INVx2_ASAP7_75t_L g426 ( .A(n_386), .Y(n_426) );
BUFx4f_ASAP7_75t_SL g477 ( .A(n_386), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_393), .Y(n_387) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVx1_ASAP7_75t_L g711 ( .A(n_390), .Y(n_711) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_394), .Y(n_472) );
INVx5_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g414 ( .A(n_395), .Y(n_414) );
INVx2_ASAP7_75t_L g504 ( .A(n_395), .Y(n_504) );
INVx2_ASAP7_75t_L g521 ( .A(n_395), .Y(n_521) );
INVx4_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g473 ( .A(n_397), .Y(n_473) );
BUFx4f_ASAP7_75t_L g519 ( .A(n_397), .Y(n_519) );
BUFx2_ASAP7_75t_L g670 ( .A(n_397), .Y(n_670) );
INVx1_ASAP7_75t_SL g837 ( .A(n_397), .Y(n_837) );
INVx1_ASAP7_75t_L g481 ( .A(n_400), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_451), .B1(n_452), .B2(n_479), .Y(n_400) );
INVx1_ASAP7_75t_SL g479 ( .A(n_401), .Y(n_479) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_427), .Y(n_405) );
INVx3_ASAP7_75t_L g618 ( .A(n_407), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_413), .C(n_415), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OA211x2_ASAP7_75t_L g501 ( .A1(n_412), .A2(n_502), .B(n_503), .C(n_505), .Y(n_501) );
BUFx3_ASAP7_75t_L g580 ( .A(n_412), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_412), .A2(n_612), .B1(n_613), .B2(n_615), .Y(n_611) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_423), .B2(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_422), .Y(n_545) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_437), .C(n_442), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx6_ASAP7_75t_SL g464 ( .A(n_436), .Y(n_464) );
INVx1_ASAP7_75t_L g602 ( .A(n_436), .Y(n_602) );
INVx1_ASAP7_75t_SL g639 ( .A(n_436), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_437) );
INVx2_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
INVx3_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
INVx2_ASAP7_75t_L g660 ( .A(n_441), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_441), .A2(n_755), .B1(n_756), .B2(n_758), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_442) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g467 ( .A(n_446), .Y(n_467) );
INVx3_ASAP7_75t_L g643 ( .A(n_446), .Y(n_643) );
BUFx3_ASAP7_75t_L g792 ( .A(n_446), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_448), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g478 ( .A(n_454), .Y(n_478) );
NAND4xp75_ASAP7_75t_L g454 ( .A(n_455), .B(n_465), .C(n_470), .D(n_475), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g705 ( .A(n_462), .Y(n_705) );
INVx1_ASAP7_75t_L g566 ( .A(n_463), .Y(n_566) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g529 ( .A(n_464), .Y(n_529) );
BUFx2_ASAP7_75t_L g706 ( .A(n_464), .Y(n_706) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g809 ( .A(n_476), .Y(n_809) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_485), .B1(n_536), .B2(n_537), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_510), .B1(n_534), .B2(n_535), .Y(n_485) );
INVx2_ASAP7_75t_SL g534 ( .A(n_486), .Y(n_534) );
XOR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_509), .Y(n_486) );
NAND4xp75_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .C(n_501), .D(n_506), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
INVx5_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_SL g679 ( .A(n_491), .Y(n_679) );
INVx4_ASAP7_75t_L g757 ( .A(n_491), .Y(n_757) );
INVx1_ASAP7_75t_L g787 ( .A(n_491), .Y(n_787) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
BUFx2_ASAP7_75t_L g844 ( .A(n_499), .Y(n_844) );
INVx2_ASAP7_75t_SL g583 ( .A(n_507), .Y(n_583) );
INVx4_ASAP7_75t_SL g535 ( .A(n_510), .Y(n_535) );
AO22x2_ASAP7_75t_SL g735 ( .A1(n_510), .A2(n_535), .B1(n_736), .B2(n_765), .Y(n_735) );
XOR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_533), .Y(n_510) );
NAND3x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_524), .C(n_530), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_514), .A2(n_655), .B(n_656), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_514), .A2(n_674), .B(n_675), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_514), .A2(n_718), .B(n_719), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g828 ( .A1(n_514), .A2(n_829), .B(n_830), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .C(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g553 ( .A(n_519), .Y(n_553) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
BUFx2_ASAP7_75t_L g797 ( .A(n_527), .Y(n_797) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_SL g537 ( .A1(n_538), .A2(n_571), .B1(n_572), .B2(n_603), .Y(n_537) );
INVx1_ASAP7_75t_L g603 ( .A(n_538), .Y(n_603) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND3x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_554), .C(n_560), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g761 ( .A(n_561), .Y(n_761) );
OAI22xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_562) );
BUFx2_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_588), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .C(n_585), .Y(n_576) );
OAI221xp5_ASAP7_75t_SL g804 ( .A1(n_580), .A2(n_613), .B1(n_805), .B2(n_806), .C(n_807), .Y(n_804) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B(n_584), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_595), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .Y(n_589) );
BUFx4f_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g794 ( .A(n_592), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_601), .Y(n_595) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g767 ( .A(n_604), .Y(n_767) );
XOR2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_687), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OA22x2_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_646), .B1(n_685), .B2(n_686), .Y(n_607) );
INVx1_ASAP7_75t_L g685 ( .A(n_608), .Y(n_685) );
INVx2_ASAP7_75t_SL g644 ( .A(n_609), .Y(n_644) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_610), .B(n_631), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_616), .C(n_622), .Y(n_610) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_619), .Y(n_616) );
BUFx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g813 ( .A(n_621), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_622) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
BUFx2_ASAP7_75t_L g748 ( .A(n_628), .Y(n_748) );
OR2x6_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND4x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .C(n_640), .D(n_641), .Y(n_631) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g686 ( .A(n_646), .Y(n_686) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_665), .Y(n_646) );
XOR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_664), .Y(n_647) );
NAND4xp75_ASAP7_75t_SL g648 ( .A(n_649), .B(n_658), .C(n_662), .D(n_663), .Y(n_648) );
NOR2xp67_ASAP7_75t_SL g649 ( .A(n_650), .B(n_654), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .C(n_653), .Y(n_650) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
XOR2x2_ASAP7_75t_SL g665 ( .A(n_666), .B(n_684), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_667), .B(n_676), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_673), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .C(n_672), .Y(n_668) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_734), .B2(n_735), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AO22x1_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_714), .B1(n_732), .B2(n_733), .Y(n_691) );
INVx1_ASAP7_75t_L g732 ( .A(n_692), .Y(n_732) );
NAND4xp75_ASAP7_75t_L g693 ( .A(n_694), .B(n_701), .C(n_707), .D(n_712), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g834 ( .A(n_711), .Y(n_834) );
INVx3_ASAP7_75t_SL g733 ( .A(n_714), .Y(n_733) );
XOR2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_731), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_716), .B(n_724), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g765 ( .A(n_736), .Y(n_765) );
INVx1_ASAP7_75t_L g763 ( .A(n_737), .Y(n_763) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_750), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .C(n_746), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .C(n_759), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_774), .Y(n_769) );
OR2x2_ASAP7_75t_SL g849 ( .A(n_770), .B(n_775), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_771), .Y(n_816) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_772), .B(n_820), .Y(n_823) );
CKINVDCx16_ASAP7_75t_R g820 ( .A(n_773), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
OAI322xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_815), .A3(n_817), .B1(n_821), .B2(n_824), .C1(n_825), .C2(n_847), .Y(n_781) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_803), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_795), .Y(n_784) );
OAI221xp5_ASAP7_75t_SL g785 ( .A1(n_786), .A2(n_788), .B1(n_789), .B2(n_790), .C(n_791), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI221xp5_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_798), .B1(n_799), .B2(n_801), .C(n_802), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_SL g803 ( .A(n_804), .B(n_808), .Y(n_803) );
OAI222xp33_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_811), .B2(n_812), .C1(n_813), .C2(n_814), .Y(n_808) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g846 ( .A(n_826), .Y(n_846) );
NAND2x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_838), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_832), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
INVx1_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_839), .B(n_842), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
endmodule