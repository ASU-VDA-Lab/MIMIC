module real_jpeg_19414_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_321, n_11, n_14, n_7, n_322, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_321;
input n_11;
input n_14;
input n_7;
input n_322;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_0),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_111),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_0),
.A2(n_58),
.B1(n_59),
.B2(n_111),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_111),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_1),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_107),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_107),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_107),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_3),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_242)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_5),
.B(n_34),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_5),
.A2(n_16),
.B(n_58),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_116),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_5),
.A2(n_95),
.B1(n_96),
.B2(n_174),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_41),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_36),
.B(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_6),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_80),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_80),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_38),
.B1(n_58),
.B2(n_59),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_7),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_277)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_10),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_113),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_113),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_113),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_12),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_118),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_118),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_118),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_13),
.A2(n_30),
.B1(n_58),
.B2(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_13),
.A2(n_30),
.B1(n_43),
.B2(n_44),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_14),
.A2(n_36),
.A3(n_44),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_16),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_16),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

BUFx3_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_86),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_22),
.B(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_27),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_32),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g115 ( 
.A(n_29),
.B(n_116),
.CON(n_115),
.SN(n_115)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_34),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_31),
.A2(n_34),
.B1(n_79),
.B2(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_32),
.B(n_36),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_33),
.A2(n_35),
.B1(n_115),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_42),
.B(n_45),
.C(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_35),
.B(n_116),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_46),
.B(n_49),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_46),
.B1(n_49),
.B2(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_46),
.B1(n_62),
.B2(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_41),
.A2(n_46),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_41),
.A2(n_46),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_42),
.A2(n_47),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_42),
.A2(n_47),
.B1(n_112),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_42),
.A2(n_47),
.B1(n_142),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_42),
.A2(n_47),
.B1(n_126),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_42),
.A2(n_47),
.B1(n_84),
.B2(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_43),
.B(n_45),
.Y(n_200)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_44),
.A2(n_56),
.B(n_116),
.C(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_61),
.C(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_53),
.A2(n_76),
.B1(n_82),
.B2(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_57),
.B(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_57),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_57),
.B1(n_101),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_54),
.A2(n_57),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_54),
.A2(n_57),
.B1(n_169),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_54),
.A2(n_57),
.B1(n_189),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_54),
.A2(n_57),
.B1(n_106),
.B2(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_54),
.A2(n_57),
.B1(n_102),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_54),
.A2(n_57),
.B1(n_244),
.B2(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_54),
.A2(n_57),
.B1(n_60),
.B2(n_277),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_57),
.B(n_116),
.Y(n_172)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_59),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_65),
.A2(n_68),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_65),
.A2(n_68),
.B1(n_124),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_65),
.A2(n_68),
.B1(n_251),
.B2(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.C(n_81),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_71),
.A2(n_72),
.B1(n_77),
.B2(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_77),
.C(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_77),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_77),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_81),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_300),
.A3(n_312),
.B1(n_318),
.B2(n_319),
.C(n_321),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_281),
.B(n_299),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_257),
.B(n_280),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_148),
.B(n_233),
.C(n_256),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_133),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_91),
.B(n_133),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_119),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_93),
.B(n_103),
.C(n_119),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_94),
.B(n_100),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_95),
.A2(n_96),
.B1(n_132),
.B2(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_95),
.A2(n_96),
.B1(n_158),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_95),
.A2(n_161),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_95),
.A2(n_96),
.B1(n_147),
.B2(n_192),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_95),
.A2(n_191),
.B(n_242),
.Y(n_275)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_98),
.B(n_116),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_114),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_128),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_121),
.B(n_127),
.C(n_128),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_131),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_134),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_145),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_140),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_144),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_232),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_227),
.B(n_231),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_213),
.B(n_226),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_194),
.B(n_212),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_181),
.B(n_193),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_170),
.B(n_180),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_162),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_166),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_175),
.B(n_179),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_202),
.B1(n_210),
.B2(n_211),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_197),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_199),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_223),
.C(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_222),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_235),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_255),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_246),
.C(n_255),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_249),
.C(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_279),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_272),
.B2(n_273),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_273),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_265),
.C(n_269),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_271),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_278),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_275),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_275),
.A2(n_292),
.B1(n_295),
.B2(n_322),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_297),
.B2(n_298),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_291),
.C(n_298),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B(n_290),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_302),
.C(n_308),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_302),
.B1(n_303),
.B2(n_317),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_310),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_309),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);


endmodule