module fake_jpeg_3653_n_78 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_20),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_27),
.B(n_26),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_37),
.B1(n_32),
.B2(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_37)
);

NAND2xp67_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_21),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_32),
.B(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_18),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_35),
.B1(n_39),
.B2(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_40),
.B1(n_39),
.B2(n_44),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_42),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_47),
.B(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_59),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_17),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_16),
.C(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_13),
.B1(n_8),
.B2(n_9),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_64)
);

A2O1A1O1Ixp25_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_7),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_47),
.B(n_5),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_4),
.C(n_6),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_69),
.B(n_61),
.Y(n_74)
);

NOR2xp67_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_69),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_73),
.B(n_72),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_64),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_12),
.Y(n_78)
);


endmodule