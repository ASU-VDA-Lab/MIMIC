module fake_jpeg_7302_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_33),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_0),
.CON(n_36),
.SN(n_36)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_18),
.B(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_24),
.B(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_27),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_29),
.B1(n_16),
.B2(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_50),
.B1(n_58),
.B2(n_63),
.Y(n_77)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

OA22x2_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_23),
.B1(n_27),
.B2(n_19),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_39),
.B1(n_40),
.B2(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_29),
.B1(n_40),
.B2(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_29),
.B1(n_21),
.B2(n_22),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_39),
.B1(n_18),
.B2(n_33),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_26),
.B1(n_32),
.B2(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_30),
.B1(n_32),
.B2(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_39),
.B1(n_0),
.B2(n_2),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_38),
.B1(n_28),
.B2(n_22),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_69),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_39),
.B1(n_23),
.B2(n_37),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_90),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_83),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_0),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_14),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_11),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_42),
.Y(n_97)
);

AO21x2_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_60),
.B(n_34),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_97),
.B1(n_78),
.B2(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_115),
.B1(n_78),
.B2(n_94),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_10),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_3),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_79),
.B1(n_88),
.B2(n_3),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_37),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_122),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_37),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_64),
.B(n_1),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_73),
.C(n_84),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_129),
.C(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_128),
.B(n_133),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_75),
.C(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_134),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_76),
.B1(n_80),
.B2(n_83),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_135),
.B1(n_137),
.B2(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_74),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_77),
.B1(n_69),
.B2(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_74),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_77),
.B1(n_85),
.B2(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_143),
.B1(n_145),
.B2(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_144),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_81),
.B1(n_88),
.B2(n_79),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_1),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_2),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_155),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_158),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_142),
.B1(n_126),
.B2(n_115),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_178),
.B1(n_180),
.B2(n_185),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_103),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_111),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_162),
.B(n_179),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_182),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_111),
.B(n_106),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_177),
.B(n_184),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_106),
.C(n_125),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_146),
.C(n_125),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_152),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_111),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_122),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_131),
.B1(n_101),
.B2(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_195),
.B1(n_204),
.B2(n_208),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_209),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_145),
.B1(n_101),
.B2(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_196),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_123),
.B1(n_122),
.B2(n_117),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_117),
.C(n_112),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_173),
.C(n_157),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_159),
.B(n_186),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_105),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_123),
.B1(n_105),
.B2(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_107),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_120),
.B1(n_124),
.B2(n_42),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_216),
.C(n_217),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_175),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_226),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_171),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_225),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_183),
.B1(n_167),
.B2(n_161),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_208),
.B1(n_124),
.B2(n_120),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_178),
.C(n_159),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_197),
.B(n_190),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_168),
.C(n_165),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_232),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_165),
.C(n_120),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_219),
.C(n_223),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_241),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_225),
.CI(n_213),
.CON(n_253),
.SN(n_253)
);

AOI221xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_206),
.B1(n_190),
.B2(n_189),
.C(n_199),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_198),
.B(n_195),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_242),
.A2(n_247),
.B(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_204),
.B1(n_165),
.B2(n_211),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_41),
.B1(n_6),
.B2(n_7),
.Y(n_261)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_249),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_228),
.B1(n_41),
.B2(n_34),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_110),
.B(n_124),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_4),
.C(n_5),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_217),
.B1(n_230),
.B2(n_221),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_248),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_247),
.B1(n_239),
.B2(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_262),
.C(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_243),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_228),
.B1(n_5),
.B2(n_6),
.Y(n_260)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_34),
.C(n_7),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_237),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_273),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_249),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_248),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_253),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_282),
.B(n_262),
.Y(n_285)
);

AOI21x1_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_235),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_279),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_269),
.A2(n_263),
.B(n_256),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_235),
.B(n_256),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_272),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_252),
.C(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_288),
.A3(n_281),
.B1(n_286),
.B2(n_253),
.C1(n_274),
.C2(n_12),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_266),
.C(n_259),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_4),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_14),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_15),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_15),
.C(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_15),
.Y(n_297)
);


endmodule