module fake_netlist_6_660_n_3395 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_951, n_783, n_106, n_725, n_952, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_969, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_360, n_945, n_603, n_119, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_797, n_666, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_589, n_860, n_481, n_788, n_819, n_939, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_561, n_33, n_477, n_549, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_941, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_355, n_426, n_317, n_149, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3395);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_969;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_945;
input n_603;
input n_119;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3395;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_3368;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_1658;
wire n_2593;
wire n_3269;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_1543;
wire n_2811;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_2831;
wire n_2998;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3247;
wire n_3069;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_1214;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3153;
wire n_1188;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_3280;
wire n_1515;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_1369;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_2750;
wire n_1164;
wire n_1627;
wire n_1295;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_2913;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_1952;
wire n_2573;
wire n_2646;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_3179;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_2435;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3306;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_1223;
wire n_2990;
wire n_1775;
wire n_1773;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_2327;
wire n_2201;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_1841;
wire n_2823;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3379;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1650;
wire n_1045;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_988;
wire n_2140;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2787;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_3215;
wire n_3336;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_2649;
wire n_2721;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3290;
wire n_1109;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_3361;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3359;
wire n_2795;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g974 ( 
.A(n_927),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_954),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_5),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_567),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_944),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_186),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_764),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_940),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_621),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_597),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_857),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_379),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_820),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_532),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_546),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_672),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_134),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_515),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_759),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_959),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_873),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_252),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_851),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_926),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_62),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_881),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_665),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_15),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_696),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_815),
.Y(n_1003)
);

CKINVDCx16_ASAP7_75t_R g1004 ( 
.A(n_938),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_832),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_621),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_386),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_966),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_264),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_839),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_769),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_871),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_916),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_260),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_825),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_426),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_461),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_819),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_8),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_378),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_178),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_387),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_785),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_941),
.Y(n_1024)
);

BUFx5_ASAP7_75t_L g1025 ( 
.A(n_674),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_945),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_803),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_6),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_967),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_681),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_291),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_22),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_110),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_863),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_823),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_746),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_969),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_662),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_930),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_166),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_667),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_288),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_446),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_747),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_594),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_874),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_935),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_229),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_149),
.Y(n_1049)
);

CKINVDCx16_ASAP7_75t_R g1050 ( 
.A(n_615),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_176),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_853),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_660),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_565),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_420),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_893),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_295),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_679),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_252),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_730),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_279),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_664),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_846),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_876),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_615),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_858),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_867),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_217),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_48),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_161),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_256),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_913),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_69),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_212),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_933),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_701),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_403),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_650),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_673),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_566),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_160),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_868),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_355),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_63),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_894),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_348),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_880),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_150),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_683),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_680),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_195),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_865),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_60),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_639),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_682),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_664),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_908),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_519),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_883),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_914),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_323),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_889),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_404),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_36),
.Y(n_1104)
);

BUFx2_ASAP7_75t_SL g1105 ( 
.A(n_879),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_387),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_796),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_306),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_182),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_593),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_268),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_310),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_188),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_388),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_878),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_121),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_934),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_862),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_431),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_8),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_512),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_668),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_158),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_905),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_419),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_379),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_627),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_95),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_224),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_953),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_131),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_283),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_482),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_160),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_350),
.Y(n_1135)
);

BUFx5_ASAP7_75t_L g1136 ( 
.A(n_711),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_535),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_833),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_929),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_113),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_33),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_294),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_423),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_904),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_13),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_671),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_168),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_544),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_656),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_675),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_875),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_676),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_275),
.Y(n_1153)
);

CKINVDCx16_ASAP7_75t_R g1154 ( 
.A(n_345),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_921),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_418),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_854),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_968),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_530),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_524),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_299),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_426),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_821),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_760),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_920),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_687),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_537),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_412),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_713),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_566),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_450),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_677),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_468),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_717),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_230),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_612),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_343),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_447),
.Y(n_1178)
);

CKINVDCx16_ASAP7_75t_R g1179 ( 
.A(n_476),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_84),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_956),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_608),
.Y(n_1182)
);

BUFx5_ASAP7_75t_L g1183 ( 
.A(n_903),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_202),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_36),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_970),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_898),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_931),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_315),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_302),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_939),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_762),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_282),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_684),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_277),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_870),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_152),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_923),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_94),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_890),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_864),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_866),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_204),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_132),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_950),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_21),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_757),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_922),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_666),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_902),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_919),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_249),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_932),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_884),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_107),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_530),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_756),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_200),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_461),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_492),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_97),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_678),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_544),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_115),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_725),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_136),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_828),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_885),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_439),
.Y(n_1229)
);

CKINVDCx14_ASAP7_75t_R g1230 ( 
.A(n_872),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_89),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_443),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_877),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_680),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_106),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_901),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_670),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_6),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_386),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_928),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_896),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_91),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_673),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_468),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_744),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_636),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_563),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_392),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_856),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_182),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_869),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_787),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_360),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_84),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_663),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_28),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_342),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_422),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_888),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_784),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_882),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_690),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_362),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_600),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_861),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_841),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_918),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_915),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_46),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_234),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_860),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_951),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_216),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_510),
.Y(n_1274)
);

INVxp33_ASAP7_75t_L g1275 ( 
.A(n_617),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_223),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_336),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_125),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_706),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_753),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_677),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_572),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_834),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_910),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_431),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_466),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_773),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_420),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_689),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_830),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_577),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_855),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_140),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_227),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_337),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_635),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_53),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_435),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_907),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_303),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_315),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_467),
.Y(n_1302)
);

BUFx10_ASAP7_75t_L g1303 ( 
.A(n_912),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_895),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_320),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_642),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_909),
.Y(n_1307)
);

BUFx10_ASAP7_75t_L g1308 ( 
.A(n_624),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_147),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_900),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_110),
.Y(n_1311)
);

BUFx8_ASAP7_75t_SL g1312 ( 
.A(n_335),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_317),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_937),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_448),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_782),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_899),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_92),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_925),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_891),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_11),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_671),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_936),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_887),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_886),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_423),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_652),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_557),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_283),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_906),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_911),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_143),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_122),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_70),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_350),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_702),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_917),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_924),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_23),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_897),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_187),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_697),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_892),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_220),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_146),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_816),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_859),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_304),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_669),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_129),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1050),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1025),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1025),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1025),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1025),
.Y(n_1355)
);

BUFx10_ASAP7_75t_L g1356 ( 
.A(n_1120),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1025),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1312),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_975),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1008),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_979),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_980),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_979),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_979),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1053),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1053),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1053),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_1265),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_984),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1112),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1065),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1065),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1065),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1104),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1104),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1104),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1135),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1135),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1135),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1029),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1141),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_986),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_992),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1272),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1154),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1141),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1141),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1195),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1067),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_996),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1195),
.Y(n_1391)
);

INVxp33_ASAP7_75t_SL g1392 ( 
.A(n_1270),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1195),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1179),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1115),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1226),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1226),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1226),
.Y(n_1398)
);

INVxp33_ASAP7_75t_SL g1399 ( 
.A(n_1006),
.Y(n_1399)
);

CKINVDCx16_ASAP7_75t_R g1400 ( 
.A(n_1315),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1156),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1260),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1234),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1152),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_989),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_978),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1287),
.Y(n_1407)
);

INVxp33_ASAP7_75t_SL g1408 ( 
.A(n_1329),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_990),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1000),
.Y(n_1410)
);

CKINVDCx14_ASAP7_75t_R g1411 ( 
.A(n_1230),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1016),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1020),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1021),
.Y(n_1414)
);

INVxp67_ASAP7_75t_SL g1415 ( 
.A(n_1060),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1272),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1028),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_997),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1031),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1002),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1352),
.A2(n_1063),
.B(n_1012),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1411),
.B(n_1292),
.Y(n_1423)
);

INVx5_ASAP7_75t_L g1424 ( 
.A(n_1384),
.Y(n_1424)
);

XOR2xp5_ASAP7_75t_L g1425 ( 
.A(n_1360),
.B(n_1319),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1380),
.B(n_1082),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1396),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1361),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_L g1429 ( 
.A(n_1359),
.B(n_977),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1362),
.B(n_993),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1384),
.Y(n_1431)
);

AND2x6_ASAP7_75t_L g1432 ( 
.A(n_1353),
.B(n_1272),
.Y(n_1432)
);

AND2x6_ASAP7_75t_L g1433 ( 
.A(n_1354),
.B(n_1279),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1363),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1400),
.B(n_974),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1384),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1369),
.B(n_1024),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1416),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1399),
.A2(n_1200),
.B1(n_1004),
.B2(n_1061),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1364),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1355),
.B(n_1158),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1416),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1382),
.B(n_1037),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1416),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1383),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1365),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1366),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1367),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1390),
.B(n_1202),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1371),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1351),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1401),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1372),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1370),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1373),
.Y(n_1455)
);

CKINVDCx6p67_ASAP7_75t_R g1456 ( 
.A(n_1385),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1374),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1375),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1408),
.A2(n_1275),
.B1(n_1127),
.B2(n_985),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1376),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1392),
.A2(n_1246),
.B1(n_983),
.B2(n_988),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1378),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1379),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1368),
.B(n_1299),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1418),
.B(n_999),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1406),
.B(n_1029),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1394),
.B(n_982),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1389),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1420),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1415),
.B(n_1249),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1452),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1436),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1442),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1451),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1445),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1469),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1468),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1465),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1431),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1456),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1425),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1430),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1454),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1437),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_R g1486 ( 
.A(n_1429),
.B(n_1395),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1443),
.Y(n_1487)
);

BUFx10_ASAP7_75t_L g1488 ( 
.A(n_1426),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1466),
.B(n_1404),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1449),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1444),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1428),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1444),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1439),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1434),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1464),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1440),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1459),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1467),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1441),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1461),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.B(n_1435),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1423),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1427),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1447),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1448),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1447),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1450),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1450),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1463),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1463),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1453),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1458),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1455),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1424),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1457),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1462),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1460),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1422),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1424),
.Y(n_1521)
);

BUFx10_ASAP7_75t_L g1522 ( 
.A(n_1432),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1421),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1432),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1432),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1433),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1433),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1433),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1445),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1445),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1452),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1465),
.B(n_1358),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1445),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1444),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1439),
.A2(n_1407),
.B1(n_1402),
.B2(n_1124),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1436),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1452),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1445),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1445),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1445),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1452),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1468),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1445),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1492),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1491),
.B(n_1405),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1482),
.B(n_1357),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1485),
.B(n_981),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1493),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1499),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1495),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1478),
.B(n_1356),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1475),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1489),
.B(n_1356),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1487),
.B(n_1046),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1504),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1490),
.B(n_994),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1534),
.B(n_1208),
.Y(n_1557)
);

NOR2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1480),
.B(n_1403),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_L g1559 ( 
.A(n_1502),
.B(n_991),
.C(n_987),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1532),
.B(n_1266),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1493),
.Y(n_1561)
);

AND2x6_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1015),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1505),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1508),
.B(n_1330),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1523),
.A2(n_1102),
.B1(n_1205),
.B2(n_1336),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1474),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1497),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1520),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1506),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1507),
.A2(n_1513),
.B1(n_1519),
.B2(n_1494),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1493),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1510),
.B(n_1409),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1500),
.B(n_1023),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1473),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1536),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1472),
.Y(n_1576)
);

AND3x1_ASAP7_75t_L g1577 ( 
.A(n_1535),
.B(n_1222),
.C(n_1001),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1509),
.B(n_1027),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1479),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1511),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1534),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1512),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1515),
.B(n_1052),
.Y(n_1583)
);

BUFx10_ASAP7_75t_L g1584 ( 
.A(n_1476),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1483),
.B(n_1410),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1496),
.B(n_1342),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1529),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1484),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1530),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1517),
.B(n_1518),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1486),
.B(n_1503),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1542),
.Y(n_1592)
);

INVxp33_ASAP7_75t_L g1593 ( 
.A(n_1471),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1521),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1531),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1537),
.Y(n_1596)
);

BUFx8_ASAP7_75t_SL g1597 ( 
.A(n_1477),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1541),
.Y(n_1598)
);

NAND2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1501),
.B(n_976),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1514),
.B(n_1412),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1488),
.B(n_1533),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1498),
.B(n_1080),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1526),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1527),
.B(n_1066),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1488),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1525),
.A2(n_1005),
.B1(n_1010),
.B2(n_1003),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1540),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1522),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1516),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1516),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1522),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1528),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1543),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1481),
.A2(n_1072),
.B1(n_1233),
.B2(n_1165),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1492),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1492),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1492),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1475),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1504),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1491),
.B(n_1413),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1492),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1489),
.B(n_1414),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1492),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1491),
.B(n_1417),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1489),
.B(n_1419),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1504),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1492),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1499),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1492),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1504),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1474),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1542),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1492),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1482),
.B(n_1092),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1482),
.B(n_1097),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1492),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1482),
.B(n_1011),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1491),
.B(n_1381),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1499),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1499),
.B(n_1081),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1505),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1499),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1499),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1504),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1499),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1474),
.Y(n_1647)
);

AND2x6_ASAP7_75t_L g1648 ( 
.A(n_1524),
.B(n_1107),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1532),
.A2(n_1346),
.B(n_1118),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1493),
.Y(n_1650)
);

BUFx10_ASAP7_75t_L g1651 ( 
.A(n_1480),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1492),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1474),
.B(n_1105),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1491),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1504),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1499),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1499),
.Y(n_1657)
);

INVxp33_ASAP7_75t_L g1658 ( 
.A(n_1474),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1478),
.B(n_1093),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1555),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1546),
.B(n_1117),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1547),
.B(n_1013),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1544),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1561),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1659),
.B(n_1055),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1556),
.B(n_1157),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1602),
.B(n_1071),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1635),
.B(n_1636),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1549),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1550),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1560),
.B(n_1164),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1567),
.A2(n_1213),
.B1(n_1214),
.B2(n_1192),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1561),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1629),
.B(n_1018),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1640),
.B(n_1026),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1569),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1578),
.A2(n_1617),
.B(n_1616),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1571),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1618),
.Y(n_1680)
);

INVxp33_ASAP7_75t_L g1681 ( 
.A(n_1641),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1622),
.B(n_1227),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1627),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1624),
.B(n_1228),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1628),
.B(n_1267),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1643),
.B(n_1079),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1630),
.A2(n_1271),
.B1(n_1289),
.B2(n_1268),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1634),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1631),
.Y(n_1689)
);

NAND2xp33_ASAP7_75t_L g1690 ( 
.A(n_1609),
.B(n_1136),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1566),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1644),
.B(n_1034),
.Y(n_1692)
);

BUFx5_ASAP7_75t_L g1693 ( 
.A(n_1637),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1290),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1646),
.B(n_1035),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1656),
.B(n_1036),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1623),
.B(n_1314),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1565),
.A2(n_1261),
.B1(n_1325),
.B2(n_1324),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1551),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1626),
.B(n_1096),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1597),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1582),
.B(n_1039),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1645),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1615),
.A2(n_1338),
.B1(n_1331),
.B2(n_1343),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1583),
.B(n_1044),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1603),
.A2(n_1593),
.B(n_1604),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1658),
.B(n_1108),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1554),
.B(n_1149),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1559),
.A2(n_1064),
.B1(n_1075),
.B2(n_1047),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1655),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1553),
.B(n_1180),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1573),
.B(n_1076),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1571),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1576),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1650),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1632),
.Y(n_1716)
);

INVx5_ASAP7_75t_L g1717 ( 
.A(n_1584),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1568),
.A2(n_1279),
.B(n_1087),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1572),
.B(n_1085),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1575),
.B(n_1099),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1595),
.A2(n_1100),
.B1(n_1138),
.B2(n_1130),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1574),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1570),
.B(n_1139),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1596),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1598),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1585),
.B(n_1144),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1638),
.B(n_1151),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1588),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1649),
.B(n_1155),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1562),
.A2(n_1183),
.B1(n_1136),
.B2(n_1279),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1562),
.B(n_1163),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1647),
.B(n_1098),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1562),
.B(n_1648),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1590),
.B(n_1189),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1579),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1581),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1648),
.B(n_1166),
.Y(n_1737)
);

AND2x6_ASAP7_75t_L g1738 ( 
.A(n_1609),
.B(n_1042),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1610),
.A2(n_1611),
.B(n_1612),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1607),
.A2(n_1599),
.B(n_1580),
.C(n_1564),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1648),
.B(n_1169),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1548),
.Y(n_1742)
);

NOR2xp67_ASAP7_75t_L g1743 ( 
.A(n_1563),
.B(n_1174),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1642),
.B(n_1608),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1613),
.B(n_1181),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1650),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1639),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1545),
.Y(n_1748)
);

OAI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1653),
.A2(n_1349),
.B1(n_1109),
.B2(n_1178),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1653),
.A2(n_1136),
.B1(n_1183),
.B2(n_1056),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1621),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1552),
.B(n_1186),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1625),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1654),
.B(n_1187),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1557),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1586),
.B(n_1591),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1606),
.A2(n_1106),
.B(n_1074),
.C(n_1077),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1605),
.B(n_1600),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1587),
.B(n_995),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1614),
.B(n_1601),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1577),
.B(n_1188),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1558),
.B(n_1191),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1589),
.B(n_998),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1619),
.B(n_1131),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1592),
.A2(n_1198),
.B1(n_1201),
.B2(n_1196),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1633),
.A2(n_1210),
.B(n_1207),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1594),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1651),
.A2(n_1084),
.B(n_1090),
.C(n_1051),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1549),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1546),
.B(n_1211),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_SL g1771 ( 
.A(n_1552),
.B(n_1056),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1546),
.B(n_1217),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_SL g1773 ( 
.A(n_1584),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1544),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1546),
.B(n_1225),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1546),
.B(n_1236),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1546),
.B(n_1240),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1546),
.B(n_1241),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1546),
.B(n_1245),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1546),
.B(n_1251),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1546),
.A2(n_1259),
.B(n_1252),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1555),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1659),
.B(n_1007),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1546),
.B(n_1262),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1659),
.B(n_1131),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1546),
.B(n_1280),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1546),
.B(n_1283),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1544),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1555),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1555),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1629),
.B(n_1386),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1597),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1546),
.B(n_1284),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1546),
.B(n_1304),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1546),
.B(n_1307),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1555),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1560),
.A2(n_1183),
.B1(n_1136),
.B2(n_1303),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1555),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1546),
.B(n_1310),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1659),
.B(n_1308),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1546),
.B(n_1316),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1659),
.B(n_1009),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1546),
.B(n_1320),
.Y(n_1803)
);

NAND2xp33_ASAP7_75t_L g1804 ( 
.A(n_1609),
.B(n_1136),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1549),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1560),
.A2(n_1323),
.B1(n_1340),
.B2(n_1337),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1546),
.B(n_1347),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1546),
.B(n_1183),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1560),
.A2(n_1017),
.B1(n_1019),
.B2(n_1014),
.Y(n_1809)
);

OAI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1615),
.A2(n_1111),
.B1(n_1114),
.B2(n_1103),
.C(n_1101),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1544),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1546),
.B(n_1303),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1546),
.B(n_1317),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1544),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1546),
.B(n_1317),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1555),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1546),
.B(n_1183),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1544),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1544),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1669),
.A2(n_1388),
.B(n_1387),
.Y(n_1820)
);

AOI33xp33_ASAP7_75t_L g1821 ( 
.A1(n_1700),
.A2(n_1132),
.A3(n_1133),
.B1(n_1146),
.B2(n_1145),
.B3(n_1123),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1678),
.A2(n_1393),
.B(n_1391),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1672),
.A2(n_1160),
.B(n_1147),
.Y(n_1823)
);

INVx5_ASAP7_75t_L g1824 ( 
.A(n_1665),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1783),
.B(n_1022),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1751),
.B(n_1162),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1665),
.Y(n_1827)
);

INVx4_ASAP7_75t_L g1828 ( 
.A(n_1717),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1668),
.B(n_1030),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1808),
.A2(n_1168),
.B(n_1167),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1666),
.A2(n_1033),
.B1(n_1038),
.B2(n_1032),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1756),
.B(n_1040),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1802),
.B(n_1041),
.Y(n_1833)
);

AOI222xp33_ASAP7_75t_L g1834 ( 
.A1(n_1708),
.A2(n_1308),
.B1(n_1322),
.B2(n_1339),
.C1(n_1294),
.C2(n_1258),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1772),
.B(n_1043),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1706),
.A2(n_1398),
.B(n_1397),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1785),
.B(n_1045),
.Y(n_1837)
);

BUFx12f_ASAP7_75t_L g1838 ( 
.A(n_1691),
.Y(n_1838)
);

NOR2xp67_ASAP7_75t_L g1839 ( 
.A(n_1717),
.B(n_685),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1775),
.B(n_1048),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1777),
.B(n_1049),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1697),
.A2(n_1172),
.B(n_1171),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1664),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1739),
.A2(n_1185),
.B(n_1173),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1817),
.A2(n_1209),
.B(n_1190),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1778),
.B(n_1057),
.Y(n_1846)
);

NOR3xp33_ASAP7_75t_L g1847 ( 
.A(n_1711),
.B(n_1686),
.C(n_1758),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1780),
.B(n_1058),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1716),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1660),
.Y(n_1850)
);

AO21x2_ASAP7_75t_L g1851 ( 
.A1(n_1729),
.A2(n_1661),
.B(n_1667),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1784),
.B(n_1059),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1699),
.B(n_1062),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1793),
.A2(n_1220),
.B(n_1215),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1670),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1799),
.A2(n_1231),
.B(n_1229),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1693),
.B(n_1068),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1671),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1681),
.B(n_1069),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1801),
.A2(n_1242),
.B(n_1238),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1705),
.A2(n_1264),
.B(n_1263),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1663),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1712),
.A2(n_1277),
.B(n_1274),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1677),
.A2(n_1070),
.B1(n_1078),
.B2(n_1073),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1679),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1800),
.B(n_1083),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1683),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1745),
.A2(n_1295),
.B(n_1281),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1680),
.B(n_1086),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1701),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1754),
.A2(n_1776),
.B(n_1770),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1688),
.A2(n_1091),
.B1(n_1094),
.B2(n_1089),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1740),
.A2(n_1302),
.B(n_1306),
.C(n_1298),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1689),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1693),
.B(n_1095),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1753),
.B(n_1311),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1734),
.A2(n_1774),
.B(n_1811),
.C(n_1788),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1814),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1818),
.A2(n_1321),
.B(n_1318),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1819),
.B(n_1110),
.Y(n_1880)
);

OAI321xp33_ASAP7_75t_L g1881 ( 
.A1(n_1749),
.A2(n_1698),
.A3(n_1809),
.B1(n_1797),
.B2(n_1810),
.C(n_1750),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1682),
.A2(n_1348),
.B(n_1328),
.Y(n_1882)
);

A2O1A1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1723),
.A2(n_1088),
.B(n_1170),
.C(n_1054),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1714),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1779),
.A2(n_1224),
.B(n_1204),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1693),
.B(n_1113),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1703),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1786),
.A2(n_1807),
.B(n_1794),
.Y(n_1888)
);

INVx3_ASAP7_75t_SL g1889 ( 
.A(n_1792),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1710),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1693),
.B(n_1116),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1679),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1732),
.B(n_1119),
.Y(n_1893)
);

NAND2x1_ASAP7_75t_L g1894 ( 
.A(n_1782),
.B(n_1250),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1787),
.A2(n_1269),
.B(n_688),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1757),
.A2(n_1122),
.B(n_1125),
.C(n_1121),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1795),
.A2(n_691),
.B(n_686),
.Y(n_1897)
);

CKINVDCx6p67_ASAP7_75t_R g1898 ( 
.A(n_1773),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1728),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1769),
.Y(n_1900)
);

OAI21xp33_ASAP7_75t_L g1901 ( 
.A1(n_1771),
.A2(n_1128),
.B(n_1126),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1719),
.B(n_1129),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1713),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1713),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1760),
.B(n_1805),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1684),
.A2(n_1137),
.B(n_1134),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1726),
.B(n_1140),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1803),
.A2(n_693),
.B(n_692),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1789),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1724),
.B(n_1142),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1725),
.B(n_1143),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1722),
.B(n_1148),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1790),
.B(n_1150),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1727),
.A2(n_1720),
.B(n_1662),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1796),
.A2(n_695),
.B(n_694),
.Y(n_1915)
);

O2A1O1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1812),
.A2(n_1159),
.B(n_1161),
.C(n_1153),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1798),
.A2(n_699),
.B(n_698),
.Y(n_1917)
);

AOI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1685),
.A2(n_703),
.B(n_700),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1816),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1735),
.B(n_1175),
.Y(n_1920)
);

BUFx8_ASAP7_75t_L g1921 ( 
.A(n_1767),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1694),
.A2(n_705),
.B(n_704),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1736),
.Y(n_1923)
);

BUFx4f_ASAP7_75t_L g1924 ( 
.A(n_1746),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1702),
.A2(n_708),
.B(n_707),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1733),
.A2(n_1737),
.B(n_1731),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1741),
.A2(n_710),
.B(n_709),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1742),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_L g1929 ( 
.A(n_1755),
.B(n_712),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1746),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1715),
.A2(n_715),
.B(n_714),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1759),
.B(n_1176),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1674),
.Y(n_1933)
);

AND2x2_ASAP7_75t_SL g1934 ( 
.A(n_1763),
.B(n_0),
.Y(n_1934)
);

AO21x1_ASAP7_75t_L g1935 ( 
.A1(n_1813),
.A2(n_1815),
.B(n_1761),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1738),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1781),
.B(n_1177),
.Y(n_1937)
);

AOI21x1_ASAP7_75t_SL g1938 ( 
.A1(n_1825),
.A2(n_1932),
.B(n_1840),
.Y(n_1938)
);

OR2x6_ASAP7_75t_L g1939 ( 
.A(n_1838),
.B(n_1744),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1833),
.B(n_1707),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1924),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1914),
.A2(n_1926),
.B(n_1871),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1849),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1847),
.B(n_1764),
.Y(n_1944)
);

BUFx12f_ASAP7_75t_L g1945 ( 
.A(n_1828),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1824),
.Y(n_1946)
);

INVxp67_ASAP7_75t_SL g1947 ( 
.A(n_1855),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1893),
.B(n_1791),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1888),
.A2(n_1804),
.B(n_1690),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1837),
.B(n_1748),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1829),
.B(n_1752),
.Y(n_1951)
);

NOR2x1_ASAP7_75t_L g1952 ( 
.A(n_1865),
.B(n_1743),
.Y(n_1952)
);

BUFx12f_ASAP7_75t_L g1953 ( 
.A(n_1921),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1900),
.B(n_1675),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1934),
.B(n_1765),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1905),
.B(n_1762),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1870),
.B(n_1747),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1843),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1858),
.Y(n_1959)
);

O2A1O1Ixp5_ASAP7_75t_L g1960 ( 
.A1(n_1935),
.A2(n_1766),
.B(n_1676),
.C(n_1695),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1892),
.Y(n_1961)
);

BUFx12f_ASAP7_75t_L g1962 ( 
.A(n_1936),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1827),
.Y(n_1963)
);

AOI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1857),
.A2(n_1886),
.B(n_1875),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1877),
.A2(n_1806),
.B1(n_1704),
.B2(n_1721),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1878),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1853),
.B(n_1692),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1851),
.A2(n_1718),
.B(n_1730),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1930),
.Y(n_1969)
);

NOR3xp33_ASAP7_75t_SL g1970 ( 
.A(n_1901),
.B(n_1768),
.C(n_1696),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1831),
.A2(n_1687),
.B(n_1673),
.C(n_1709),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1884),
.A2(n_1899),
.B1(n_1841),
.B2(n_1846),
.Y(n_1972)
);

NOR3xp33_ASAP7_75t_SL g1973 ( 
.A(n_1832),
.B(n_1184),
.C(n_1182),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1919),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1824),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1866),
.B(n_1859),
.Y(n_1976)
);

O2A1O1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1873),
.A2(n_1738),
.B(n_1194),
.C(n_1197),
.Y(n_1977)
);

AOI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1834),
.A2(n_1738),
.B1(n_1199),
.B2(n_1203),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1824),
.B(n_716),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1835),
.B(n_1193),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1827),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1848),
.B(n_1206),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1903),
.B(n_718),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1850),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1852),
.A2(n_1891),
.B(n_1830),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1907),
.B(n_1902),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1904),
.Y(n_1987)
);

AO22x1_ASAP7_75t_L g1988 ( 
.A1(n_1879),
.A2(n_1216),
.B1(n_1218),
.B2(n_1212),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1933),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1862),
.A2(n_1221),
.B1(n_1223),
.B2(n_1219),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1867),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1869),
.B(n_1232),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1874),
.Y(n_1993)
);

O2A1O1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1823),
.A2(n_1237),
.B(n_1239),
.C(n_1235),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1911),
.B(n_1243),
.Y(n_1995)
);

INVx4_ASAP7_75t_L g1996 ( 
.A(n_1904),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1889),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1895),
.A2(n_720),
.B(n_719),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1887),
.Y(n_1999)
);

A2O1A1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1881),
.A2(n_1247),
.B(n_1253),
.C(n_1248),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1890),
.A2(n_1254),
.B1(n_1255),
.B2(n_1244),
.Y(n_2001)
);

A2O1A1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1896),
.A2(n_1257),
.B(n_1276),
.C(n_1273),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1826),
.B(n_1256),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1898),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1882),
.A2(n_1282),
.B1(n_1285),
.B2(n_1278),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1923),
.B(n_1286),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1906),
.A2(n_1876),
.B1(n_1909),
.B2(n_1880),
.Y(n_2007)
);

NOR3xp33_ASAP7_75t_SL g2008 ( 
.A(n_1883),
.B(n_1291),
.C(n_1288),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1821),
.B(n_1293),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1928),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1910),
.B(n_1296),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1937),
.A2(n_722),
.B(n_721),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1912),
.A2(n_1300),
.B1(n_1301),
.B2(n_1297),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1920),
.B(n_1305),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1927),
.A2(n_724),
.B(n_723),
.Y(n_2015)
);

AOI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1897),
.A2(n_1908),
.B(n_1915),
.Y(n_2016)
);

AND3x1_ASAP7_75t_SL g2017 ( 
.A(n_1864),
.B(n_1313),
.C(n_1309),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1913),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1929),
.A2(n_1327),
.B1(n_1332),
.B2(n_1326),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1872),
.B(n_1333),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1854),
.B(n_1334),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1856),
.B(n_1335),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1917),
.A2(n_727),
.B(n_726),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1860),
.B(n_1341),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1868),
.B(n_1344),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1925),
.A2(n_729),
.B(n_728),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1922),
.A2(n_732),
.B(n_731),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1894),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1931),
.A2(n_734),
.B(n_733),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1836),
.A2(n_736),
.B(n_735),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1916),
.B(n_1345),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1918),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1842),
.B(n_1350),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1863),
.A2(n_738),
.B(n_737),
.Y(n_2034)
);

AOI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1861),
.A2(n_740),
.B(n_739),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1844),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1822),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1820),
.Y(n_2038)
);

BUFx12f_ASAP7_75t_L g2039 ( 
.A(n_1839),
.Y(n_2039)
);

AOI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1845),
.A2(n_742),
.B(n_741),
.Y(n_2040)
);

A2O1A1Ixp33_ASAP7_75t_L g2041 ( 
.A1(n_1885),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1833),
.B(n_1),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1833),
.B(n_2),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_SL g2044 ( 
.A(n_1833),
.B(n_3),
.C(n_4),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_1833),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2045)
);

NOR3xp33_ASAP7_75t_L g2046 ( 
.A(n_1833),
.B(n_7),
.C(n_9),
.Y(n_2046)
);

OAI21x1_ASAP7_75t_L g2047 ( 
.A1(n_1926),
.A2(n_745),
.B(n_743),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1847),
.B(n_7),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1833),
.B(n_9),
.Y(n_2049)
);

AND2x6_ASAP7_75t_L g2050 ( 
.A(n_1843),
.B(n_748),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1914),
.A2(n_750),
.B(n_749),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1833),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1833),
.B(n_10),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1924),
.Y(n_2054)
);

OAI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1833),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1914),
.A2(n_752),
.B(n_751),
.Y(n_2056)
);

NOR2xp67_ASAP7_75t_L g2057 ( 
.A(n_1855),
.B(n_754),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1843),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1847),
.B(n_14),
.Y(n_2059)
);

OAI22x1_ASAP7_75t_L g2060 ( 
.A1(n_1833),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1914),
.A2(n_758),
.B(n_755),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1833),
.B(n_15),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1838),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1847),
.B(n_16),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1833),
.B(n_17),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1914),
.A2(n_763),
.B(n_761),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1833),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1942),
.A2(n_958),
.B(n_957),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1940),
.B(n_765),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1958),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_2047),
.A2(n_767),
.B(n_766),
.Y(n_2071)
);

OAI21x1_ASAP7_75t_L g2072 ( 
.A1(n_2016),
.A2(n_770),
.B(n_768),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1943),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_1961),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1959),
.Y(n_2075)
);

OR2x6_ASAP7_75t_L g2076 ( 
.A(n_2054),
.B(n_771),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1948),
.B(n_19),
.Y(n_2077)
);

OAI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_1967),
.A2(n_20),
.B(n_21),
.Y(n_2078)
);

INVx6_ASAP7_75t_L g2079 ( 
.A(n_1996),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1976),
.B(n_22),
.Y(n_2080)
);

OAI21x1_ASAP7_75t_L g2081 ( 
.A1(n_1968),
.A2(n_774),
.B(n_772),
.Y(n_2081)
);

AOI221x1_ASAP7_75t_L g2082 ( 
.A1(n_2046),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.C(n_26),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1941),
.B(n_775),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1997),
.B(n_776),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1950),
.B(n_24),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_1985),
.A2(n_25),
.B(n_26),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2018),
.B(n_27),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1951),
.B(n_27),
.Y(n_2088)
);

OAI21x1_ASAP7_75t_L g2089 ( 
.A1(n_2051),
.A2(n_778),
.B(n_777),
.Y(n_2089)
);

AO31x2_ASAP7_75t_L g2090 ( 
.A1(n_1949),
.A2(n_780),
.A3(n_781),
.B(n_779),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1982),
.B(n_28),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_1963),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1986),
.B(n_29),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_SL g2094 ( 
.A(n_2039),
.B(n_783),
.Y(n_2094)
);

AOI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_1965),
.A2(n_972),
.B(n_971),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1966),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1947),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_2036),
.A2(n_973),
.B(n_788),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_1954),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1972),
.A2(n_949),
.B(n_948),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1957),
.B(n_786),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2058),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_2056),
.A2(n_2066),
.B(n_2061),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2010),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_1955),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1974),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2014),
.B(n_30),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_2037),
.A2(n_790),
.B(n_789),
.Y(n_2108)
);

AOI211x1_ASAP7_75t_L g2109 ( 
.A1(n_2055),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_2042),
.B(n_32),
.Y(n_2110)
);

AO21x2_ASAP7_75t_L g2111 ( 
.A1(n_1964),
.A2(n_792),
.B(n_791),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2044),
.B(n_34),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_2015),
.A2(n_964),
.B(n_963),
.Y(n_2113)
);

OAI21x1_ASAP7_75t_L g2114 ( 
.A1(n_2040),
.A2(n_794),
.B(n_793),
.Y(n_2114)
);

NOR2xp67_ASAP7_75t_L g2115 ( 
.A(n_1989),
.B(n_795),
.Y(n_2115)
);

O2A1O1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_2043),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2049),
.B(n_35),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2053),
.B(n_37),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2062),
.B(n_38),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1984),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_2023),
.A2(n_955),
.B(n_952),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_1969),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2024),
.B(n_38),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1991),
.Y(n_2124)
);

OAI21x1_ASAP7_75t_L g2125 ( 
.A1(n_1938),
.A2(n_798),
.B(n_797),
.Y(n_2125)
);

O2A1O1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_2065),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_1981),
.Y(n_2127)
);

AOI21x1_ASAP7_75t_SL g2128 ( 
.A1(n_2009),
.A2(n_39),
.B(n_40),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2029),
.A2(n_961),
.B(n_960),
.Y(n_2129)
);

AOI21xp5_ASAP7_75t_L g2130 ( 
.A1(n_2038),
.A2(n_965),
.B(n_962),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1944),
.B(n_2007),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1960),
.A2(n_800),
.B(n_799),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_2027),
.A2(n_802),
.B(n_801),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_1956),
.A2(n_2026),
.B(n_1998),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1981),
.Y(n_2135)
);

AO21x2_ASAP7_75t_L g2136 ( 
.A1(n_2002),
.A2(n_2030),
.B(n_2012),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1980),
.B(n_41),
.Y(n_2137)
);

AOI21x1_ASAP7_75t_L g2138 ( 
.A1(n_2028),
.A2(n_2059),
.B(n_2048),
.Y(n_2138)
);

A2O1A1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_2031),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2139)
);

AOI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_1971),
.A2(n_943),
.B(n_942),
.Y(n_2140)
);

NAND3xp33_ASAP7_75t_SL g2141 ( 
.A(n_1994),
.B(n_42),
.C(n_43),
.Y(n_2141)
);

AOI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_1977),
.A2(n_947),
.B(n_946),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1953),
.Y(n_2143)
);

OAI21x1_ASAP7_75t_L g2144 ( 
.A1(n_2034),
.A2(n_805),
.B(n_804),
.Y(n_2144)
);

INVx5_ASAP7_75t_L g2145 ( 
.A(n_1945),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_1992),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_2146)
);

AO31x2_ASAP7_75t_L g2147 ( 
.A1(n_2041),
.A2(n_807),
.A3(n_808),
.B(n_806),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_SL g2148 ( 
.A(n_2004),
.Y(n_2148)
);

NOR4xp25_ASAP7_75t_L g2149 ( 
.A(n_2064),
.B(n_54),
.C(n_62),
.D(n_45),
.Y(n_2149)
);

BUFx8_ASAP7_75t_SL g2150 ( 
.A(n_2004),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2070),
.Y(n_2151)
);

NOR2x1_ASAP7_75t_SL g2152 ( 
.A(n_2111),
.B(n_2032),
.Y(n_2152)
);

O2A1O1Ixp33_ASAP7_75t_SL g2153 ( 
.A1(n_2139),
.A2(n_2067),
.B(n_2000),
.C(n_2022),
.Y(n_2153)
);

NAND2x1p5_ASAP7_75t_L g2154 ( 
.A(n_2097),
.B(n_1946),
.Y(n_2154)
);

AO21x2_ASAP7_75t_L g2155 ( 
.A1(n_2086),
.A2(n_2132),
.B(n_2134),
.Y(n_2155)
);

OAI21x1_ASAP7_75t_L g2156 ( 
.A1(n_2103),
.A2(n_2035),
.B(n_1993),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2080),
.B(n_2060),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2075),
.Y(n_2158)
);

OAI21x1_ASAP7_75t_L g2159 ( 
.A1(n_2072),
.A2(n_1952),
.B(n_1999),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2102),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2074),
.B(n_1957),
.Y(n_2161)
);

INVx1_ASAP7_75t_SL g2162 ( 
.A(n_2099),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_SL g2163 ( 
.A1(n_2078),
.A2(n_2050),
.B1(n_1995),
.B2(n_2020),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_2081),
.A2(n_2021),
.B(n_2032),
.Y(n_2164)
);

OAI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2091),
.A2(n_2107),
.B1(n_2088),
.B2(n_2082),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2095),
.A2(n_2011),
.B(n_2057),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2123),
.B(n_1973),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2106),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_2141),
.A2(n_2045),
.B1(n_2052),
.B2(n_2025),
.Y(n_2169)
);

OA21x2_ASAP7_75t_L g2170 ( 
.A1(n_2125),
.A2(n_2008),
.B(n_1970),
.Y(n_2170)
);

NOR2xp67_ASAP7_75t_L g2171 ( 
.A(n_2145),
.B(n_1962),
.Y(n_2171)
);

OAI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_2140),
.A2(n_2100),
.B(n_2069),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_2092),
.B(n_2063),
.Y(n_2173)
);

AO31x2_ASAP7_75t_L g2174 ( 
.A1(n_2068),
.A2(n_2019),
.A3(n_2013),
.B(n_2006),
.Y(n_2174)
);

OAI21x1_ASAP7_75t_L g2175 ( 
.A1(n_2114),
.A2(n_2071),
.B(n_2089),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_L g2176 ( 
.A1(n_2108),
.A2(n_2033),
.B(n_2001),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_2144),
.A2(n_1990),
.B(n_1975),
.Y(n_2177)
);

INVx4_ASAP7_75t_L g2178 ( 
.A(n_2135),
.Y(n_2178)
);

BUFx2_ASAP7_75t_L g2179 ( 
.A(n_2073),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_2079),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2120),
.Y(n_2181)
);

OAI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_2093),
.A2(n_1978),
.B1(n_1939),
.B2(n_1988),
.Y(n_2182)
);

AND2x4_ASAP7_75t_L g2183 ( 
.A(n_2101),
.B(n_1979),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2142),
.A2(n_2005),
.B(n_2003),
.Y(n_2184)
);

NOR2x1_ASAP7_75t_R g2185 ( 
.A(n_2143),
.B(n_1983),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_2122),
.Y(n_2186)
);

OAI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2137),
.A2(n_1939),
.B1(n_1987),
.B2(n_2017),
.C(n_2050),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2096),
.Y(n_2188)
);

OAI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2131),
.A2(n_2050),
.B(n_47),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_2133),
.A2(n_810),
.B(n_809),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2124),
.Y(n_2191)
);

AO31x2_ASAP7_75t_L g2192 ( 
.A1(n_2121),
.A2(n_2129),
.A3(n_2113),
.B(n_2130),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2117),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2193)
);

INVx5_ASAP7_75t_L g2194 ( 
.A(n_2150),
.Y(n_2194)
);

BUFx6f_ASAP7_75t_L g2195 ( 
.A(n_2135),
.Y(n_2195)
);

O2A1O1Ixp33_ASAP7_75t_SL g2196 ( 
.A1(n_2110),
.A2(n_51),
.B(n_52),
.C(n_50),
.Y(n_2196)
);

AO21x2_ASAP7_75t_L g2197 ( 
.A1(n_2136),
.A2(n_49),
.B(n_50),
.Y(n_2197)
);

OAI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_2138),
.A2(n_51),
.B(n_52),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_2195),
.Y(n_2199)
);

OA21x2_ASAP7_75t_L g2200 ( 
.A1(n_2198),
.A2(n_2119),
.B(n_2118),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_2195),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2186),
.B(n_2104),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_L g2203 ( 
.A1(n_2175),
.A2(n_2128),
.B(n_2098),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2179),
.B(n_2112),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2160),
.Y(n_2205)
);

CKINVDCx6p67_ASAP7_75t_R g2206 ( 
.A(n_2194),
.Y(n_2206)
);

AO31x2_ASAP7_75t_L g2207 ( 
.A1(n_2152),
.A2(n_2105),
.A3(n_2146),
.B(n_2094),
.Y(n_2207)
);

AO31x2_ASAP7_75t_L g2208 ( 
.A1(n_2166),
.A2(n_2077),
.A3(n_2109),
.B(n_2149),
.Y(n_2208)
);

AOI222xp33_ASAP7_75t_L g2209 ( 
.A1(n_2169),
.A2(n_2087),
.B1(n_2085),
.B2(n_2084),
.C1(n_2083),
.C2(n_2148),
.Y(n_2209)
);

AO21x2_ASAP7_75t_L g2210 ( 
.A1(n_2172),
.A2(n_2126),
.B(n_2116),
.Y(n_2210)
);

OA21x2_ASAP7_75t_L g2211 ( 
.A1(n_2159),
.A2(n_2115),
.B(n_2090),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2168),
.Y(n_2212)
);

AOI21x1_ASAP7_75t_L g2213 ( 
.A1(n_2189),
.A2(n_2170),
.B(n_2177),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_2194),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2155),
.A2(n_2076),
.B(n_2147),
.Y(n_2215)
);

OAI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2163),
.A2(n_2076),
.B1(n_2145),
.B2(n_2079),
.Y(n_2216)
);

BUFx2_ASAP7_75t_L g2217 ( 
.A(n_2154),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2181),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2157),
.B(n_2147),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2153),
.A2(n_2090),
.B(n_2127),
.Y(n_2220)
);

AOI21x1_ASAP7_75t_L g2221 ( 
.A1(n_2184),
.A2(n_53),
.B(n_54),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2158),
.Y(n_2222)
);

A2O1A1Ixp33_ASAP7_75t_L g2223 ( 
.A1(n_2187),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2188),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2191),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2151),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_L g2227 ( 
.A1(n_2156),
.A2(n_812),
.B(n_811),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_2162),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_2167),
.B(n_55),
.Y(n_2229)
);

AOI21x1_ASAP7_75t_L g2230 ( 
.A1(n_2190),
.A2(n_56),
.B(n_57),
.Y(n_2230)
);

AOI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_2197),
.A2(n_814),
.B(n_813),
.Y(n_2231)
);

NOR2x1_ASAP7_75t_SL g2232 ( 
.A(n_2180),
.B(n_817),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2164),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_2176),
.A2(n_822),
.B(n_818),
.Y(n_2234)
);

OAI21x1_ASAP7_75t_L g2235 ( 
.A1(n_2192),
.A2(n_826),
.B(n_824),
.Y(n_2235)
);

INVx2_ASAP7_75t_SL g2236 ( 
.A(n_2173),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2161),
.B(n_58),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2185),
.B(n_58),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2178),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2165),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2240)
);

OAI21x1_ASAP7_75t_SL g2241 ( 
.A1(n_2193),
.A2(n_59),
.B(n_61),
.Y(n_2241)
);

AO31x2_ASAP7_75t_L g2242 ( 
.A1(n_2192),
.A2(n_65),
.A3(n_63),
.B(n_64),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2196),
.Y(n_2243)
);

AOI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2182),
.A2(n_829),
.B(n_827),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2174),
.Y(n_2245)
);

NAND2x1p5_ASAP7_75t_L g2246 ( 
.A(n_2171),
.B(n_831),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2183),
.B(n_835),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2174),
.A2(n_837),
.B(n_836),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2160),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2225),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2205),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2204),
.B(n_64),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2212),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2228),
.B(n_65),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2218),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2249),
.Y(n_2256)
);

AO21x2_ASAP7_75t_L g2257 ( 
.A1(n_2245),
.A2(n_66),
.B(n_67),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2222),
.Y(n_2258)
);

OAI21x1_ASAP7_75t_L g2259 ( 
.A1(n_2203),
.A2(n_840),
.B(n_838),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2224),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2202),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2226),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2201),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2242),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2242),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2233),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2217),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2219),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2200),
.B(n_66),
.Y(n_2269)
);

AO21x2_ASAP7_75t_L g2270 ( 
.A1(n_2215),
.A2(n_67),
.B(n_68),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2236),
.B(n_68),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2221),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2210),
.B(n_69),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2213),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2208),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2206),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2208),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2230),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2239),
.B(n_842),
.Y(n_2279)
);

INVx3_ASAP7_75t_L g2280 ( 
.A(n_2199),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2237),
.B(n_70),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_2214),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2243),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2211),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2234),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2220),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2235),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2227),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2229),
.B(n_71),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2207),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2207),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_2246),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2232),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_2238),
.Y(n_2294)
);

OAI21x1_ASAP7_75t_L g2295 ( 
.A1(n_2248),
.A2(n_844),
.B(n_843),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2216),
.Y(n_2296)
);

OAI21x1_ASAP7_75t_L g2297 ( 
.A1(n_2231),
.A2(n_847),
.B(n_845),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2247),
.B(n_71),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2241),
.Y(n_2299)
);

AOI21x1_ASAP7_75t_L g2300 ( 
.A1(n_2244),
.A2(n_72),
.B(n_73),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2209),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2240),
.B(n_72),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2223),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2228),
.B(n_73),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2205),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2225),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2205),
.Y(n_2307)
);

OA21x2_ASAP7_75t_L g2308 ( 
.A1(n_2215),
.A2(n_74),
.B(n_75),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2202),
.B(n_74),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_2214),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2202),
.B(n_75),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2205),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2225),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2205),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2225),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2225),
.Y(n_2316)
);

AO21x2_ASAP7_75t_L g2317 ( 
.A1(n_2245),
.A2(n_76),
.B(n_77),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2225),
.Y(n_2318)
);

OR2x2_ASAP7_75t_L g2319 ( 
.A(n_2225),
.B(n_76),
.Y(n_2319)
);

CKINVDCx20_ASAP7_75t_R g2320 ( 
.A(n_2206),
.Y(n_2320)
);

BUFx3_ASAP7_75t_L g2321 ( 
.A(n_2214),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2205),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2202),
.B(n_77),
.Y(n_2323)
);

INVx5_ASAP7_75t_L g2324 ( 
.A(n_2199),
.Y(n_2324)
);

OAI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2244),
.A2(n_78),
.B(n_79),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2303),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2326)
);

INVx2_ASAP7_75t_SL g2327 ( 
.A(n_2282),
.Y(n_2327)
);

CKINVDCx20_ASAP7_75t_R g2328 ( 
.A(n_2320),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2261),
.B(n_80),
.Y(n_2329)
);

INVx1_ASAP7_75t_SL g2330 ( 
.A(n_2276),
.Y(n_2330)
);

NOR2x1_ASAP7_75t_SL g2331 ( 
.A(n_2324),
.B(n_2286),
.Y(n_2331)
);

OAI221xp5_ASAP7_75t_L g2332 ( 
.A1(n_2325),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.C(n_85),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_SL g2333 ( 
.A1(n_2301),
.A2(n_83),
.B1(n_85),
.B2(n_82),
.Y(n_2333)
);

AOI221xp5_ASAP7_75t_L g2334 ( 
.A1(n_2273),
.A2(n_87),
.B1(n_81),
.B2(n_86),
.C(n_88),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2251),
.Y(n_2335)
);

AOI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2296),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2302),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2267),
.B(n_90),
.Y(n_2338)
);

OAI22xp33_ASAP7_75t_L g2339 ( 
.A1(n_2269),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_2339)
);

AOI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2295),
.A2(n_849),
.B(n_848),
.Y(n_2340)
);

OR2x6_ASAP7_75t_L g2341 ( 
.A(n_2293),
.B(n_93),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_L g2342 ( 
.A1(n_2270),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2342)
);

OA21x2_ASAP7_75t_L g2343 ( 
.A1(n_2284),
.A2(n_96),
.B(n_98),
.Y(n_2343)
);

AOI22xp33_ASAP7_75t_SL g2344 ( 
.A1(n_2298),
.A2(n_100),
.B1(n_101),
.B2(n_99),
.Y(n_2344)
);

AOI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2289),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_2292),
.B(n_101),
.Y(n_2346)
);

OAI221xp5_ASAP7_75t_L g2347 ( 
.A1(n_2299),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.C(n_105),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2253),
.Y(n_2348)
);

OAI21x1_ASAP7_75t_SL g2349 ( 
.A1(n_2283),
.A2(n_102),
.B(n_103),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_2272),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2255),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2268),
.B(n_107),
.Y(n_2352)
);

AND2x2_ASAP7_75t_SL g2353 ( 
.A(n_2308),
.B(n_108),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2300),
.A2(n_111),
.B1(n_108),
.B2(n_109),
.Y(n_2354)
);

OAI33xp33_ASAP7_75t_L g2355 ( 
.A1(n_2275),
.A2(n_112),
.A3(n_114),
.B1(n_109),
.B2(n_111),
.B3(n_113),
.Y(n_2355)
);

AOI222xp33_ASAP7_75t_L g2356 ( 
.A1(n_2309),
.A2(n_115),
.B1(n_117),
.B2(n_112),
.C1(n_114),
.C2(n_116),
.Y(n_2356)
);

OAI22xp33_ASAP7_75t_L g2357 ( 
.A1(n_2300),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_L g2358 ( 
.A1(n_2294),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2256),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_SL g2360 ( 
.A1(n_2308),
.A2(n_121),
.B1(n_122),
.B2(n_120),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2297),
.A2(n_852),
.B(n_850),
.Y(n_2361)
);

OAI22xp5_ASAP7_75t_L g2362 ( 
.A1(n_2280),
.A2(n_124),
.B1(n_119),
.B2(n_123),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2324),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2363)
);

AOI22xp33_ASAP7_75t_L g2364 ( 
.A1(n_2257),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2252),
.B(n_126),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2305),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2316),
.B(n_127),
.Y(n_2367)
);

OAI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_2324),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2307),
.Y(n_2369)
);

AOI22xp33_ASAP7_75t_L g2370 ( 
.A1(n_2317),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2277),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2250),
.B(n_133),
.Y(n_2372)
);

OAI211xp5_ASAP7_75t_L g2373 ( 
.A1(n_2311),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2312),
.Y(n_2374)
);

AOI221xp5_ASAP7_75t_L g2375 ( 
.A1(n_2323),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.C(n_140),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2314),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2322),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2319),
.A2(n_2306),
.B1(n_2315),
.B2(n_2313),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2318),
.Y(n_2379)
);

OAI21xp33_ASAP7_75t_L g2380 ( 
.A1(n_2290),
.A2(n_138),
.B(n_139),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2262),
.Y(n_2381)
);

INVx4_ASAP7_75t_L g2382 ( 
.A(n_2310),
.Y(n_2382)
);

AOI22xp33_ASAP7_75t_L g2383 ( 
.A1(n_2285),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2258),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2279),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_2385)
);

AOI222xp33_ASAP7_75t_L g2386 ( 
.A1(n_2254),
.A2(n_146),
.B1(n_148),
.B2(n_144),
.C1(n_145),
.C2(n_147),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2260),
.Y(n_2387)
);

AOI22xp33_ASAP7_75t_L g2388 ( 
.A1(n_2278),
.A2(n_149),
.B1(n_145),
.B2(n_148),
.Y(n_2388)
);

OR2x6_ASAP7_75t_L g2389 ( 
.A(n_2321),
.B(n_150),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2266),
.Y(n_2390)
);

OAI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2291),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2274),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2264),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2263),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2265),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2287),
.Y(n_2396)
);

OAI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2259),
.A2(n_155),
.B(n_156),
.Y(n_2397)
);

OAI221xp5_ASAP7_75t_L g2398 ( 
.A1(n_2304),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_2398)
);

OAI22xp33_ASAP7_75t_L g2399 ( 
.A1(n_2288),
.A2(n_161),
.B1(n_157),
.B2(n_159),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2263),
.A2(n_163),
.B1(n_159),
.B2(n_162),
.Y(n_2400)
);

OAI21x1_ASAP7_75t_L g2401 ( 
.A1(n_2271),
.A2(n_162),
.B(n_163),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2281),
.B(n_164),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2251),
.Y(n_2403)
);

AOI221xp5_ASAP7_75t_L g2404 ( 
.A1(n_2303),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2303),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_2405)
);

AOI22xp33_ASAP7_75t_L g2406 ( 
.A1(n_2303),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_2406)
);

OAI211xp5_ASAP7_75t_L g2407 ( 
.A1(n_2303),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2276),
.B(n_172),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2256),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2303),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_2410)
);

AOI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2303),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2267),
.B(n_175),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2256),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2303),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2267),
.B(n_177),
.Y(n_2415)
);

OAI211xp5_ASAP7_75t_SL g2416 ( 
.A1(n_2273),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_2416)
);

AO21x2_ASAP7_75t_L g2417 ( 
.A1(n_2290),
.A2(n_179),
.B(n_180),
.Y(n_2417)
);

OAI221xp5_ASAP7_75t_L g2418 ( 
.A1(n_2303),
.A2(n_184),
.B1(n_181),
.B2(n_183),
.C(n_185),
.Y(n_2418)
);

AOI22xp5_ASAP7_75t_L g2419 ( 
.A1(n_2303),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2256),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2263),
.Y(n_2421)
);

AOI22xp33_ASAP7_75t_L g2422 ( 
.A1(n_2303),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2276),
.B(n_189),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2395),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2332),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2393),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2335),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2353),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2378),
.B(n_192),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2327),
.B(n_193),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2379),
.B(n_2384),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2392),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2348),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2351),
.B(n_193),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2390),
.Y(n_2435)
);

HB1xp67_ASAP7_75t_L g2436 ( 
.A(n_2396),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2421),
.B(n_194),
.Y(n_2437)
);

INVx5_ASAP7_75t_L g2438 ( 
.A(n_2389),
.Y(n_2438)
);

BUFx2_ASAP7_75t_L g2439 ( 
.A(n_2382),
.Y(n_2439)
);

AND2x4_ASAP7_75t_L g2440 ( 
.A(n_2403),
.B(n_194),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2381),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2359),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2387),
.B(n_195),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2366),
.B(n_196),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2369),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_2330),
.B(n_196),
.Y(n_2446)
);

OR2x2_ASAP7_75t_L g2447 ( 
.A(n_2376),
.B(n_197),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2374),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2341),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2377),
.B(n_197),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2409),
.B(n_198),
.Y(n_2451)
);

BUFx2_ASAP7_75t_L g2452 ( 
.A(n_2343),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2413),
.B(n_198),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2420),
.B(n_199),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2372),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2367),
.B(n_199),
.Y(n_2456)
);

BUFx2_ASAP7_75t_L g2457 ( 
.A(n_2341),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2331),
.Y(n_2458)
);

BUFx2_ASAP7_75t_SL g2459 ( 
.A(n_2328),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2343),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2329),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2352),
.B(n_200),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2338),
.B(n_201),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2412),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2415),
.B(n_201),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2417),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2401),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2349),
.Y(n_2468)
);

AOI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2356),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2402),
.B(n_203),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2365),
.B(n_205),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2354),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2389),
.B(n_205),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2346),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2346),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2408),
.B(n_206),
.Y(n_2476)
);

INVx3_ASAP7_75t_L g2477 ( 
.A(n_2423),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2397),
.B(n_206),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2391),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2357),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2363),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2360),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2385),
.B(n_207),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2340),
.B(n_207),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2339),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2334),
.B(n_208),
.Y(n_2486)
);

OR2x2_ASAP7_75t_L g2487 ( 
.A(n_2337),
.B(n_208),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2361),
.B(n_209),
.Y(n_2488)
);

OR2x2_ASAP7_75t_L g2489 ( 
.A(n_2398),
.B(n_209),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2380),
.B(n_210),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2342),
.B(n_210),
.Y(n_2491)
);

AOI22xp33_ASAP7_75t_SL g2492 ( 
.A1(n_2407),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2416),
.Y(n_2493)
);

HB1xp67_ASAP7_75t_L g2494 ( 
.A(n_2368),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2347),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2364),
.B(n_211),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2419),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2362),
.Y(n_2498)
);

INVxp67_ASAP7_75t_L g2499 ( 
.A(n_2418),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2375),
.B(n_213),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2370),
.B(n_214),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2373),
.B(n_214),
.Y(n_2502)
);

HB1xp67_ASAP7_75t_L g2503 ( 
.A(n_2414),
.Y(n_2503)
);

INVx2_ASAP7_75t_SL g2504 ( 
.A(n_2336),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2344),
.B(n_215),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2399),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2386),
.B(n_215),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2333),
.B(n_216),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_L g2509 ( 
.A(n_2394),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2400),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2404),
.B(n_217),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2350),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2383),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2345),
.B(n_218),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2371),
.B(n_2358),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2355),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2326),
.B(n_219),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2388),
.Y(n_2518)
);

HB1xp67_ASAP7_75t_L g2519 ( 
.A(n_2405),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2406),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2410),
.Y(n_2521)
);

HB1xp67_ASAP7_75t_L g2522 ( 
.A(n_2411),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2422),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2392),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2382),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2379),
.B(n_221),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_SL g2527 ( 
.A1(n_2332),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2395),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2395),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2379),
.B(n_222),
.Y(n_2530)
);

AND2x4_ASAP7_75t_SL g2531 ( 
.A(n_2382),
.B(n_224),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2327),
.B(n_225),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2327),
.B(n_225),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2395),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2393),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2379),
.B(n_226),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2392),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2392),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2395),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2382),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2327),
.B(n_226),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2327),
.B(n_227),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2395),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2395),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2379),
.B(n_228),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2327),
.B(n_228),
.Y(n_2546)
);

NOR2x1_ASAP7_75t_SL g2547 ( 
.A(n_2341),
.B(n_229),
.Y(n_2547)
);

AOI22xp33_ASAP7_75t_L g2548 ( 
.A1(n_2332),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2424),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2458),
.B(n_231),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2441),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2467),
.B(n_2439),
.Y(n_2552)
);

NOR3xp33_ASAP7_75t_SL g2553 ( 
.A(n_2507),
.B(n_232),
.C(n_233),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2449),
.B(n_233),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2457),
.B(n_234),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2528),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2455),
.B(n_235),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2529),
.Y(n_2558)
);

INVxp67_ASAP7_75t_L g2559 ( 
.A(n_2494),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2534),
.Y(n_2560)
);

AND2x4_ASAP7_75t_SL g2561 ( 
.A(n_2525),
.B(n_2540),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_2474),
.B(n_235),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2475),
.B(n_236),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2461),
.B(n_2472),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2432),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2539),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2464),
.B(n_236),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2524),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2445),
.B(n_237),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2503),
.B(n_237),
.Y(n_2570)
);

HB1xp67_ASAP7_75t_L g2571 ( 
.A(n_2535),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2468),
.B(n_238),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2499),
.B(n_238),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2543),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2544),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2427),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2537),
.B(n_2538),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2466),
.B(n_2498),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2433),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2435),
.B(n_239),
.Y(n_2580)
);

INVx2_ASAP7_75t_SL g2581 ( 
.A(n_2438),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2480),
.B(n_239),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2436),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2442),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2438),
.B(n_240),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2460),
.B(n_240),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2452),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2448),
.Y(n_2588)
);

OR2x2_ASAP7_75t_L g2589 ( 
.A(n_2452),
.B(n_241),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2426),
.B(n_2438),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2431),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2450),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2497),
.B(n_241),
.Y(n_2593)
);

INVx4_ASAP7_75t_L g2594 ( 
.A(n_2531),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2485),
.B(n_242),
.Y(n_2595)
);

BUFx3_ASAP7_75t_L g2596 ( 
.A(n_2446),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2506),
.B(n_2481),
.Y(n_2597)
);

HB1xp67_ASAP7_75t_L g2598 ( 
.A(n_2447),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2509),
.B(n_2443),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2477),
.B(n_242),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2459),
.B(n_2444),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2451),
.Y(n_2602)
);

INVx1_ASAP7_75t_SL g2603 ( 
.A(n_2546),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2454),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2453),
.B(n_243),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2526),
.B(n_243),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2434),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2530),
.B(n_244),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2536),
.B(n_244),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2545),
.Y(n_2610)
);

NAND2x1_ASAP7_75t_SL g2611 ( 
.A(n_2482),
.B(n_2493),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2429),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2510),
.B(n_245),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2478),
.B(n_245),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2504),
.B(n_246),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2440),
.B(n_246),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2430),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2532),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2479),
.B(n_247),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2533),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2541),
.Y(n_2621)
);

BUFx2_ASAP7_75t_L g2622 ( 
.A(n_2542),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2437),
.Y(n_2623)
);

HB1xp67_ASAP7_75t_L g2624 ( 
.A(n_2519),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2547),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2520),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2518),
.B(n_247),
.Y(n_2627)
);

NAND3xp33_ASAP7_75t_L g2628 ( 
.A(n_2527),
.B(n_248),
.C(n_249),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2521),
.B(n_248),
.Y(n_2629)
);

AND2x4_ASAP7_75t_L g2630 ( 
.A(n_2484),
.B(n_250),
.Y(n_2630)
);

AND2x4_ASAP7_75t_L g2631 ( 
.A(n_2488),
.B(n_250),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2463),
.B(n_251),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2523),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2522),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2495),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_SL g2636 ( 
.A(n_2502),
.B(n_251),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2465),
.B(n_253),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2473),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2512),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2456),
.B(n_253),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2471),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2513),
.B(n_254),
.Y(n_2642)
);

AOI221xp5_ASAP7_75t_L g2643 ( 
.A1(n_2469),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.C(n_257),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2462),
.B(n_255),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2483),
.B(n_257),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_2470),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2476),
.B(n_258),
.Y(n_2647)
);

AND2x4_ASAP7_75t_L g2648 ( 
.A(n_2487),
.B(n_258),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2489),
.B(n_259),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2490),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2516),
.B(n_259),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2505),
.B(n_260),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2515),
.Y(n_2653)
);

INVxp67_ASAP7_75t_SL g2654 ( 
.A(n_2508),
.Y(n_2654)
);

AND2x4_ASAP7_75t_L g2655 ( 
.A(n_2491),
.B(n_261),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2428),
.B(n_261),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2486),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2496),
.B(n_262),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2501),
.B(n_262),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2511),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2500),
.B(n_263),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2492),
.B(n_263),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2517),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2514),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2425),
.B(n_264),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2548),
.B(n_265),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2441),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2458),
.B(n_265),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2461),
.B(n_266),
.Y(n_2669)
);

NAND3xp33_ASAP7_75t_SL g2670 ( 
.A(n_2452),
.B(n_266),
.C(n_267),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2424),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2461),
.B(n_267),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2424),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2441),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2441),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2458),
.B(n_268),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2458),
.B(n_269),
.Y(n_2677)
);

OR2x2_ASAP7_75t_L g2678 ( 
.A(n_2455),
.B(n_269),
.Y(n_2678)
);

INVxp67_ASAP7_75t_SL g2679 ( 
.A(n_2547),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2458),
.B(n_270),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2424),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2461),
.B(n_270),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2458),
.B(n_271),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2461),
.B(n_271),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2441),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2461),
.B(n_272),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2458),
.B(n_272),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2461),
.B(n_273),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2441),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2439),
.B(n_273),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2424),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2438),
.B(n_274),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2455),
.B(n_274),
.Y(n_2693)
);

AND2x4_ASAP7_75t_L g2694 ( 
.A(n_2439),
.B(n_275),
.Y(n_2694)
);

HB1xp67_ASAP7_75t_L g2695 ( 
.A(n_2535),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2458),
.B(n_276),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2458),
.B(n_276),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2458),
.B(n_277),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2535),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2424),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2441),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2438),
.B(n_278),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2458),
.B(n_278),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2424),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2424),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2424),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2458),
.B(n_279),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2458),
.B(n_280),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2424),
.Y(n_2709)
);

OR2x2_ASAP7_75t_L g2710 ( 
.A(n_2455),
.B(n_280),
.Y(n_2710)
);

INVxp67_ASAP7_75t_SL g2711 ( 
.A(n_2547),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_L g2712 ( 
.A(n_2499),
.B(n_281),
.C(n_282),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2424),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2439),
.B(n_281),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2458),
.B(n_284),
.Y(n_2715)
);

INVxp67_ASAP7_75t_SL g2716 ( 
.A(n_2547),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2441),
.Y(n_2717)
);

INVxp67_ASAP7_75t_L g2718 ( 
.A(n_2449),
.Y(n_2718)
);

OAI31xp33_ASAP7_75t_L g2719 ( 
.A1(n_2624),
.A2(n_286),
.A3(n_284),
.B(n_285),
.Y(n_2719)
);

AO21x2_ASAP7_75t_L g2720 ( 
.A1(n_2587),
.A2(n_285),
.B(n_286),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2561),
.B(n_2718),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2571),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2549),
.Y(n_2723)
);

AOI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2634),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_2724)
);

OAI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2553),
.A2(n_287),
.B(n_289),
.Y(n_2725)
);

INVxp67_ASAP7_75t_SL g2726 ( 
.A(n_2611),
.Y(n_2726)
);

NOR2x1_ASAP7_75t_L g2727 ( 
.A(n_2589),
.B(n_290),
.Y(n_2727)
);

HB1xp67_ASAP7_75t_L g2728 ( 
.A(n_2695),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2599),
.B(n_290),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2638),
.B(n_291),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2556),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2653),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_2732)
);

OAI221xp5_ASAP7_75t_SL g2733 ( 
.A1(n_2643),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.C(n_296),
.Y(n_2733)
);

OAI22xp5_ASAP7_75t_SL g2734 ( 
.A1(n_2679),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2558),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_SL g2736 ( 
.A(n_2581),
.B(n_2711),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2692),
.A2(n_297),
.B(n_298),
.Y(n_2737)
);

AOI22xp33_ASAP7_75t_L g2738 ( 
.A1(n_2660),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_2738)
);

AOI21xp33_ASAP7_75t_L g2739 ( 
.A1(n_2716),
.A2(n_300),
.B(n_301),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2699),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2560),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2559),
.B(n_302),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2566),
.Y(n_2743)
);

AOI22xp33_ASAP7_75t_L g2744 ( 
.A1(n_2628),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2635),
.B(n_305),
.Y(n_2745)
);

NAND3xp33_ASAP7_75t_L g2746 ( 
.A(n_2578),
.B(n_306),
.C(n_307),
.Y(n_2746)
);

OAI21xp33_ASAP7_75t_L g2747 ( 
.A1(n_2636),
.A2(n_307),
.B(n_308),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2622),
.B(n_308),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2622),
.B(n_309),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2626),
.B(n_309),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2574),
.Y(n_2751)
);

AND2x4_ASAP7_75t_SL g2752 ( 
.A(n_2594),
.B(n_310),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2575),
.Y(n_2753)
);

OR2x2_ASAP7_75t_L g2754 ( 
.A(n_2633),
.B(n_311),
.Y(n_2754)
);

AOI22xp33_ASAP7_75t_L g2755 ( 
.A1(n_2657),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_2755)
);

OAI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2702),
.A2(n_312),
.B(n_313),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2576),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2590),
.Y(n_2758)
);

BUFx2_ASAP7_75t_L g2759 ( 
.A(n_2625),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2597),
.B(n_314),
.Y(n_2760)
);

AND2x4_ASAP7_75t_L g2761 ( 
.A(n_2601),
.B(n_314),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2646),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2552),
.B(n_316),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2646),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2641),
.B(n_316),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2612),
.B(n_317),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2579),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2671),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2673),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2598),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2654),
.B(n_318),
.Y(n_2771)
);

AOI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2639),
.A2(n_2663),
.B1(n_2664),
.B2(n_2651),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2604),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2623),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2681),
.Y(n_2775)
);

OAI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2564),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2617),
.B(n_319),
.Y(n_2777)
);

NOR3xp33_ASAP7_75t_L g2778 ( 
.A(n_2670),
.B(n_321),
.C(n_322),
.Y(n_2778)
);

HB1xp67_ASAP7_75t_L g2779 ( 
.A(n_2583),
.Y(n_2779)
);

AOI21xp33_ASAP7_75t_L g2780 ( 
.A1(n_2665),
.A2(n_321),
.B(n_322),
.Y(n_2780)
);

INVx4_ASAP7_75t_L g2781 ( 
.A(n_2585),
.Y(n_2781)
);

INVx2_ASAP7_75t_SL g2782 ( 
.A(n_2596),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2691),
.Y(n_2783)
);

OAI31xp33_ASAP7_75t_L g2784 ( 
.A1(n_2712),
.A2(n_325),
.A3(n_323),
.B(n_324),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2607),
.B(n_324),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2700),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2704),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2551),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_2584),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2667),
.B(n_325),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2705),
.Y(n_2791)
);

OR2x2_ASAP7_75t_L g2792 ( 
.A(n_2610),
.B(n_326),
.Y(n_2792)
);

OR2x6_ASAP7_75t_L g2793 ( 
.A(n_2554),
.B(n_326),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2706),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2674),
.B(n_327),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2586),
.B(n_327),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2650),
.B(n_328),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2675),
.B(n_328),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2709),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2685),
.B(n_329),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2689),
.B(n_2701),
.Y(n_2801)
);

AO21x2_ASAP7_75t_L g2802 ( 
.A1(n_2570),
.A2(n_329),
.B(n_330),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2717),
.B(n_2592),
.Y(n_2803)
);

INVxp67_ASAP7_75t_SL g2804 ( 
.A(n_2642),
.Y(n_2804)
);

OAI22xp33_ASAP7_75t_L g2805 ( 
.A1(n_2603),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2614),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_2806)
);

AOI21xp33_ASAP7_75t_L g2807 ( 
.A1(n_2656),
.A2(n_333),
.B(n_334),
.Y(n_2807)
);

AOI31xp33_ASAP7_75t_L g2808 ( 
.A1(n_2662),
.A2(n_336),
.A3(n_334),
.B(n_335),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2577),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2565),
.Y(n_2810)
);

AND2x4_ASAP7_75t_L g2811 ( 
.A(n_2618),
.B(n_337),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2568),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2713),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2620),
.Y(n_2814)
);

AND4x1_ASAP7_75t_L g2815 ( 
.A(n_2573),
.B(n_340),
.C(n_338),
.D(n_339),
.Y(n_2815)
);

NAND3xp33_ASAP7_75t_L g2816 ( 
.A(n_2661),
.B(n_338),
.C(n_339),
.Y(n_2816)
);

AO21x2_ASAP7_75t_L g2817 ( 
.A1(n_2669),
.A2(n_340),
.B(n_341),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2588),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2629),
.Y(n_2819)
);

INVx1_ASAP7_75t_SL g2820 ( 
.A(n_2555),
.Y(n_2820)
);

NAND2x1p5_ASAP7_75t_SL g2821 ( 
.A(n_2550),
.B(n_2668),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2591),
.Y(n_2822)
);

INVx4_ASAP7_75t_L g2823 ( 
.A(n_2690),
.Y(n_2823)
);

INVx4_ASAP7_75t_L g2824 ( 
.A(n_2694),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2602),
.Y(n_2825)
);

NAND4xp25_ASAP7_75t_L g2826 ( 
.A(n_2593),
.B(n_343),
.C(n_344),
.D(n_342),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2621),
.Y(n_2827)
);

AOI221xp5_ASAP7_75t_L g2828 ( 
.A1(n_2619),
.A2(n_345),
.B1(n_341),
.B2(n_344),
.C(n_346),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2613),
.B(n_346),
.Y(n_2829)
);

OAI31xp33_ASAP7_75t_SL g2830 ( 
.A1(n_2649),
.A2(n_2582),
.A3(n_2666),
.B(n_2659),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2580),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2676),
.B(n_347),
.Y(n_2832)
);

HB1xp67_ASAP7_75t_L g2833 ( 
.A(n_2678),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2569),
.Y(n_2834)
);

OR2x2_ASAP7_75t_L g2835 ( 
.A(n_2693),
.B(n_347),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2557),
.B(n_348),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2714),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2710),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2672),
.B(n_349),
.Y(n_2839)
);

NOR3xp33_ASAP7_75t_L g2840 ( 
.A(n_2682),
.B(n_349),
.C(n_351),
.Y(n_2840)
);

INVx1_ASAP7_75t_SL g2841 ( 
.A(n_2615),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2770),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2721),
.B(n_2677),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2781),
.B(n_2680),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2752),
.Y(n_2845)
);

INVx2_ASAP7_75t_SL g2846 ( 
.A(n_2837),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2820),
.B(n_2841),
.Y(n_2847)
);

AND2x4_ASAP7_75t_L g2848 ( 
.A(n_2758),
.B(n_2683),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2782),
.B(n_2687),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2722),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2823),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2759),
.B(n_2696),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2728),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2762),
.B(n_2697),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2764),
.B(n_2698),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2804),
.B(n_2572),
.Y(n_2856)
);

OAI211xp5_ASAP7_75t_SL g2857 ( 
.A1(n_2772),
.A2(n_2645),
.B(n_2606),
.C(n_2609),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2740),
.Y(n_2858)
);

AND2x4_ASAP7_75t_L g2859 ( 
.A(n_2824),
.B(n_2703),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2831),
.B(n_2707),
.Y(n_2860)
);

O2A1O1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2808),
.A2(n_2684),
.B(n_2688),
.C(n_2686),
.Y(n_2861)
);

INVxp67_ASAP7_75t_SL g2862 ( 
.A(n_2726),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2830),
.B(n_2708),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2779),
.Y(n_2864)
);

OR2x2_ASAP7_75t_L g2865 ( 
.A(n_2833),
.B(n_2608),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2834),
.B(n_2715),
.Y(n_2866)
);

INVx1_ASAP7_75t_SL g2867 ( 
.A(n_2748),
.Y(n_2867)
);

INVx1_ASAP7_75t_SL g2868 ( 
.A(n_2749),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2819),
.B(n_2595),
.Y(n_2869)
);

NAND2xp33_ASAP7_75t_R g2870 ( 
.A(n_2725),
.B(n_2648),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2821),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2809),
.B(n_2567),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2761),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2838),
.B(n_2627),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2803),
.B(n_2630),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2802),
.B(n_2631),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2789),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2736),
.B(n_2600),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2723),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2731),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2788),
.B(n_2652),
.Y(n_2881)
);

OAI222xp33_ASAP7_75t_L g2882 ( 
.A1(n_2733),
.A2(n_2640),
.B1(n_2658),
.B2(n_2605),
.C1(n_2644),
.C2(n_2655),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2817),
.B(n_2562),
.Y(n_2883)
);

OR2x2_ASAP7_75t_L g2884 ( 
.A(n_2773),
.B(n_2563),
.Y(n_2884)
);

OAI31xp33_ASAP7_75t_L g2885 ( 
.A1(n_2734),
.A2(n_2616),
.A3(n_2647),
.B(n_2637),
.Y(n_2885)
);

BUFx2_ASAP7_75t_L g2886 ( 
.A(n_2727),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2735),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2763),
.B(n_2632),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2840),
.B(n_2814),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2774),
.B(n_351),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2729),
.B(n_352),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2720),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2760),
.B(n_352),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2810),
.Y(n_2894)
);

NAND3xp33_ASAP7_75t_L g2895 ( 
.A(n_2778),
.B(n_353),
.C(n_354),
.Y(n_2895)
);

OR2x2_ASAP7_75t_L g2896 ( 
.A(n_2827),
.B(n_353),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2741),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2743),
.Y(n_2898)
);

NAND3xp33_ASAP7_75t_L g2899 ( 
.A(n_2784),
.B(n_354),
.C(n_355),
.Y(n_2899)
);

INVx1_ASAP7_75t_SL g2900 ( 
.A(n_2793),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2797),
.B(n_356),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2900),
.B(n_2825),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2862),
.B(n_2730),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2851),
.B(n_2801),
.Y(n_2904)
);

INVx3_ASAP7_75t_SL g2905 ( 
.A(n_2845),
.Y(n_2905)
);

CKINVDCx16_ASAP7_75t_R g2906 ( 
.A(n_2870),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2886),
.B(n_2766),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2843),
.B(n_2793),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2842),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2852),
.B(n_2812),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2867),
.B(n_2745),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2868),
.B(n_2765),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2850),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2853),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2859),
.Y(n_2915)
);

INVxp67_ASAP7_75t_L g2916 ( 
.A(n_2892),
.Y(n_2916)
);

OR2x2_ASAP7_75t_L g2917 ( 
.A(n_2871),
.B(n_2771),
.Y(n_2917)
);

AOI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2899),
.A2(n_2846),
.B1(n_2878),
.B2(n_2859),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2844),
.B(n_2832),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2882),
.B(n_2839),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2885),
.B(n_2719),
.Y(n_2921)
);

INVx2_ASAP7_75t_SL g2922 ( 
.A(n_2849),
.Y(n_2922)
);

INVx3_ASAP7_75t_L g2923 ( 
.A(n_2848),
.Y(n_2923)
);

OR2x2_ASAP7_75t_L g2924 ( 
.A(n_2874),
.B(n_2742),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2875),
.B(n_2790),
.Y(n_2925)
);

AOI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2895),
.A2(n_2747),
.B1(n_2746),
.B2(n_2776),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2848),
.B(n_2751),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2858),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2854),
.B(n_2795),
.Y(n_2929)
);

INVx1_ASAP7_75t_SL g2930 ( 
.A(n_2883),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2864),
.Y(n_2931)
);

CKINVDCx11_ASAP7_75t_R g2932 ( 
.A(n_2873),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2888),
.B(n_2822),
.Y(n_2933)
);

INVxp67_ASAP7_75t_L g2934 ( 
.A(n_2904),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2902),
.Y(n_2935)
);

OAI22xp33_ASAP7_75t_R g2936 ( 
.A1(n_2920),
.A2(n_2865),
.B1(n_2877),
.B2(n_2884),
.Y(n_2936)
);

OR2x2_ASAP7_75t_L g2937 ( 
.A(n_2903),
.B(n_2930),
.Y(n_2937)
);

INVx2_ASAP7_75t_SL g2938 ( 
.A(n_2905),
.Y(n_2938)
);

OAI22xp33_ASAP7_75t_SL g2939 ( 
.A1(n_2906),
.A2(n_2863),
.B1(n_2889),
.B2(n_2876),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2923),
.Y(n_2940)
);

OR2x2_ASAP7_75t_L g2941 ( 
.A(n_2907),
.B(n_2912),
.Y(n_2941)
);

HB1xp67_ASAP7_75t_L g2942 ( 
.A(n_2915),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2908),
.B(n_2855),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2921),
.A2(n_2869),
.B1(n_2881),
.B2(n_2847),
.Y(n_2944)
);

OAI21xp5_ASAP7_75t_SL g2945 ( 
.A1(n_2926),
.A2(n_2744),
.B(n_2756),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2909),
.Y(n_2946)
);

A2O1A1Ixp33_ASAP7_75t_L g2947 ( 
.A1(n_2918),
.A2(n_2861),
.B(n_2737),
.C(n_2739),
.Y(n_2947)
);

A2O1A1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2916),
.A2(n_2816),
.B(n_2828),
.C(n_2807),
.Y(n_2948)
);

OR2x2_ASAP7_75t_L g2949 ( 
.A(n_2917),
.B(n_2856),
.Y(n_2949)
);

AND2x4_ASAP7_75t_L g2950 ( 
.A(n_2922),
.B(n_2860),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2913),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2919),
.B(n_2872),
.Y(n_2952)
);

INVx1_ASAP7_75t_SL g2953 ( 
.A(n_2932),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2942),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2953),
.Y(n_2955)
);

INVxp67_ASAP7_75t_L g2956 ( 
.A(n_2938),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2950),
.B(n_2929),
.Y(n_2957)
);

O2A1O1Ixp5_ASAP7_75t_L g2958 ( 
.A1(n_2947),
.A2(n_2940),
.B(n_2948),
.C(n_2914),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2943),
.B(n_2925),
.Y(n_2959)
);

INVx2_ASAP7_75t_SL g2960 ( 
.A(n_2937),
.Y(n_2960)
);

INVxp67_ASAP7_75t_L g2961 ( 
.A(n_2952),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2936),
.A2(n_2910),
.B1(n_2924),
.B2(n_2928),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2949),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2955),
.B(n_2934),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2959),
.B(n_2944),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2954),
.Y(n_2966)
);

AOI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2956),
.A2(n_2945),
.B1(n_2939),
.B2(n_2935),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2960),
.Y(n_2968)
);

AOI221xp5_ASAP7_75t_L g2969 ( 
.A1(n_2958),
.A2(n_2931),
.B1(n_2951),
.B2(n_2946),
.C(n_2927),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2963),
.B(n_2927),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2957),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2961),
.Y(n_2972)
);

AOI221xp5_ASAP7_75t_L g2973 ( 
.A1(n_2969),
.A2(n_2962),
.B1(n_2933),
.B2(n_2911),
.C(n_2898),
.Y(n_2973)
);

AOI322xp5_ASAP7_75t_L g2974 ( 
.A1(n_2967),
.A2(n_2805),
.A3(n_2780),
.B1(n_2901),
.B2(n_2724),
.C1(n_2879),
.C2(n_2887),
.Y(n_2974)
);

AOI21xp33_ASAP7_75t_SL g2975 ( 
.A1(n_2965),
.A2(n_2941),
.B(n_2896),
.Y(n_2975)
);

AOI322xp5_ASAP7_75t_L g2976 ( 
.A1(n_2968),
.A2(n_2880),
.A3(n_2897),
.B1(n_2732),
.B2(n_2755),
.C1(n_2738),
.C2(n_2866),
.Y(n_2976)
);

AOI311xp33_ASAP7_75t_L g2977 ( 
.A1(n_2966),
.A2(n_2806),
.A3(n_2767),
.B(n_2768),
.C(n_2757),
.Y(n_2977)
);

AOI221x1_ASAP7_75t_L g2978 ( 
.A1(n_2964),
.A2(n_2971),
.B1(n_2972),
.B2(n_2970),
.C(n_2894),
.Y(n_2978)
);

AOI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2965),
.A2(n_2857),
.B(n_2829),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2970),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2970),
.B(n_2891),
.Y(n_2981)
);

NOR4xp25_ASAP7_75t_L g2982 ( 
.A(n_2969),
.B(n_2890),
.C(n_2826),
.D(n_2796),
.Y(n_2982)
);

AOI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2968),
.A2(n_2753),
.B1(n_2775),
.B2(n_2769),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2970),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2970),
.B(n_2893),
.Y(n_2985)
);

NAND4xp25_ASAP7_75t_L g2986 ( 
.A(n_2967),
.B(n_2836),
.C(n_2792),
.D(n_2785),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2970),
.B(n_2783),
.Y(n_2987)
);

O2A1O1Ixp5_ASAP7_75t_L g2988 ( 
.A1(n_2965),
.A2(n_2787),
.B(n_2791),
.C(n_2786),
.Y(n_2988)
);

OAI211xp5_ASAP7_75t_L g2989 ( 
.A1(n_2967),
.A2(n_2835),
.B(n_2754),
.C(n_2750),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2970),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2980),
.B(n_2794),
.Y(n_2991)
);

OAI321xp33_ASAP7_75t_L g2992 ( 
.A1(n_2973),
.A2(n_2800),
.A3(n_2798),
.B1(n_2818),
.B2(n_2813),
.C(n_2799),
.Y(n_2992)
);

OAI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2979),
.A2(n_2974),
.B(n_2981),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2990),
.B(n_2777),
.Y(n_2994)
);

AOI21xp33_ASAP7_75t_L g2995 ( 
.A1(n_2989),
.A2(n_2811),
.B(n_2815),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2984),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_2996)
);

OAI221xp5_ASAP7_75t_SL g2997 ( 
.A1(n_2983),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.C(n_360),
.Y(n_2997)
);

A2O1A1Ixp33_ASAP7_75t_L g2998 ( 
.A1(n_2976),
.A2(n_362),
.B(n_363),
.C(n_361),
.Y(n_2998)
);

AOI21xp33_ASAP7_75t_L g2999 ( 
.A1(n_2985),
.A2(n_363),
.B(n_361),
.Y(n_2999)
);

AOI322xp5_ASAP7_75t_L g3000 ( 
.A1(n_2987),
.A2(n_368),
.A3(n_367),
.B1(n_365),
.B2(n_359),
.C1(n_364),
.C2(n_366),
.Y(n_3000)
);

INVxp33_ASAP7_75t_L g3001 ( 
.A(n_2986),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2988),
.Y(n_3002)
);

OAI22xp5_ASAP7_75t_L g3003 ( 
.A1(n_2975),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_3003)
);

OAI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2978),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2977),
.A2(n_2982),
.B1(n_371),
.B2(n_369),
.Y(n_3005)
);

OAI21xp5_ASAP7_75t_L g3006 ( 
.A1(n_2979),
.A2(n_370),
.B(n_371),
.Y(n_3006)
);

OAI211xp5_ASAP7_75t_L g3007 ( 
.A1(n_2973),
.A2(n_373),
.B(n_370),
.C(n_372),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2981),
.B(n_372),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2980),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3009)
);

NAND4xp25_ASAP7_75t_L g3010 ( 
.A(n_2973),
.B(n_376),
.C(n_374),
.D(n_375),
.Y(n_3010)
);

A2O1A1Ixp33_ASAP7_75t_L g3011 ( 
.A1(n_2995),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2994),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_3003),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_3002),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_3008),
.Y(n_3015)
);

AOI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2993),
.A2(n_3004),
.B(n_2992),
.Y(n_3016)
);

NOR4xp25_ASAP7_75t_SL g3017 ( 
.A(n_2998),
.B(n_381),
.C(n_377),
.D(n_380),
.Y(n_3017)
);

AOI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_3010),
.A2(n_3001),
.B1(n_3007),
.B2(n_3005),
.Y(n_3018)
);

OAI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2991),
.A2(n_382),
.B1(n_383),
.B2(n_381),
.Y(n_3019)
);

OAI221xp5_ASAP7_75t_SL g3020 ( 
.A1(n_3000),
.A2(n_383),
.B1(n_380),
.B2(n_382),
.C(n_384),
.Y(n_3020)
);

O2A1O1Ixp33_ASAP7_75t_L g3021 ( 
.A1(n_3006),
.A2(n_388),
.B(n_384),
.C(n_385),
.Y(n_3021)
);

AOI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_3009),
.A2(n_390),
.B1(n_385),
.B2(n_389),
.Y(n_3022)
);

AOI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2999),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_3023)
);

XOR2x2_ASAP7_75t_L g3024 ( 
.A(n_2997),
.B(n_391),
.Y(n_3024)
);

AOI21xp33_ASAP7_75t_SL g3025 ( 
.A1(n_2996),
.A2(n_392),
.B(n_393),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_3005),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_3026)
);

OAI21xp33_ASAP7_75t_L g3027 ( 
.A1(n_3001),
.A2(n_394),
.B(n_395),
.Y(n_3027)
);

INVx1_ASAP7_75t_SL g3028 ( 
.A(n_2994),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2994),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2994),
.B(n_396),
.Y(n_3030)
);

AOI22xp33_ASAP7_75t_L g3031 ( 
.A1(n_3001),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_3005),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3032)
);

AOI221xp5_ASAP7_75t_L g3033 ( 
.A1(n_3026),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.C(n_402),
.Y(n_3033)
);

OA22x2_ASAP7_75t_L g3034 ( 
.A1(n_3018),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_3028),
.B(n_403),
.Y(n_3035)
);

XNOR2xp5_ASAP7_75t_L g3036 ( 
.A(n_3024),
.B(n_404),
.Y(n_3036)
);

OAI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_3016),
.A2(n_3011),
.B(n_3032),
.Y(n_3037)
);

A2O1A1Ixp33_ASAP7_75t_L g3038 ( 
.A1(n_3021),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_3030),
.Y(n_3039)
);

OAI221xp5_ASAP7_75t_L g3040 ( 
.A1(n_3014),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.C(n_408),
.Y(n_3040)
);

XNOR2xp5_ASAP7_75t_L g3041 ( 
.A(n_3029),
.B(n_408),
.Y(n_3041)
);

NAND5xp2_ASAP7_75t_L g3042 ( 
.A(n_3013),
.B(n_411),
.C(n_409),
.D(n_410),
.E(n_412),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_3012),
.B(n_409),
.Y(n_3043)
);

AOI22xp33_ASAP7_75t_L g3044 ( 
.A1(n_3015),
.A2(n_413),
.B1(n_410),
.B2(n_411),
.Y(n_3044)
);

INVx1_ASAP7_75t_SL g3045 ( 
.A(n_3022),
.Y(n_3045)
);

NAND3xp33_ASAP7_75t_SL g3046 ( 
.A(n_3017),
.B(n_413),
.C(n_414),
.Y(n_3046)
);

AOI22xp5_ASAP7_75t_L g3047 ( 
.A1(n_3027),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_3023),
.Y(n_3048)
);

AOI21xp33_ASAP7_75t_L g3049 ( 
.A1(n_3019),
.A2(n_415),
.B(n_416),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_3031),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_3050)
);

O2A1O1Ixp33_ASAP7_75t_L g3051 ( 
.A1(n_3020),
.A2(n_422),
.B(n_417),
.C(n_421),
.Y(n_3051)
);

HB1xp67_ASAP7_75t_L g3052 ( 
.A(n_3025),
.Y(n_3052)
);

OAI21xp33_ASAP7_75t_SL g3053 ( 
.A1(n_3018),
.A2(n_421),
.B(n_424),
.Y(n_3053)
);

AND2x4_ASAP7_75t_L g3054 ( 
.A(n_3012),
.B(n_425),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_3028),
.B(n_424),
.Y(n_3055)
);

AOI221xp5_ASAP7_75t_L g3056 ( 
.A1(n_3026),
.A2(n_428),
.B1(n_425),
.B2(n_427),
.C(n_429),
.Y(n_3056)
);

AOI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_3028),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_3028),
.B(n_430),
.Y(n_3058)
);

OAI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_3016),
.A2(n_433),
.B(n_432),
.Y(n_3059)
);

AOI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_3028),
.A2(n_433),
.B1(n_430),
.B2(n_432),
.Y(n_3060)
);

INVxp67_ASAP7_75t_L g3061 ( 
.A(n_3030),
.Y(n_3061)
);

AOI21xp33_ASAP7_75t_SL g3062 ( 
.A1(n_3026),
.A2(n_434),
.B(n_435),
.Y(n_3062)
);

XNOR2x1_ASAP7_75t_L g3063 ( 
.A(n_3024),
.B(n_434),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_3012),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_3064)
);

OAI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_3018),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_3065)
);

CKINVDCx16_ASAP7_75t_R g3066 ( 
.A(n_3018),
.Y(n_3066)
);

INVxp33_ASAP7_75t_SL g3067 ( 
.A(n_3018),
.Y(n_3067)
);

AOI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_3028),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_3068)
);

NOR3xp33_ASAP7_75t_L g3069 ( 
.A(n_3029),
.B(n_442),
.C(n_441),
.Y(n_3069)
);

AOI31xp33_ASAP7_75t_L g3070 ( 
.A1(n_3028),
.A2(n_449),
.A3(n_457),
.B(n_440),
.Y(n_3070)
);

A2O1A1Ixp33_ASAP7_75t_L g3071 ( 
.A1(n_3016),
.A2(n_444),
.B(n_442),
.C(n_443),
.Y(n_3071)
);

AOI22xp5_ASAP7_75t_L g3072 ( 
.A1(n_3067),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_3072)
);

OAI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_3066),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_3073)
);

AOI31xp33_ASAP7_75t_L g3074 ( 
.A1(n_3046),
.A2(n_451),
.A3(n_449),
.B(n_450),
.Y(n_3074)
);

AO22x2_ASAP7_75t_SL g3075 ( 
.A1(n_3069),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3041),
.Y(n_3076)
);

NOR2xp67_ASAP7_75t_L g3077 ( 
.A(n_3042),
.B(n_452),
.Y(n_3077)
);

AOI31xp33_ASAP7_75t_L g3078 ( 
.A1(n_3036),
.A2(n_455),
.A3(n_453),
.B(n_454),
.Y(n_3078)
);

INVxp33_ASAP7_75t_L g3079 ( 
.A(n_3063),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_3034),
.Y(n_3080)
);

OR2x2_ASAP7_75t_L g3081 ( 
.A(n_3035),
.B(n_454),
.Y(n_3081)
);

AO22x2_ASAP7_75t_L g3082 ( 
.A1(n_3045),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_3082)
);

HB1xp67_ASAP7_75t_L g3083 ( 
.A(n_3054),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_3054),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3070),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_3052),
.B(n_456),
.Y(n_3086)
);

OAI22xp5_ASAP7_75t_L g3087 ( 
.A1(n_3047),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_3087)
);

AOI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_3048),
.A2(n_3050),
.B1(n_3053),
.B2(n_3059),
.Y(n_3088)
);

NOR2x1_ASAP7_75t_L g3089 ( 
.A(n_3058),
.B(n_458),
.Y(n_3089)
);

NOR2x1_ASAP7_75t_L g3090 ( 
.A(n_3055),
.B(n_459),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3043),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3037),
.B(n_460),
.Y(n_3092)
);

AOI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_3065),
.A2(n_3061),
.B1(n_3039),
.B2(n_3056),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3057),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_3060),
.Y(n_3095)
);

INVx1_ASAP7_75t_SL g3096 ( 
.A(n_3068),
.Y(n_3096)
);

OAI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_3071),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3051),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3062),
.B(n_462),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3038),
.Y(n_3100)
);

NOR2x1_ASAP7_75t_L g3101 ( 
.A(n_3040),
.B(n_463),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_3033),
.B(n_464),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3064),
.Y(n_3103)
);

AND3x4_ASAP7_75t_L g3104 ( 
.A(n_3049),
.B(n_465),
.C(n_466),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3044),
.Y(n_3105)
);

NOR2x1_ASAP7_75t_L g3106 ( 
.A(n_3046),
.B(n_465),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3052),
.B(n_467),
.Y(n_3107)
);

NOR2xp67_ASAP7_75t_L g3108 ( 
.A(n_3046),
.B(n_469),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_3052),
.B(n_469),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_3067),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_3110)
);

AOI22xp5_ASAP7_75t_L g3111 ( 
.A1(n_3067),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_3111)
);

AND2x4_ASAP7_75t_L g3112 ( 
.A(n_3035),
.B(n_473),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3041),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_3067),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_3114)
);

NOR2x1_ASAP7_75t_L g3115 ( 
.A(n_3046),
.B(n_474),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3041),
.Y(n_3116)
);

INVxp33_ASAP7_75t_L g3117 ( 
.A(n_3041),
.Y(n_3117)
);

NOR2x1_ASAP7_75t_L g3118 ( 
.A(n_3046),
.B(n_475),
.Y(n_3118)
);

NOR2x1_ASAP7_75t_L g3119 ( 
.A(n_3046),
.B(n_476),
.Y(n_3119)
);

BUFx3_ASAP7_75t_L g3120 ( 
.A(n_3084),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_3092),
.B(n_477),
.Y(n_3121)
);

NOR2x1_ASAP7_75t_L g3122 ( 
.A(n_3090),
.B(n_477),
.Y(n_3122)
);

OAI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_3072),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_3082),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3082),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_3110),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_3126)
);

AOI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_3077),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_3074),
.B(n_481),
.Y(n_3128)
);

NOR2x1_ASAP7_75t_L g3129 ( 
.A(n_3106),
.B(n_483),
.Y(n_3129)
);

AOI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_3108),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_3130)
);

NOR2xp33_ASAP7_75t_L g3131 ( 
.A(n_3078),
.B(n_484),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3083),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3075),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_3086),
.B(n_485),
.Y(n_3134)
);

NOR3xp33_ASAP7_75t_L g3135 ( 
.A(n_3098),
.B(n_494),
.C(n_486),
.Y(n_3135)
);

NOR2x1p5_ASAP7_75t_L g3136 ( 
.A(n_3085),
.B(n_487),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3107),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3109),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_3081),
.B(n_487),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_3112),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3115),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3118),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_3119),
.B(n_488),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_3080),
.B(n_489),
.Y(n_3144)
);

NAND4xp75_ASAP7_75t_L g3145 ( 
.A(n_3089),
.B(n_490),
.C(n_488),
.D(n_489),
.Y(n_3145)
);

INVx1_ASAP7_75t_SL g3146 ( 
.A(n_3099),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3073),
.Y(n_3147)
);

NOR2x1_ASAP7_75t_L g3148 ( 
.A(n_3104),
.B(n_490),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3111),
.Y(n_3149)
);

AND2x4_ASAP7_75t_L g3150 ( 
.A(n_3076),
.B(n_491),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_3117),
.B(n_491),
.Y(n_3151)
);

AOI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_3096),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_SL g3153 ( 
.A(n_3097),
.B(n_493),
.Y(n_3153)
);

NAND4xp75_ASAP7_75t_L g3154 ( 
.A(n_3101),
.B(n_3093),
.C(n_3102),
.D(n_3113),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3114),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3088),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3094),
.Y(n_3157)
);

XOR2x1_ASAP7_75t_L g3158 ( 
.A(n_3116),
.B(n_495),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3095),
.Y(n_3159)
);

HB1xp67_ASAP7_75t_L g3160 ( 
.A(n_3087),
.Y(n_3160)
);

NOR2x1_ASAP7_75t_L g3161 ( 
.A(n_3100),
.B(n_495),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3103),
.Y(n_3162)
);

XNOR2xp5_ASAP7_75t_L g3163 ( 
.A(n_3079),
.B(n_496),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3105),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3091),
.B(n_496),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3082),
.Y(n_3166)
);

XOR2xp5_ASAP7_75t_L g3167 ( 
.A(n_3117),
.B(n_497),
.Y(n_3167)
);

NAND4xp75_ASAP7_75t_L g3168 ( 
.A(n_3090),
.B(n_499),
.C(n_497),
.D(n_498),
.Y(n_3168)
);

NOR2x1_ASAP7_75t_L g3169 ( 
.A(n_3090),
.B(n_498),
.Y(n_3169)
);

NOR2x1_ASAP7_75t_L g3170 ( 
.A(n_3090),
.B(n_499),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3092),
.B(n_500),
.Y(n_3171)
);

INVx2_ASAP7_75t_SL g3172 ( 
.A(n_3083),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_3077),
.B(n_500),
.Y(n_3173)
);

XNOR2xp5_ASAP7_75t_L g3174 ( 
.A(n_3077),
.B(n_501),
.Y(n_3174)
);

NAND4xp75_ASAP7_75t_L g3175 ( 
.A(n_3090),
.B(n_503),
.C(n_501),
.D(n_502),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3082),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3082),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3082),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3082),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3082),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_3074),
.B(n_502),
.Y(n_3181)
);

AO22x2_ASAP7_75t_L g3182 ( 
.A1(n_3125),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_3182)
);

OAI211xp5_ASAP7_75t_SL g3183 ( 
.A1(n_3132),
.A2(n_506),
.B(n_504),
.C(n_505),
.Y(n_3183)
);

AOI221xp5_ASAP7_75t_L g3184 ( 
.A1(n_3172),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.C(n_509),
.Y(n_3184)
);

OAI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_3127),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.Y(n_3185)
);

NAND3xp33_ASAP7_75t_L g3186 ( 
.A(n_3135),
.B(n_510),
.C(n_511),
.Y(n_3186)
);

OAI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_3130),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_3187)
);

AOI21xp33_ASAP7_75t_SL g3188 ( 
.A1(n_3166),
.A2(n_513),
.B(n_514),
.Y(n_3188)
);

OAI211xp5_ASAP7_75t_SL g3189 ( 
.A1(n_3156),
.A2(n_516),
.B(n_514),
.C(n_515),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_L g3190 ( 
.A1(n_3120),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3167),
.Y(n_3191)
);

OAI221xp5_ASAP7_75t_L g3192 ( 
.A1(n_3144),
.A2(n_3174),
.B1(n_3173),
.B2(n_3133),
.C(n_3153),
.Y(n_3192)
);

OAI22xp5_ASAP7_75t_SL g3193 ( 
.A1(n_3141),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_3193)
);

AOI31xp33_ASAP7_75t_L g3194 ( 
.A1(n_3129),
.A2(n_522),
.A3(n_520),
.B(n_521),
.Y(n_3194)
);

NOR3xp33_ASAP7_75t_SL g3195 ( 
.A(n_3154),
.B(n_3142),
.C(n_3162),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_3151),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_3196)
);

OAI221xp5_ASAP7_75t_L g3197 ( 
.A1(n_3176),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.C(n_526),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3148),
.B(n_523),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3163),
.Y(n_3199)
);

NAND3xp33_ASAP7_75t_SL g3200 ( 
.A(n_3178),
.B(n_3180),
.C(n_3179),
.Y(n_3200)
);

NAND3xp33_ASAP7_75t_L g3201 ( 
.A(n_3122),
.B(n_525),
.C(n_526),
.Y(n_3201)
);

NAND4xp75_ASAP7_75t_L g3202 ( 
.A(n_3161),
.B(n_529),
.C(n_527),
.D(n_528),
.Y(n_3202)
);

NOR3x2_ASAP7_75t_L g3203 ( 
.A(n_3168),
.B(n_527),
.C(n_528),
.Y(n_3203)
);

XNOR2xp5_ASAP7_75t_L g3204 ( 
.A(n_3158),
.B(n_529),
.Y(n_3204)
);

NAND3xp33_ASAP7_75t_SL g3205 ( 
.A(n_3124),
.B(n_531),
.C(n_532),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3157),
.A2(n_534),
.B1(n_531),
.B2(n_533),
.Y(n_3206)
);

NAND4xp25_ASAP7_75t_L g3207 ( 
.A(n_3164),
.B(n_535),
.C(n_533),
.D(n_534),
.Y(n_3207)
);

INVx1_ASAP7_75t_SL g3208 ( 
.A(n_3175),
.Y(n_3208)
);

OAI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_3143),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_3209)
);

OR3x2_ASAP7_75t_L g3210 ( 
.A(n_3137),
.B(n_536),
.C(n_538),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_3139),
.B(n_539),
.Y(n_3211)
);

AO22x2_ASAP7_75t_L g3212 ( 
.A1(n_3177),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3169),
.Y(n_3213)
);

OAI21xp33_ASAP7_75t_SL g3214 ( 
.A1(n_3170),
.A2(n_540),
.B(n_541),
.Y(n_3214)
);

OAI211xp5_ASAP7_75t_L g3215 ( 
.A1(n_3128),
.A2(n_545),
.B(n_542),
.C(n_543),
.Y(n_3215)
);

OAI211xp5_ASAP7_75t_L g3216 ( 
.A1(n_3181),
.A2(n_545),
.B(n_542),
.C(n_543),
.Y(n_3216)
);

AOI221xp5_ASAP7_75t_L g3217 ( 
.A1(n_3147),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.C(n_549),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_3150),
.Y(n_3218)
);

O2A1O1Ixp33_ASAP7_75t_L g3219 ( 
.A1(n_3131),
.A2(n_549),
.B(n_547),
.C(n_548),
.Y(n_3219)
);

O2A1O1Ixp33_ASAP7_75t_L g3220 ( 
.A1(n_3160),
.A2(n_3165),
.B(n_3159),
.C(n_3123),
.Y(n_3220)
);

NOR2x1_ASAP7_75t_L g3221 ( 
.A(n_3145),
.B(n_550),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_3152),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.Y(n_3222)
);

XOR2xp5_ASAP7_75t_L g3223 ( 
.A(n_3138),
.B(n_551),
.Y(n_3223)
);

OAI211xp5_ASAP7_75t_SL g3224 ( 
.A1(n_3146),
.A2(n_554),
.B(n_552),
.C(n_553),
.Y(n_3224)
);

NAND4xp25_ASAP7_75t_SL g3225 ( 
.A(n_3149),
.B(n_555),
.C(n_553),
.D(n_554),
.Y(n_3225)
);

OAI22xp5_ASAP7_75t_L g3226 ( 
.A1(n_3134),
.A2(n_3140),
.B1(n_3155),
.B2(n_3136),
.Y(n_3226)
);

OAI221xp5_ASAP7_75t_SL g3227 ( 
.A1(n_3121),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.C(n_558),
.Y(n_3227)
);

AND4x1_ASAP7_75t_L g3228 ( 
.A(n_3171),
.B(n_559),
.C(n_556),
.D(n_558),
.Y(n_3228)
);

A2O1A1Ixp33_ASAP7_75t_L g3229 ( 
.A1(n_3126),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_3229)
);

AOI221xp5_ASAP7_75t_L g3230 ( 
.A1(n_3150),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.C(n_563),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3144),
.B(n_562),
.Y(n_3231)
);

NOR2xp33_ASAP7_75t_L g3232 ( 
.A(n_3172),
.B(n_564),
.Y(n_3232)
);

NAND3xp33_ASAP7_75t_SL g3233 ( 
.A(n_3130),
.B(n_564),
.C(n_565),
.Y(n_3233)
);

NOR3xp33_ASAP7_75t_L g3234 ( 
.A(n_3172),
.B(n_567),
.C(n_568),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_3127),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.Y(n_3235)
);

NOR4xp25_ASAP7_75t_L g3236 ( 
.A(n_3125),
.B(n_571),
.C(n_569),
.D(n_570),
.Y(n_3236)
);

OAI22xp33_ASAP7_75t_SL g3237 ( 
.A1(n_3125),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.Y(n_3237)
);

OAI22xp5_ASAP7_75t_L g3238 ( 
.A1(n_3127),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.Y(n_3238)
);

OAI221xp5_ASAP7_75t_L g3239 ( 
.A1(n_3127),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.C(n_577),
.Y(n_3239)
);

NOR2x1p5_ASAP7_75t_L g3240 ( 
.A(n_3202),
.B(n_576),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3223),
.Y(n_3241)
);

AND4x1_ASAP7_75t_L g3242 ( 
.A(n_3195),
.B(n_580),
.C(n_578),
.D(n_579),
.Y(n_3242)
);

OAI22x1_ASAP7_75t_L g3243 ( 
.A1(n_3228),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_3243)
);

OR3x2_ASAP7_75t_L g3244 ( 
.A(n_3199),
.B(n_581),
.C(n_582),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_3182),
.Y(n_3245)
);

AOI22xp5_ASAP7_75t_SL g3246 ( 
.A1(n_3204),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_3182),
.Y(n_3247)
);

XNOR2xp5_ASAP7_75t_L g3248 ( 
.A(n_3203),
.B(n_583),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3212),
.Y(n_3249)
);

NAND2x1p5_ASAP7_75t_L g3250 ( 
.A(n_3213),
.B(n_584),
.Y(n_3250)
);

XNOR2x1_ASAP7_75t_L g3251 ( 
.A(n_3221),
.B(n_584),
.Y(n_3251)
);

AND2x4_ASAP7_75t_L g3252 ( 
.A(n_3218),
.B(n_585),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3236),
.B(n_585),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3212),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3194),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3211),
.Y(n_3256)
);

AND2x4_ASAP7_75t_L g3257 ( 
.A(n_3191),
.B(n_586),
.Y(n_3257)
);

AOI22xp5_ASAP7_75t_L g3258 ( 
.A1(n_3200),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3210),
.Y(n_3259)
);

OAI22x1_ASAP7_75t_L g3260 ( 
.A1(n_3225),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3188),
.B(n_3232),
.Y(n_3261)
);

INVx3_ASAP7_75t_L g3262 ( 
.A(n_3198),
.Y(n_3262)
);

OA22x2_ASAP7_75t_L g3263 ( 
.A1(n_3208),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3231),
.Y(n_3264)
);

HB1xp67_ASAP7_75t_L g3265 ( 
.A(n_3193),
.Y(n_3265)
);

XNOR2x1_ASAP7_75t_L g3266 ( 
.A(n_3226),
.B(n_590),
.Y(n_3266)
);

NOR2xp33_ASAP7_75t_L g3267 ( 
.A(n_3214),
.B(n_591),
.Y(n_3267)
);

HB1xp67_ASAP7_75t_L g3268 ( 
.A(n_3201),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3197),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3206),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_3237),
.B(n_3234),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_3186),
.B(n_592),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3219),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3205),
.Y(n_3274)
);

INVxp67_ASAP7_75t_L g3275 ( 
.A(n_3207),
.Y(n_3275)
);

AOI21x1_ASAP7_75t_L g3276 ( 
.A1(n_3215),
.A2(n_592),
.B(n_593),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3216),
.Y(n_3277)
);

XOR2x1_ASAP7_75t_L g3278 ( 
.A(n_3209),
.B(n_594),
.Y(n_3278)
);

NAND2x1p5_ASAP7_75t_L g3279 ( 
.A(n_3196),
.B(n_3192),
.Y(n_3279)
);

NOR2x1p5_ASAP7_75t_L g3280 ( 
.A(n_3233),
.B(n_595),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_3185),
.B(n_3235),
.Y(n_3281)
);

AND4x1_ASAP7_75t_L g3282 ( 
.A(n_3220),
.B(n_3217),
.C(n_3229),
.D(n_3184),
.Y(n_3282)
);

AND2x4_ASAP7_75t_L g3283 ( 
.A(n_3190),
.B(n_595),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3230),
.B(n_596),
.Y(n_3284)
);

HB1xp67_ASAP7_75t_L g3285 ( 
.A(n_3238),
.Y(n_3285)
);

NOR2x1p5_ASAP7_75t_L g3286 ( 
.A(n_3278),
.B(n_3189),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3244),
.Y(n_3287)
);

NOR3xp33_ASAP7_75t_SL g3288 ( 
.A(n_3267),
.B(n_3239),
.C(n_3224),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3263),
.Y(n_3289)
);

O2A1O1Ixp33_ASAP7_75t_SL g3290 ( 
.A1(n_3253),
.A2(n_3183),
.B(n_3222),
.C(n_3187),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3250),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3252),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3243),
.Y(n_3293)
);

NAND2x1p5_ASAP7_75t_L g3294 ( 
.A(n_3242),
.B(n_3227),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3257),
.Y(n_3295)
);

XNOR2x1_ASAP7_75t_L g3296 ( 
.A(n_3251),
.B(n_596),
.Y(n_3296)
);

HB1xp67_ASAP7_75t_L g3297 ( 
.A(n_3260),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3276),
.Y(n_3298)
);

AOI22xp33_ASAP7_75t_L g3299 ( 
.A1(n_3240),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_3299)
);

AOI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_3259),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_3300)
);

XNOR2x1_ASAP7_75t_L g3301 ( 
.A(n_3266),
.B(n_601),
.Y(n_3301)
);

BUFx2_ASAP7_75t_L g3302 ( 
.A(n_3245),
.Y(n_3302)
);

INVx2_ASAP7_75t_SL g3303 ( 
.A(n_3280),
.Y(n_3303)
);

OR2x6_ASAP7_75t_L g3304 ( 
.A(n_3249),
.B(n_3254),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3271),
.A2(n_601),
.B(n_602),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3246),
.B(n_602),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3247),
.B(n_603),
.Y(n_3307)
);

NAND3xp33_ASAP7_75t_L g3308 ( 
.A(n_3258),
.B(n_603),
.C(n_604),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_3255),
.B(n_604),
.Y(n_3309)
);

XNOR2xp5_ASAP7_75t_L g3310 ( 
.A(n_3248),
.B(n_605),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3262),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3265),
.Y(n_3312)
);

OR3x2_ASAP7_75t_L g3313 ( 
.A(n_3274),
.B(n_605),
.C(n_606),
.Y(n_3313)
);

XNOR2xp5_ASAP7_75t_L g3314 ( 
.A(n_3282),
.B(n_606),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3283),
.Y(n_3315)
);

INVxp67_ASAP7_75t_SL g3316 ( 
.A(n_3261),
.Y(n_3316)
);

INVx3_ASAP7_75t_L g3317 ( 
.A(n_3272),
.Y(n_3317)
);

XOR2xp5_ASAP7_75t_L g3318 ( 
.A(n_3241),
.B(n_607),
.Y(n_3318)
);

NAND3xp33_ASAP7_75t_SL g3319 ( 
.A(n_3284),
.B(n_607),
.C(n_608),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3256),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3268),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3318),
.Y(n_3322)
);

OAI21x1_ASAP7_75t_SL g3323 ( 
.A1(n_3305),
.A2(n_3273),
.B(n_3277),
.Y(n_3323)
);

OAI22x1_ASAP7_75t_L g3324 ( 
.A1(n_3314),
.A2(n_3275),
.B1(n_3279),
.B2(n_3269),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3290),
.A2(n_3285),
.B(n_3270),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3293),
.B(n_3264),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_3294),
.B(n_3281),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3307),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_R g3329 ( 
.A(n_3319),
.B(n_609),
.Y(n_3329)
);

XNOR2xp5_ASAP7_75t_L g3330 ( 
.A(n_3310),
.B(n_609),
.Y(n_3330)
);

OA22x2_ASAP7_75t_L g3331 ( 
.A1(n_3304),
.A2(n_3298),
.B1(n_3312),
.B2(n_3289),
.Y(n_3331)
);

AOI31xp33_ASAP7_75t_L g3332 ( 
.A1(n_3296),
.A2(n_612),
.A3(n_610),
.B(n_611),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3313),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3297),
.B(n_610),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3309),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3306),
.A2(n_611),
.B(n_613),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3299),
.B(n_613),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3301),
.Y(n_3338)
);

OAI22x1_ASAP7_75t_L g3339 ( 
.A1(n_3286),
.A2(n_3302),
.B1(n_3287),
.B2(n_3308),
.Y(n_3339)
);

OAI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3325),
.A2(n_3334),
.B(n_3331),
.Y(n_3340)
);

XOR2xp5_ASAP7_75t_L g3341 ( 
.A(n_3330),
.B(n_3321),
.Y(n_3341)
);

NAND2x1p5_ASAP7_75t_L g3342 ( 
.A(n_3327),
.B(n_3291),
.Y(n_3342)
);

AOI22x1_ASAP7_75t_L g3343 ( 
.A1(n_3339),
.A2(n_3320),
.B1(n_3311),
.B2(n_3316),
.Y(n_3343)
);

HB1xp67_ASAP7_75t_L g3344 ( 
.A(n_3329),
.Y(n_3344)
);

NOR2xp67_ASAP7_75t_L g3345 ( 
.A(n_3336),
.B(n_3300),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3332),
.B(n_3292),
.Y(n_3346)
);

XOR2xp5_ASAP7_75t_L g3347 ( 
.A(n_3324),
.B(n_3295),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3333),
.B(n_3303),
.Y(n_3348)
);

INVx4_ASAP7_75t_L g3349 ( 
.A(n_3326),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3335),
.Y(n_3350)
);

AO22x2_ASAP7_75t_L g3351 ( 
.A1(n_3323),
.A2(n_3315),
.B1(n_3317),
.B2(n_3304),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3322),
.A2(n_3288),
.B1(n_617),
.B2(n_614),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3337),
.B(n_614),
.Y(n_3353)
);

CKINVDCx5p33_ASAP7_75t_R g3354 ( 
.A(n_3349),
.Y(n_3354)
);

INVx2_ASAP7_75t_SL g3355 ( 
.A(n_3342),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3351),
.Y(n_3356)
);

HB1xp67_ASAP7_75t_L g3357 ( 
.A(n_3340),
.Y(n_3357)
);

OAI22xp5_ASAP7_75t_SL g3358 ( 
.A1(n_3347),
.A2(n_3338),
.B1(n_3328),
.B2(n_619),
.Y(n_3358)
);

OAI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3352),
.A2(n_619),
.B1(n_616),
.B2(n_618),
.Y(n_3359)
);

OAI22x1_ASAP7_75t_L g3360 ( 
.A1(n_3343),
.A2(n_620),
.B1(n_616),
.B2(n_618),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3353),
.Y(n_3361)
);

INVx2_ASAP7_75t_SL g3362 ( 
.A(n_3350),
.Y(n_3362)
);

OAI22x1_ASAP7_75t_L g3363 ( 
.A1(n_3341),
.A2(n_3344),
.B1(n_3346),
.B2(n_3348),
.Y(n_3363)
);

XNOR2x1_ASAP7_75t_L g3364 ( 
.A(n_3345),
.B(n_620),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_SL g3365 ( 
.A1(n_3342),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3355),
.A2(n_625),
.B1(n_622),
.B2(n_623),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3364),
.B(n_625),
.Y(n_3367)
);

INVxp33_ASAP7_75t_L g3368 ( 
.A(n_3365),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3356),
.B(n_626),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3360),
.B(n_3357),
.Y(n_3370)
);

BUFx2_ASAP7_75t_L g3371 ( 
.A(n_3354),
.Y(n_3371)
);

AOI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3362),
.A2(n_626),
.B(n_627),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3363),
.A2(n_628),
.B(n_629),
.Y(n_3373)
);

OAI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3358),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3359),
.A2(n_630),
.B(n_631),
.Y(n_3375)
);

OAI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_3361),
.A2(n_631),
.B(n_632),
.Y(n_3376)
);

AOI221xp5_ASAP7_75t_L g3377 ( 
.A1(n_3373),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.C(n_635),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3369),
.A2(n_636),
.B1(n_633),
.B2(n_634),
.Y(n_3378)
);

OAI22xp5_ASAP7_75t_L g3379 ( 
.A1(n_3367),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3370),
.A2(n_637),
.B(n_638),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_3371),
.A2(n_3368),
.B1(n_3375),
.B2(n_3374),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_3372),
.A2(n_640),
.B(n_641),
.Y(n_3382)
);

AOI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3366),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3376),
.A2(n_643),
.B(n_644),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_L g3385 ( 
.A1(n_3381),
.A2(n_643),
.B(n_644),
.Y(n_3385)
);

OAI222xp33_ASAP7_75t_L g3386 ( 
.A1(n_3382),
.A2(n_647),
.B1(n_649),
.B2(n_645),
.C1(n_646),
.C2(n_648),
.Y(n_3386)
);

AOI222xp33_ASAP7_75t_SL g3387 ( 
.A1(n_3379),
.A2(n_647),
.B1(n_649),
.B2(n_645),
.C1(n_646),
.C2(n_648),
.Y(n_3387)
);

AOI222xp33_ASAP7_75t_SL g3388 ( 
.A1(n_3378),
.A2(n_652),
.B1(n_654),
.B2(n_650),
.C1(n_651),
.C2(n_653),
.Y(n_3388)
);

AOI321xp33_ASAP7_75t_L g3389 ( 
.A1(n_3384),
.A2(n_654),
.A3(n_656),
.B1(n_651),
.B2(n_653),
.C(n_655),
.Y(n_3389)
);

AOI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3387),
.A2(n_3377),
.B1(n_3383),
.B2(n_3380),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_SL g3391 ( 
.A1(n_3385),
.A2(n_658),
.B1(n_655),
.B2(n_657),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3391),
.B(n_3388),
.Y(n_3392)
);

AO21x2_ASAP7_75t_L g3393 ( 
.A1(n_3390),
.A2(n_3386),
.B(n_3389),
.Y(n_3393)
);

AOI21xp33_ASAP7_75t_L g3394 ( 
.A1(n_3393),
.A2(n_657),
.B(n_658),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3394),
.A2(n_3392),
.B1(n_661),
.B2(n_659),
.Y(n_3395)
);


endmodule