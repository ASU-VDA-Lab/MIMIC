module fake_jpeg_29775_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_55),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_42),
.B1(n_35),
.B2(n_38),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_68),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_38),
.B1(n_47),
.B2(n_36),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_48),
.B1(n_39),
.B2(n_45),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_39),
.CI(n_43),
.CON(n_71),
.SN(n_71)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_3),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_81),
.Y(n_86)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_16),
.B1(n_34),
.B2(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_83),
.Y(n_92)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_20),
.B1(n_24),
.B2(n_9),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_4),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_5),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_17),
.A3(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_93),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_15),
.C(n_26),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_96),
.B(n_14),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_19),
.B(n_23),
.C(n_11),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_87),
.C(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_106),
.B1(n_94),
.B2(n_21),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_91),
.B1(n_96),
.B2(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_113),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_109),
.Y(n_117)
);

INVxp33_ASAP7_75t_SL g116 ( 
.A(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_118),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_112),
.B(n_110),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_114),
.C(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_107),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_106),
.B(n_101),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_124),
.Y(n_125)
);


endmodule