module fake_netlist_1_2184_n_14 (n_3, n_1, n_2, n_0, n_14);
input n_3;
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_3), .B(n_2), .Y(n_4) );
INVx3_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
NAND3xp33_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .C(n_1), .Y(n_7) );
OR2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_5), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
OAI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_7), .B1(n_4), .B2(n_2), .Y(n_10) );
NOR4xp75_ASAP7_75t_SL g11 ( .A(n_10), .B(n_0), .C(n_1), .D(n_2), .Y(n_11) );
OR2x2_ASAP7_75t_L g12 ( .A(n_10), .B(n_9), .Y(n_12) );
BUFx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_11), .B1(n_1), .B2(n_3), .Y(n_14) );
endmodule