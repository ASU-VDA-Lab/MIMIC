module fake_jpeg_1056_n_471 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_51),
.B(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_8),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_54),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_21),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_56),
.A2(n_78),
.B1(n_27),
.B2(n_34),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_67),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_16),
.B(n_8),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_35),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_30),
.B(n_7),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_83),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12f_ASAP7_75t_SL g136 ( 
.A(n_84),
.Y(n_136)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_93),
.Y(n_129)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_36),
.B(n_6),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_100),
.Y(n_152)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_103),
.Y(n_109)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_36),
.B(n_6),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_101),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_18),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_64),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_106),
.B(n_155),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_50),
.B1(n_49),
.B2(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_108),
.A2(n_112),
.B1(n_146),
.B2(n_151),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_62),
.A2(n_50),
.B1(n_49),
.B2(n_43),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_50),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_116),
.A2(n_134),
.B1(n_84),
.B2(n_26),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_50),
.C(n_49),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_23),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_139),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_56),
.A2(n_55),
.B1(n_43),
.B2(n_49),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_70),
.B(n_23),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_57),
.A2(n_43),
.B1(n_40),
.B2(n_29),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_58),
.B1(n_101),
.B2(n_61),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_40),
.B1(n_29),
.B2(n_34),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_76),
.B(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_159),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_40),
.B1(n_29),
.B2(n_27),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_75),
.A2(n_29),
.B1(n_40),
.B2(n_39),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_89),
.B1(n_84),
.B2(n_93),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_65),
.B(n_22),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_76),
.B(n_22),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_163),
.B(n_179),
.Y(n_231)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_32),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_165),
.B(n_186),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_42),
.B1(n_17),
.B2(n_122),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_166),
.A2(n_183),
.B1(n_185),
.B2(n_112),
.Y(n_238)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_167),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_168),
.A2(n_197),
.B1(n_157),
.B2(n_142),
.Y(n_245)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

CKINVDCx6p67_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_182),
.A2(n_116),
.B1(n_150),
.B2(n_119),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_17),
.B1(n_96),
.B2(n_94),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_123),
.B(n_37),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_192),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_134),
.A2(n_59),
.B1(n_90),
.B2(n_83),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_105),
.B(n_32),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_130),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_87),
.B1(n_66),
.B2(n_74),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_104),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_129),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_204),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_107),
.B(n_39),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_206),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_117),
.B(n_26),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_116),
.Y(n_239)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_147),
.B(n_37),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_SL g271 ( 
.A1(n_218),
.A2(n_136),
.B(n_205),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_121),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_130),
.C(n_114),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_165),
.B(n_116),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_169),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_153),
.B1(n_128),
.B2(n_156),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_245),
.B1(n_234),
.B2(n_175),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_129),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_236),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_173),
.A2(n_194),
.B1(n_188),
.B2(n_196),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_173),
.B1(n_197),
.B2(n_182),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_175),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_147),
.Y(n_270)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_253),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_261),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_212),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_254),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_173),
.B1(n_168),
.B2(n_180),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_252),
.B1(n_258),
.B2(n_214),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_177),
.B1(n_157),
.B2(n_202),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_210),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_264),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_259),
.B1(n_249),
.B2(n_251),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_257),
.B(n_268),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_181),
.B1(n_162),
.B2(n_203),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_232),
.A2(n_146),
.B1(n_151),
.B2(n_154),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_219),
.C(n_227),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_228),
.C(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_234),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_269),
.Y(n_288)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_175),
.B(n_170),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_136),
.B(n_228),
.Y(n_289)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_271),
.B1(n_276),
.B2(n_150),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_223),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_223),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_133),
.C(n_148),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_277),
.C(n_171),
.Y(n_302)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_153),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_243),
.B(n_230),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_278),
.A2(n_287),
.B(n_305),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_281),
.A2(n_303),
.B1(n_208),
.B2(n_162),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_284),
.A2(n_289),
.B(n_298),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_291),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_256),
.B(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_246),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_211),
.B1(n_213),
.B2(n_176),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_263),
.B1(n_222),
.B2(n_240),
.Y(n_316)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_235),
.C(n_233),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_296),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_256),
.A2(n_229),
.B(n_221),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_244),
.B(n_253),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_247),
.B(n_230),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_272),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_193),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_252),
.A2(n_211),
.B1(n_187),
.B2(n_164),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_257),
.A2(n_216),
.B1(n_244),
.B2(n_222),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_258),
.B1(n_267),
.B2(n_269),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_229),
.B(n_221),
.C(n_224),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_288),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_323),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_308),
.A2(n_318),
.B1(n_321),
.B2(n_303),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_260),
.B1(n_274),
.B2(n_277),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_309),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_248),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_310),
.B(n_326),
.C(n_279),
.Y(n_355)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_313),
.A2(n_332),
.B(n_305),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_280),
.A2(n_276),
.B1(n_275),
.B2(n_226),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_226),
.B1(n_240),
.B2(n_222),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_280),
.A2(n_201),
.B1(n_198),
.B2(n_178),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_235),
.Y(n_319)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_319),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_331),
.C(n_302),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_220),
.B1(n_118),
.B2(n_195),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_220),
.Y(n_324)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_281),
.A2(n_224),
.B1(n_119),
.B2(n_167),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_328),
.B1(n_304),
.B2(n_287),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_172),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_288),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_297),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_128),
.C(n_161),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_206),
.B(n_174),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_353),
.B1(n_313),
.B2(n_332),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_283),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_340),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_319),
.B(n_286),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_336),
.B(n_348),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_310),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_349),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_342),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_285),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_285),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_291),
.C(n_301),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_347),
.C(n_350),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_344),
.A2(n_328),
.B1(n_325),
.B2(n_317),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_301),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_359),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_289),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_307),
.B(n_293),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_331),
.B(n_292),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_297),
.C(n_293),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_312),
.B(n_290),
.Y(n_351)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_312),
.A2(n_297),
.B1(n_292),
.B2(n_279),
.Y(n_353)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_306),
.B(n_294),
.C(n_191),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_329),
.C(n_332),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_358),
.A2(n_313),
.B(n_330),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_142),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_346),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_362),
.B(n_378),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_341),
.A2(n_329),
.B1(n_328),
.B2(n_323),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_363),
.A2(n_98),
.B1(n_77),
.B2(n_103),
.Y(n_399)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_324),
.Y(n_366)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_381),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_327),
.C(n_315),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_334),
.C(n_350),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_372),
.A2(n_156),
.B1(n_150),
.B2(n_118),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_358),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_376),
.A2(n_379),
.B1(n_344),
.B2(n_359),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_333),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_341),
.A2(n_308),
.B1(n_318),
.B2(n_316),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_325),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_321),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_383),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_386),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_340),
.C(n_347),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_393),
.C(n_365),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_392),
.A2(n_396),
.B1(n_402),
.B2(n_381),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_342),
.C(n_125),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_368),
.A2(n_363),
.B1(n_360),
.B2(n_367),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_394),
.A2(n_399),
.B1(n_372),
.B2(n_374),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_366),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_370),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_379),
.A2(n_33),
.B1(n_28),
.B2(n_143),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_365),
.B(n_65),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_380),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_412),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_401),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_410),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_417),
.B1(n_398),
.B2(n_388),
.Y(n_421)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_369),
.C(n_361),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_396),
.B1(n_388),
.B2(n_403),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_361),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_414),
.C(n_415),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_383),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_377),
.C(n_371),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_377),
.C(n_364),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_419),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_386),
.A2(n_125),
.B(n_33),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_28),
.Y(n_419)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

AOI211xp5_ASAP7_75t_L g422 ( 
.A1(n_418),
.A2(n_398),
.B(n_397),
.C(n_400),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_L g435 ( 
.A1(n_422),
.A2(n_413),
.B(n_404),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_406),
.A2(n_397),
.B1(n_400),
.B2(n_399),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_429),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_428),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_409),
.A2(n_143),
.B(n_11),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_415),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_10),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_430),
.A2(n_433),
.B(n_11),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_410),
.A2(n_31),
.B1(n_41),
.B2(n_10),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_434),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_10),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_435),
.A2(n_441),
.B(n_428),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_414),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_440),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_442),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_412),
.C(n_41),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_424),
.A2(n_31),
.B(n_41),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_31),
.B(n_41),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_434),
.C(n_425),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_446),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_6),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_436),
.A2(n_426),
.B(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_448),
.B(n_443),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_444),
.B(n_426),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_452),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_443),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_439),
.A2(n_422),
.B1(n_430),
.B2(n_433),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_5),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_453),
.B(n_455),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_5),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_451),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_456),
.A2(n_458),
.B(n_459),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_445),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_460),
.A2(n_447),
.B(n_11),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_450),
.C(n_440),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_462),
.A2(n_463),
.B(n_464),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_457),
.A2(n_12),
.B(n_14),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_14),
.C(n_12),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_466),
.A2(n_0),
.B(n_2),
.Y(n_468)
);

HAxp5_ASAP7_75t_SL g469 ( 
.A(n_468),
.B(n_4),
.CON(n_469),
.SN(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_467),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_470),
.Y(n_471)
);


endmodule