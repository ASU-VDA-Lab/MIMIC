module real_aes_16338_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1994;
wire n_1225;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1583;
wire n_1095;
wire n_1987;
wire n_859;
wire n_1465;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1632;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_1940;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_1648;
wire n_724;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1973;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1812;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_1971;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1691;
wire n_640;
wire n_1721;
wire n_1176;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_1280;
wire n_1369;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g814 ( .A(n_0), .Y(n_814) );
OAI211xp5_ASAP7_75t_L g1389 ( .A1(n_1), .A2(n_477), .B(n_1386), .C(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1), .Y(n_1403) );
INVx1_ASAP7_75t_L g1644 ( .A(n_2), .Y(n_1644) );
OAI22xp33_ASAP7_75t_L g1656 ( .A1(n_2), .A2(n_370), .B1(n_705), .B2(n_934), .Y(n_1656) );
AOI221xp5_ASAP7_75t_L g1639 ( .A1(n_3), .A2(n_194), .B1(n_591), .B2(n_596), .C(n_1640), .Y(n_1639) );
AOI222xp33_ASAP7_75t_L g1664 ( .A1(n_3), .A2(n_125), .B1(n_337), .B2(n_568), .C1(n_672), .C2(n_881), .Y(n_1664) );
INVx1_ASAP7_75t_L g389 ( .A(n_4), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_4), .B(n_399), .Y(n_513) );
AND2x2_ASAP7_75t_L g588 ( .A(n_4), .B(n_437), .Y(n_588) );
AND2x2_ASAP7_75t_L g605 ( .A(n_4), .B(n_282), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g840 ( .A1(n_5), .A2(n_415), .B(n_538), .C(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g855 ( .A(n_5), .Y(n_855) );
INVx1_ASAP7_75t_L g888 ( .A(n_6), .Y(n_888) );
INVx1_ASAP7_75t_L g1260 ( .A(n_7), .Y(n_1260) );
INVx1_ASAP7_75t_L g1964 ( .A(n_8), .Y(n_1964) );
INVx1_ASAP7_75t_L g1506 ( .A(n_9), .Y(n_1506) );
AOI22xp5_ASAP7_75t_L g1730 ( .A1(n_10), .A2(n_71), .B1(n_1681), .B2(n_1685), .Y(n_1730) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_11), .A2(n_84), .B1(n_671), .B2(n_1258), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1275 ( .A1(n_11), .A2(n_18), .B1(n_954), .B2(n_1276), .C(n_1278), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_12), .A2(n_26), .B1(n_1122), .B2(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1191 ( .A(n_12), .Y(n_1191) );
INVx1_ASAP7_75t_L g1987 ( .A(n_13), .Y(n_1987) );
OAI211xp5_ASAP7_75t_L g1992 ( .A1(n_13), .A2(n_477), .B(n_1608), .C(n_1993), .Y(n_1992) );
INVx1_ASAP7_75t_L g1422 ( .A(n_14), .Y(n_1422) );
INVx1_ASAP7_75t_L g1307 ( .A(n_15), .Y(n_1307) );
INVx1_ASAP7_75t_L g1563 ( .A(n_16), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_17), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g1267 ( .A1(n_18), .A2(n_266), .B1(n_672), .B2(n_1155), .Y(n_1267) );
INVx1_ASAP7_75t_L g1967 ( .A(n_19), .Y(n_1967) );
INVx2_ASAP7_75t_L g465 ( .A(n_20), .Y(n_465) );
OAI22xp33_ASAP7_75t_L g1533 ( .A1(n_21), .A2(n_255), .B1(n_496), .B2(n_794), .Y(n_1533) );
OAI22xp5_ASAP7_75t_L g1540 ( .A1(n_21), .A2(n_255), .B1(n_913), .B2(n_1010), .Y(n_1540) );
INVx1_ASAP7_75t_L g651 ( .A(n_22), .Y(n_651) );
INVx1_ASAP7_75t_L g819 ( .A(n_23), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_24), .A2(n_248), .B1(n_490), .B2(n_1527), .Y(n_1526) );
OAI22xp33_ASAP7_75t_L g1535 ( .A1(n_24), .A2(n_248), .B1(n_1008), .B2(n_1536), .Y(n_1535) );
AOI221xp5_ASAP7_75t_L g1556 ( .A1(n_25), .A2(n_240), .B1(n_967), .B2(n_1078), .C(n_1217), .Y(n_1556) );
INVxp67_ASAP7_75t_SL g1567 ( .A(n_25), .Y(n_1567) );
AOI221xp5_ASAP7_75t_L g1170 ( .A1(n_26), .A2(n_46), .B1(n_1171), .B2(n_1173), .C(n_1174), .Y(n_1170) );
INVx1_ASAP7_75t_L g1264 ( .A(n_27), .Y(n_1264) );
INVx1_ASAP7_75t_L g1670 ( .A(n_28), .Y(n_1670) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_29), .A2(n_316), .B1(n_457), .B2(n_794), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_29), .A2(n_346), .B1(n_433), .B2(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g1712 ( .A1(n_30), .A2(n_245), .B1(n_1688), .B2(n_1691), .Y(n_1712) );
INVx1_ASAP7_75t_L g1973 ( .A(n_31), .Y(n_1973) );
OA222x2_ASAP7_75t_L g1066 ( .A1(n_32), .A2(n_91), .B1(n_276), .B2(n_1067), .C1(n_1069), .C2(n_1073), .Y(n_1066) );
INVx1_ASAP7_75t_L g1120 ( .A(n_32), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_33), .Y(n_384) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_33), .B(n_382), .Y(n_1682) );
AOI22xp5_ASAP7_75t_L g1729 ( .A1(n_34), .A2(n_222), .B1(n_1688), .B2(n_1691), .Y(n_1729) );
INVx1_ASAP7_75t_L g1589 ( .A(n_35), .Y(n_1589) );
XNOR2xp5_ASAP7_75t_L g1634 ( .A(n_36), .B(n_1635), .Y(n_1634) );
INVx1_ASAP7_75t_L g1482 ( .A(n_37), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_38), .A2(n_350), .B1(n_586), .B2(n_955), .Y(n_1213) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_38), .Y(n_1230) );
INVx1_ASAP7_75t_L g1903 ( .A(n_39), .Y(n_1903) );
OAI211xp5_ASAP7_75t_L g1912 ( .A1(n_39), .A2(n_615), .B(n_1913), .C(n_1919), .Y(n_1912) );
AOI221xp5_ASAP7_75t_L g1548 ( .A1(n_40), .A2(n_110), .B1(n_596), .B2(n_1078), .C(n_1549), .Y(n_1548) );
AOI22xp33_ASAP7_75t_L g1577 ( .A1(n_40), .A2(n_117), .B1(n_1232), .B2(n_1578), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_41), .A2(n_241), .B1(n_674), .B2(n_985), .Y(n_1156) );
INVx1_ASAP7_75t_L g1176 ( .A(n_41), .Y(n_1176) );
AOI22xp5_ASAP7_75t_L g1704 ( .A1(n_42), .A2(n_307), .B1(n_1688), .B2(n_1691), .Y(n_1704) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_43), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_44), .A2(n_302), .B1(n_1008), .B2(n_1310), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_44), .A2(n_201), .B1(n_457), .B2(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1015 ( .A(n_45), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g1160 ( .A1(n_46), .A2(n_342), .B1(n_688), .B2(n_1155), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1927 ( .A1(n_47), .A2(n_333), .B1(n_591), .B2(n_634), .C(n_1640), .Y(n_1927) );
INVxp67_ASAP7_75t_SL g1935 ( .A(n_47), .Y(n_1935) );
INVxp67_ASAP7_75t_SL g1263 ( .A(n_48), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_48), .A2(n_191), .B1(n_627), .B2(n_1284), .Y(n_1283) );
AOI22xp5_ASAP7_75t_L g1722 ( .A1(n_49), .A2(n_132), .B1(n_1688), .B2(n_1691), .Y(n_1722) );
INVx1_ASAP7_75t_L g1532 ( .A(n_50), .Y(n_1532) );
OAI211xp5_ASAP7_75t_L g1537 ( .A1(n_50), .A2(n_415), .B(n_895), .C(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1909 ( .A(n_51), .Y(n_1909) );
OAI22xp5_ASAP7_75t_L g1928 ( .A1(n_51), .A2(n_237), .B1(n_1637), .B2(n_1929), .Y(n_1928) );
AOI22xp33_ASAP7_75t_SL g1321 ( .A1(n_52), .A2(n_147), .B1(n_1322), .B2(n_1323), .Y(n_1321) );
AOI22xp33_ASAP7_75t_SL g1350 ( .A1(n_52), .A2(n_281), .B1(n_1232), .B2(n_1345), .Y(n_1350) );
INVx1_ASAP7_75t_L g1022 ( .A(n_53), .Y(n_1022) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_54), .A2(n_411), .B(n_415), .C(n_420), .Y(n_410) );
INVx1_ASAP7_75t_L g486 ( .A(n_54), .Y(n_486) );
INVx1_ASAP7_75t_L g1418 ( .A(n_55), .Y(n_1418) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_56), .Y(n_1090) );
INVx1_ASAP7_75t_L g1271 ( .A(n_57), .Y(n_1271) );
INVx1_ASAP7_75t_L g1559 ( .A(n_58), .Y(n_1559) );
INVx1_ASAP7_75t_L g882 ( .A(n_59), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g1720 ( .A1(n_60), .A2(n_193), .B1(n_1681), .B2(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g1562 ( .A(n_61), .Y(n_1562) );
OAI322xp33_ASAP7_75t_L g1565 ( .A1(n_61), .A2(n_570), .A3(n_867), .B1(n_937), .B2(n_1566), .C1(n_1569), .C2(n_1574), .Y(n_1565) );
AOI22xp33_ASAP7_75t_SL g1218 ( .A1(n_62), .A2(n_289), .B1(n_955), .B2(n_1219), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_62), .A2(n_272), .B1(n_1111), .B2(n_1232), .Y(n_1231) );
INVxp67_ASAP7_75t_SL g1926 ( .A(n_63), .Y(n_1926) );
AOI22xp33_ASAP7_75t_L g1945 ( .A1(n_63), .A2(n_162), .B1(n_1258), .B2(n_1946), .Y(n_1945) );
CKINVDCx5p33_ASAP7_75t_R g1262 ( .A(n_64), .Y(n_1262) );
INVx1_ASAP7_75t_L g1293 ( .A(n_65), .Y(n_1293) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_66), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_67), .A2(n_81), .B1(n_683), .B2(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1175 ( .A(n_67), .Y(n_1175) );
INVx1_ASAP7_75t_L g525 ( .A(n_68), .Y(n_525) );
OAI22xp33_ASAP7_75t_SL g1209 ( .A1(n_69), .A2(n_278), .B1(n_536), .B2(n_1089), .Y(n_1209) );
INVx1_ASAP7_75t_L g1246 ( .A(n_69), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_70), .A2(n_120), .B1(n_598), .B2(n_602), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_70), .A2(n_260), .B1(n_674), .B2(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g1486 ( .A(n_72), .Y(n_1486) );
INVx1_ASAP7_75t_L g1617 ( .A(n_73), .Y(n_1617) );
AOI21xp33_ASAP7_75t_L g966 ( .A1(n_74), .A2(n_967), .B(n_968), .Y(n_966) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_74), .A2(n_296), .B1(n_985), .B2(n_990), .C(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g1596 ( .A(n_75), .Y(n_1596) );
INVx1_ASAP7_75t_L g1597 ( .A(n_76), .Y(n_1597) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_77), .Y(n_1147) );
XOR2x2_ASAP7_75t_L g580 ( .A(n_78), .B(n_581), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_79), .A2(n_137), .B1(n_391), .B2(n_768), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_79), .A2(n_137), .B1(n_457), .B2(n_786), .Y(n_785) );
OAI222xp33_ASAP7_75t_L g928 ( .A1(n_80), .A2(n_89), .B1(n_96), .B2(n_657), .C1(n_929), .C2(n_935), .Y(n_928) );
INVx1_ASAP7_75t_L g1195 ( .A(n_81), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1680 ( .A1(n_82), .A2(n_269), .B1(n_1681), .B2(n_1685), .Y(n_1680) );
INVx1_ASAP7_75t_L g1443 ( .A(n_83), .Y(n_1443) );
OAI211xp5_ASAP7_75t_L g1449 ( .A1(n_83), .A2(n_988), .B(n_1049), .C(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1292 ( .A(n_84), .Y(n_1292) );
INVx1_ASAP7_75t_L g885 ( .A(n_85), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g1009 ( .A1(n_86), .A2(n_90), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_86), .A2(n_90), .B1(n_496), .B2(n_1056), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_87), .Y(n_947) );
INVx1_ASAP7_75t_L g1417 ( .A(n_88), .Y(n_1417) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_91), .A2(n_214), .B1(n_1105), .B2(n_1107), .C(n_1109), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_92), .A2(n_326), .B1(n_441), .B2(n_627), .Y(n_1184) );
INVx1_ASAP7_75t_L g1197 ( .A(n_92), .Y(n_1197) );
INVx1_ASAP7_75t_L g1080 ( .A(n_93), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_93), .A2(n_159), .B1(n_677), .B2(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1031 ( .A(n_94), .Y(n_1031) );
XOR2x2_ASAP7_75t_L g1458 ( .A(n_95), .B(n_1459), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_96), .A2(n_369), .B1(n_979), .B2(n_981), .Y(n_978) );
OR2x2_ASAP7_75t_L g1907 ( .A(n_97), .B(n_643), .Y(n_1907) );
INVx1_ASAP7_75t_L g1517 ( .A(n_98), .Y(n_1517) );
OAI211xp5_ASAP7_75t_L g1529 ( .A1(n_99), .A2(n_477), .B(n_1386), .C(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1539 ( .A(n_99), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g1700 ( .A1(n_100), .A2(n_196), .B1(n_1681), .B2(n_1688), .Y(n_1700) );
OAI221xp5_ASAP7_75t_L g1920 ( .A1(n_101), .A2(n_233), .B1(n_1921), .B2(n_1923), .C(n_1924), .Y(n_1920) );
OAI322xp33_ASAP7_75t_L g1933 ( .A1(n_101), .A2(n_805), .A3(n_1934), .B1(n_1937), .B2(n_1941), .C1(n_1943), .C2(n_1947), .Y(n_1933) );
INVx1_ASAP7_75t_L g1513 ( .A(n_102), .Y(n_1513) );
INVx1_ASAP7_75t_L g807 ( .A(n_103), .Y(n_807) );
INVx1_ASAP7_75t_L g842 ( .A(n_104), .Y(n_842) );
INVx1_ASAP7_75t_L g1463 ( .A(n_105), .Y(n_1463) );
XOR2x2_ASAP7_75t_L g863 ( .A(n_106), .B(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1699 ( .A1(n_106), .A2(n_325), .B1(n_1685), .B2(n_1691), .Y(n_1699) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_107), .A2(n_183), .B1(n_970), .B2(n_971), .Y(n_969) );
INVx1_ASAP7_75t_L g987 ( .A(n_107), .Y(n_987) );
XNOR2xp5_ASAP7_75t_L g1408 ( .A(n_108), .B(n_1409), .Y(n_1408) );
AOI22xp5_ASAP7_75t_L g1706 ( .A1(n_108), .A2(n_182), .B1(n_1681), .B2(n_1707), .Y(n_1706) );
CKINVDCx5p33_ASAP7_75t_R g1270 ( .A(n_109), .Y(n_1270) );
INVx1_ASAP7_75t_L g1573 ( .A(n_110), .Y(n_1573) );
INVx1_ASAP7_75t_L g1531 ( .A(n_111), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_112), .A2(n_347), .B1(n_675), .B2(n_1158), .Y(n_1266) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_112), .A2(n_235), .B1(n_955), .B2(n_1173), .C(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1925 ( .A(n_113), .Y(n_1925) );
AOI22xp33_ASAP7_75t_L g1687 ( .A1(n_114), .A2(n_358), .B1(n_1688), .B2(n_1691), .Y(n_1687) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_115), .A2(n_181), .B1(n_459), .B2(n_786), .Y(n_1388) );
OAI22xp33_ASAP7_75t_L g1398 ( .A1(n_115), .A2(n_181), .B1(n_391), .B2(n_445), .Y(n_1398) );
INVx1_ASAP7_75t_L g1199 ( .A(n_116), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_117), .A2(n_363), .B1(n_1173), .B2(n_1558), .Y(n_1557) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_118), .A2(n_172), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_118), .A2(n_172), .B1(n_850), .B2(n_1046), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1982 ( .A1(n_119), .A2(n_124), .B1(n_768), .B2(n_847), .Y(n_1982) );
OAI22xp33_ASAP7_75t_L g1990 ( .A1(n_119), .A2(n_124), .B1(n_1046), .B2(n_1448), .Y(n_1990) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_120), .A2(n_145), .B1(n_680), .B2(n_683), .Y(n_679) );
INVx1_ASAP7_75t_L g1365 ( .A(n_121), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g1648 ( .A(n_122), .Y(n_1648) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_122), .A2(n_194), .B1(n_1113), .B2(n_1155), .Y(n_1668) );
INVx1_ASAP7_75t_L g382 ( .A(n_123), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g1641 ( .A1(n_125), .A2(n_341), .B1(n_1339), .B2(n_1558), .Y(n_1641) );
OAI22xp5_ASAP7_75t_L g1602 ( .A1(n_126), .A2(n_340), .B1(n_1007), .B2(n_1008), .Y(n_1602) );
OAI22xp5_ASAP7_75t_L g1632 ( .A1(n_126), .A2(n_340), .B1(n_786), .B2(n_1527), .Y(n_1632) );
INVx1_ASAP7_75t_L g1599 ( .A(n_127), .Y(n_1599) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_128), .A2(n_190), .B1(n_653), .B2(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g870 ( .A(n_129), .Y(n_870) );
OAI211xp5_ASAP7_75t_L g1461 ( .A1(n_130), .A2(n_415), .B(n_756), .C(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1471 ( .A(n_130), .Y(n_1471) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_131), .A2(n_372), .B1(n_433), .B2(n_438), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_131), .A2(n_144), .B1(n_457), .B2(n_466), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g1444 ( .A1(n_133), .A2(n_180), .B1(n_1405), .B2(n_1406), .Y(n_1444) );
OAI22xp33_ASAP7_75t_L g1453 ( .A1(n_133), .A2(n_180), .B1(n_1394), .B2(n_1454), .Y(n_1453) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_134), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_134), .A2(n_308), .B1(n_671), .B2(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_135), .A2(n_176), .B1(n_1081), .B2(n_1082), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g1250 ( .A(n_135), .B(n_466), .Y(n_1250) );
INVx1_ASAP7_75t_L g825 ( .A(n_136), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_138), .Y(n_1166) );
INVx1_ASAP7_75t_L g821 ( .A(n_139), .Y(n_821) );
INVx1_ASAP7_75t_L g1377 ( .A(n_140), .Y(n_1377) );
INVx1_ASAP7_75t_L g823 ( .A(n_141), .Y(n_823) );
OAI211xp5_ASAP7_75t_SL g1636 ( .A1(n_142), .A2(n_1637), .B(n_1638), .C(n_1642), .Y(n_1636) );
OAI22xp5_ASAP7_75t_L g1654 ( .A1(n_142), .A2(n_362), .B1(n_657), .B2(n_1655), .Y(n_1654) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_143), .A2(n_155), .B1(n_435), .B2(n_438), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_143), .A2(n_155), .B1(n_794), .B2(n_857), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_144), .A2(n_345), .B1(n_391), .B2(n_445), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_145), .A2(n_260), .B1(n_594), .B2(n_632), .C(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g1489 ( .A(n_146), .Y(n_1489) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_147), .A2(n_262), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
CKINVDCx20_ASAP7_75t_R g1647 ( .A(n_148), .Y(n_1647) );
OAI22xp5_ASAP7_75t_L g1988 ( .A1(n_149), .A2(n_320), .B1(n_438), .B2(n_1405), .Y(n_1988) );
OAI22xp5_ASAP7_75t_L g1991 ( .A1(n_149), .A2(n_320), .B1(n_1056), .B2(n_1394), .Y(n_1991) );
INVx1_ASAP7_75t_L g1986 ( .A(n_150), .Y(n_1986) );
INVx1_ASAP7_75t_L g844 ( .A(n_151), .Y(n_844) );
OAI211xp5_ASAP7_75t_L g851 ( .A1(n_151), .A2(n_477), .B(n_852), .C(n_854), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_152), .A2(n_346), .B1(n_490), .B2(n_496), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_152), .A2(n_316), .B1(n_391), .B2(n_768), .Y(n_911) );
INVx1_ASAP7_75t_L g810 ( .A(n_153), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g1703 ( .A1(n_154), .A2(n_239), .B1(n_1681), .B2(n_1685), .Y(n_1703) );
INVx1_ASAP7_75t_L g1512 ( .A(n_156), .Y(n_1512) );
INVx1_ASAP7_75t_L g1442 ( .A(n_157), .Y(n_1442) );
INVx1_ASAP7_75t_L g1601 ( .A(n_158), .Y(n_1601) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_159), .A2(n_197), .B1(n_598), .B2(n_602), .Y(n_1091) );
INVx1_ASAP7_75t_L g1413 ( .A(n_160), .Y(n_1413) );
INVxp67_ASAP7_75t_SL g1606 ( .A(n_161), .Y(n_1606) );
AOI22xp33_ASAP7_75t_L g1621 ( .A1(n_161), .A2(n_309), .B1(n_1558), .B2(n_1622), .Y(n_1621) );
AOI221xp5_ASAP7_75t_L g1917 ( .A1(n_162), .A2(n_247), .B1(n_1640), .B2(n_1650), .C(n_1918), .Y(n_1917) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_163), .A2(n_308), .B1(n_591), .B2(n_592), .C(n_596), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_163), .A2(n_263), .B1(n_669), .B2(n_672), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_164), .A2(n_357), .B1(n_1405), .B2(n_1406), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1468 ( .A1(n_164), .A2(n_357), .B1(n_466), .B2(n_857), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_165), .A2(n_214), .B1(n_654), .B2(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1121 ( .A(n_165), .Y(n_1121) );
INVx1_ASAP7_75t_L g1367 ( .A(n_166), .Y(n_1367) );
INVx1_ASAP7_75t_L g1369 ( .A(n_167), .Y(n_1369) );
OAI211xp5_ASAP7_75t_L g769 ( .A1(n_168), .A2(n_415), .B(n_770), .C(n_774), .Y(n_769) );
INVx1_ASAP7_75t_L g792 ( .A(n_168), .Y(n_792) );
OAI22xp33_ASAP7_75t_L g1466 ( .A1(n_169), .A2(n_203), .B1(n_768), .B2(n_847), .Y(n_1466) );
OAI22xp33_ASAP7_75t_L g1472 ( .A1(n_169), .A2(n_203), .B1(n_459), .B2(n_1448), .Y(n_1472) );
OAI22xp33_ASAP7_75t_L g846 ( .A1(n_170), .A2(n_273), .B1(n_445), .B2(n_847), .Y(n_846) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_170), .A2(n_273), .B1(n_459), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g1025 ( .A(n_171), .Y(n_1025) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_173), .A2(n_352), .B1(n_756), .B2(n_1223), .C(n_1225), .Y(n_1222) );
INVx1_ASAP7_75t_L g1243 ( .A(n_173), .Y(n_1243) );
INVx1_ASAP7_75t_L g1211 ( .A(n_174), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_174), .A2(n_289), .B1(n_1111), .B2(n_1237), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g1215 ( .A(n_175), .Y(n_1215) );
INVx1_ASAP7_75t_L g1245 ( .A(n_176), .Y(n_1245) );
INVx1_ASAP7_75t_L g1306 ( .A(n_177), .Y(n_1306) );
OAI211xp5_ASAP7_75t_L g1315 ( .A1(n_177), .A2(n_470), .B(n_1049), .C(n_1316), .Y(n_1315) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_178), .A2(n_470), .B(n_477), .C(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g920 ( .A(n_178), .Y(n_920) );
INVx1_ASAP7_75t_L g1970 ( .A(n_179), .Y(n_1970) );
INVxp67_ASAP7_75t_SL g993 ( .A(n_183), .Y(n_993) );
INVx1_ASAP7_75t_L g1391 ( .A(n_184), .Y(n_1391) );
INVx1_ASAP7_75t_L g1615 ( .A(n_185), .Y(n_1615) );
OAI211xp5_ASAP7_75t_L g1983 ( .A1(n_186), .A2(n_532), .B(n_1984), .C(n_1985), .Y(n_1983) );
INVx1_ASAP7_75t_L g1994 ( .A(n_186), .Y(n_1994) );
INVx1_ASAP7_75t_L g1425 ( .A(n_187), .Y(n_1425) );
INVx1_ASAP7_75t_L g1372 ( .A(n_188), .Y(n_1372) );
AOI221xp5_ASAP7_75t_L g1649 ( .A1(n_189), .A2(n_337), .B1(n_967), .B2(n_1217), .C(n_1650), .Y(n_1649) );
INVxp67_ASAP7_75t_SL g1666 ( .A(n_189), .Y(n_1666) );
OAI211xp5_ASAP7_75t_L g583 ( .A1(n_190), .A2(n_584), .B(n_589), .C(n_606), .Y(n_583) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_191), .Y(n_1273) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_192), .Y(n_1088) );
INVx1_ASAP7_75t_L g1202 ( .A(n_193), .Y(n_1202) );
INVx1_ASAP7_75t_L g519 ( .A(n_195), .Y(n_519) );
INVx1_ASAP7_75t_L g1134 ( .A(n_197), .Y(n_1134) );
INVx1_ASAP7_75t_L g421 ( .A(n_198), .Y(n_421) );
INVx1_ASAP7_75t_L g1424 ( .A(n_199), .Y(n_1424) );
INVx1_ASAP7_75t_L g1485 ( .A(n_200), .Y(n_1485) );
INVx1_ASAP7_75t_L g1304 ( .A(n_201), .Y(n_1304) );
INVx1_ASAP7_75t_L g1464 ( .A(n_202), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1469 ( .A1(n_202), .A2(n_477), .B(n_852), .C(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g965 ( .A(n_204), .Y(n_965) );
AOI221x1_ASAP7_75t_SL g984 ( .A1(n_204), .A2(n_291), .B1(n_680), .B2(n_985), .C(n_986), .Y(n_984) );
INVx1_ASAP7_75t_L g1963 ( .A(n_205), .Y(n_1963) );
AOI221x1_ASAP7_75t_SL g1075 ( .A1(n_206), .A2(n_287), .B1(n_1076), .B2(n_1077), .C(n_1079), .Y(n_1075) );
AOI21xp33_ASAP7_75t_L g1136 ( .A1(n_206), .A2(n_563), .B(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g607 ( .A(n_207), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_207), .A2(n_328), .B1(n_702), .B2(n_705), .Y(n_701) );
INVxp67_ASAP7_75t_SL g1618 ( .A(n_208), .Y(n_1618) );
AOI22xp33_ASAP7_75t_L g1624 ( .A1(n_208), .A2(n_215), .B1(n_586), .B2(n_1552), .Y(n_1624) );
AOI21xp33_ASAP7_75t_L g974 ( .A1(n_209), .A2(n_975), .B(n_976), .Y(n_974) );
INVx1_ASAP7_75t_L g994 ( .A(n_209), .Y(n_994) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_210), .A2(n_288), .B1(n_615), .B2(n_619), .C(n_624), .Y(n_614) );
INVx1_ASAP7_75t_L g691 ( .A(n_210), .Y(n_691) );
INVx2_ASAP7_75t_L g1684 ( .A(n_211), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_211), .B(n_323), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_211), .B(n_1690), .Y(n_1692) );
INVx1_ASAP7_75t_L g531 ( .A(n_212), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g1932 ( .A(n_213), .Y(n_1932) );
INVxp67_ASAP7_75t_SL g1612 ( .A(n_215), .Y(n_1612) );
INVx1_ASAP7_75t_L g537 ( .A(n_216), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_217), .A2(n_313), .B1(n_971), .B2(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1576 ( .A(n_217), .Y(n_1576) );
INVx1_ASAP7_75t_L g1600 ( .A(n_218), .Y(n_1600) );
INVx1_ASAP7_75t_L g1308 ( .A(n_219), .Y(n_1308) );
INVx1_ASAP7_75t_L g1004 ( .A(n_220), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g1714 ( .A1(n_221), .A2(n_279), .B1(n_1681), .B2(n_1691), .Y(n_1714) );
INVx1_ASAP7_75t_L g907 ( .A(n_223), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_224), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1715 ( .A1(n_225), .A2(n_230), .B1(n_1688), .B2(n_1707), .Y(n_1715) );
INVx1_ASAP7_75t_L g547 ( .A(n_226), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_227), .A2(n_360), .B1(n_1325), .B2(n_1326), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_227), .A2(n_234), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
XNOR2xp5_ASAP7_75t_L g1957 ( .A(n_228), .B(n_1958), .Y(n_1957) );
OAI211xp5_ASAP7_75t_L g1002 ( .A1(n_229), .A2(n_895), .B(n_921), .C(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1054 ( .A(n_229), .Y(n_1054) );
INVx1_ASAP7_75t_L g1392 ( .A(n_231), .Y(n_1392) );
OAI211xp5_ASAP7_75t_L g1399 ( .A1(n_231), .A2(n_957), .B(n_1400), .C(n_1402), .Y(n_1399) );
XOR2x2_ASAP7_75t_L g715 ( .A(n_232), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1901 ( .A(n_233), .Y(n_1901) );
AOI22xp33_ASAP7_75t_SL g1338 ( .A1(n_234), .A2(n_354), .B1(n_1325), .B2(n_1339), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_235), .A2(n_330), .B1(n_680), .B2(n_683), .Y(n_1256) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_236), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g1905 ( .A(n_237), .Y(n_1905) );
INVx1_ASAP7_75t_L g890 ( .A(n_238), .Y(n_890) );
INVx1_ASAP7_75t_L g1948 ( .A(n_239), .Y(n_1948) );
AOI22xp33_ASAP7_75t_L g1952 ( .A1(n_239), .A2(n_1953), .B1(n_1956), .B2(n_1995), .Y(n_1952) );
INVx1_ASAP7_75t_L g1575 ( .A(n_240), .Y(n_1575) );
INVx1_ASAP7_75t_L g1193 ( .A(n_241), .Y(n_1193) );
INVx2_ASAP7_75t_L g503 ( .A(n_242), .Y(n_503) );
INVx1_ASAP7_75t_L g575 ( .A(n_242), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_242), .B(n_465), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g1708 ( .A1(n_243), .A2(n_366), .B1(n_1688), .B2(n_1691), .Y(n_1708) );
INVx1_ASAP7_75t_L g1974 ( .A(n_244), .Y(n_1974) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_246), .A2(n_256), .B1(n_781), .B2(n_782), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_246), .A2(n_256), .B1(n_794), .B2(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g1940 ( .A(n_247), .Y(n_1940) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_249), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g1560 ( .A(n_250), .B(n_620), .Y(n_1560) );
INVxp67_ASAP7_75t_SL g1585 ( .A(n_250), .Y(n_1585) );
INVx1_ASAP7_75t_L g926 ( .A(n_251), .Y(n_926) );
INVx1_ASAP7_75t_L g1916 ( .A(n_252), .Y(n_1916) );
INVx1_ASAP7_75t_L g550 ( .A(n_253), .Y(n_550) );
INVx1_ASAP7_75t_L g1968 ( .A(n_254), .Y(n_1968) );
OAI22xp33_ASAP7_75t_L g1439 ( .A1(n_257), .A2(n_285), .B1(n_391), .B2(n_445), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_257), .A2(n_285), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
BUFx3_ASAP7_75t_L g461 ( .A(n_258), .Y(n_461) );
INVx1_ASAP7_75t_L g1545 ( .A(n_259), .Y(n_1545) );
INVx1_ASAP7_75t_L g1607 ( .A(n_261), .Y(n_1607) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_262), .A2(n_281), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_263), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1582 ( .A(n_264), .Y(n_1582) );
OAI22xp5_ASAP7_75t_SL g949 ( .A1(n_265), .A2(n_310), .B1(n_644), .B2(n_656), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_265), .Y(n_960) );
INVx1_ASAP7_75t_L g1291 ( .A(n_266), .Y(n_1291) );
INVx1_ASAP7_75t_L g1478 ( .A(n_267), .Y(n_1478) );
INVx1_ASAP7_75t_L g1554 ( .A(n_268), .Y(n_1554) );
XOR2xp5_ASAP7_75t_L g1500 ( .A(n_269), .B(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1508 ( .A(n_270), .Y(n_1508) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_271), .Y(n_725) );
AOI21xp33_ASAP7_75t_L g1212 ( .A1(n_272), .A2(n_975), .B(n_976), .Y(n_1212) );
INVx1_ASAP7_75t_L g877 ( .A(n_274), .Y(n_877) );
INVx1_ASAP7_75t_L g1020 ( .A(n_275), .Y(n_1020) );
INVx1_ASAP7_75t_L g1110 ( .A(n_276), .Y(n_1110) );
INVx1_ASAP7_75t_L g1610 ( .A(n_277), .Y(n_1610) );
INVx1_ASAP7_75t_L g1249 ( .A(n_278), .Y(n_1249) );
INVx1_ASAP7_75t_L g515 ( .A(n_280), .Y(n_515) );
BUFx3_ASAP7_75t_L g399 ( .A(n_282), .Y(n_399) );
INVx1_ASAP7_75t_L g437 ( .A(n_282), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g1633 ( .A(n_283), .Y(n_1633) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_284), .A2(n_327), .B1(n_1318), .B2(n_1394), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_284), .A2(n_327), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
XNOR2xp5_ASAP7_75t_L g801 ( .A(n_286), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g1133 ( .A(n_287), .Y(n_1133) );
INVx1_ASAP7_75t_L g696 ( .A(n_288), .Y(n_696) );
INVx1_ASAP7_75t_L g1064 ( .A(n_290), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_291), .A2(n_296), .B1(n_970), .B2(n_971), .Y(n_977) );
INVx1_ASAP7_75t_L g817 ( .A(n_292), .Y(n_817) );
INVx1_ASAP7_75t_L g1005 ( .A(n_293), .Y(n_1005) );
OAI211xp5_ASAP7_75t_L g1048 ( .A1(n_293), .A2(n_558), .B(n_1049), .C(n_1050), .Y(n_1048) );
OAI221xp5_ASAP7_75t_L g1645 ( .A1(n_294), .A2(n_361), .B1(n_615), .B2(n_619), .C(n_1646), .Y(n_1645) );
OAI22xp5_ASAP7_75t_L g1658 ( .A1(n_294), .A2(n_361), .B1(n_946), .B2(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g871 ( .A(n_295), .Y(n_871) );
INVx1_ASAP7_75t_L g1420 ( .A(n_297), .Y(n_1420) );
INVx1_ASAP7_75t_L g1481 ( .A(n_298), .Y(n_1481) );
INVx1_ASAP7_75t_L g1510 ( .A(n_299), .Y(n_1510) );
INVx1_ASAP7_75t_L g1914 ( .A(n_300), .Y(n_1914) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_301), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_302), .A2(n_374), .B1(n_857), .B2(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1026 ( .A(n_303), .Y(n_1026) );
INVx1_ASAP7_75t_L g1375 ( .A(n_304), .Y(n_1375) );
INVx1_ASAP7_75t_L g1505 ( .A(n_305), .Y(n_1505) );
CKINVDCx5p33_ASAP7_75t_R g1168 ( .A(n_306), .Y(n_1168) );
INVx1_ASAP7_75t_L g1614 ( .A(n_309), .Y(n_1614) );
INVx1_ASAP7_75t_L g953 ( .A(n_310), .Y(n_953) );
INVx1_ASAP7_75t_L g463 ( .A(n_311), .Y(n_463) );
INVx1_ASAP7_75t_L g475 ( .A(n_311), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_312), .Y(n_776) );
INVxp67_ASAP7_75t_SL g1568 ( .A(n_313), .Y(n_1568) );
INVx1_ASAP7_75t_L g873 ( .A(n_314), .Y(n_873) );
OAI211xp5_ASAP7_75t_L g1440 ( .A1(n_315), .A2(n_917), .B(n_921), .C(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1452 ( .A(n_315), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_317), .Y(n_727) );
INVx1_ASAP7_75t_L g973 ( .A(n_318), .Y(n_973) );
INVx1_ASAP7_75t_L g1378 ( .A(n_319), .Y(n_1378) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_321), .A2(n_999), .B1(n_1000), .B2(n_1057), .Y(n_998) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_321), .Y(n_1057) );
AOI22xp5_ASAP7_75t_SL g1711 ( .A1(n_321), .A2(n_371), .B1(n_1681), .B2(n_1707), .Y(n_1711) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_322), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_323), .B(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1690 ( .A(n_323), .Y(n_1690) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_324), .Y(n_742) );
INVx1_ASAP7_75t_L g1150 ( .A(n_326), .Y(n_1150) );
INVx1_ASAP7_75t_L g610 ( .A(n_328), .Y(n_610) );
INVx1_ASAP7_75t_L g1476 ( .A(n_329), .Y(n_1476) );
INVx1_ASAP7_75t_L g1280 ( .A(n_330), .Y(n_1280) );
INVx1_ASAP7_75t_L g539 ( .A(n_331), .Y(n_539) );
INVx1_ASAP7_75t_L g426 ( .A(n_332), .Y(n_426) );
OAI211xp5_ASAP7_75t_L g469 ( .A1(n_332), .A2(n_470), .B(n_477), .C(n_481), .Y(n_469) );
INVxp67_ASAP7_75t_SL g1944 ( .A(n_333), .Y(n_1944) );
INVx1_ASAP7_75t_L g1221 ( .A(n_334), .Y(n_1221) );
INVx1_ASAP7_75t_L g779 ( .A(n_335), .Y(n_779) );
OAI211xp5_ASAP7_75t_L g787 ( .A1(n_335), .A2(n_477), .B(n_788), .C(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g1414 ( .A(n_336), .Y(n_1414) );
INVx1_ASAP7_75t_L g1515 ( .A(n_338), .Y(n_1515) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_339), .A2(n_1297), .B1(n_1351), .B2(n_1352), .Y(n_1296) );
INVxp67_ASAP7_75t_SL g1352 ( .A(n_339), .Y(n_1352) );
INVx1_ASAP7_75t_L g1667 ( .A(n_341), .Y(n_1667) );
AOI211xp5_ASAP7_75t_SL g1188 ( .A1(n_342), .A2(n_1189), .B(n_1190), .C(n_1192), .Y(n_1188) );
INVx1_ASAP7_75t_L g1971 ( .A(n_343), .Y(n_1971) );
AOI21xp5_ASAP7_75t_SL g1216 ( .A1(n_344), .A2(n_975), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1229 ( .A(n_344), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_345), .A2(n_372), .B1(n_490), .B2(n_496), .Y(n_489) );
INVx1_ASAP7_75t_L g1279 ( .A(n_347), .Y(n_1279) );
INVx1_ASAP7_75t_L g1362 ( .A(n_348), .Y(n_1362) );
XOR2x2_ASAP7_75t_L g1357 ( .A(n_349), .B(n_1358), .Y(n_1357) );
INVxp67_ASAP7_75t_L g1235 ( .A(n_350), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_351), .Y(n_721) );
INVxp67_ASAP7_75t_SL g1248 ( .A(n_352), .Y(n_1248) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_353), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g1344 ( .A1(n_354), .A2(n_360), .B1(n_675), .B2(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1018 ( .A(n_355), .Y(n_1018) );
INVx1_ASAP7_75t_L g1032 ( .A(n_356), .Y(n_1032) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_359), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g1570 ( .A(n_363), .Y(n_1570) );
INVx1_ASAP7_75t_L g1488 ( .A(n_364), .Y(n_1488) );
INVx1_ASAP7_75t_L g908 ( .A(n_365), .Y(n_908) );
OAI211xp5_ASAP7_75t_L g916 ( .A1(n_365), .A2(n_917), .B(n_918), .C(n_921), .Y(n_916) );
INVx1_ASAP7_75t_L g454 ( .A(n_367), .Y(n_454) );
INVx2_ASAP7_75t_L g512 ( .A(n_367), .Y(n_512) );
INVx1_ASAP7_75t_L g574 ( .A(n_367), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_368), .Y(n_1102) );
INVx1_ASAP7_75t_L g948 ( .A(n_369), .Y(n_948) );
INVx1_ASAP7_75t_L g1643 ( .A(n_370), .Y(n_1643) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_373), .Y(n_1152) );
INVx1_ASAP7_75t_L g1302 ( .A(n_374), .Y(n_1302) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_400), .B(n_1675), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1951 ( .A(n_379), .B(n_388), .Y(n_1951) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1955 ( .A(n_381), .B(n_384), .Y(n_1955) );
INVx1_ASAP7_75t_L g1997 ( .A(n_381), .Y(n_1997) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1999 ( .A(n_384), .B(n_1997), .Y(n_1999) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g450 ( .A(n_388), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g545 ( .A(n_389), .B(n_399), .Y(n_545) );
AND2x4_ASAP7_75t_L g635 ( .A(n_389), .B(n_398), .Y(n_635) );
INVx1_ASAP7_75t_L g1007 ( .A(n_390), .Y(n_1007) );
INVxp67_ASAP7_75t_SL g1310 ( .A(n_390), .Y(n_1310) );
INVx1_ASAP7_75t_L g1536 ( .A(n_390), .Y(n_1536) );
AND2x4_ASAP7_75t_SL g1950 ( .A(n_390), .B(n_1951), .Y(n_1950) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
OR2x6_ASAP7_75t_L g435 ( .A(n_392), .B(n_436), .Y(n_435) );
BUFx4f_ASAP7_75t_L g838 ( .A(n_392), .Y(n_838) );
INVx1_ASAP7_75t_L g901 ( .A(n_392), .Y(n_901) );
INVxp67_ASAP7_75t_L g1364 ( .A(n_392), .Y(n_1364) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx4f_ASAP7_75t_L g518 ( .A(n_393), .Y(n_518) );
INVx3_ASAP7_75t_L g627 ( .A(n_393), .Y(n_627) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2x1_ASAP7_75t_L g414 ( .A(n_395), .B(n_396), .Y(n_414) );
AND2x2_ASAP7_75t_L g419 ( .A(n_395), .B(n_396), .Y(n_419) );
INVx1_ASAP7_75t_L g431 ( .A(n_395), .Y(n_431) );
INVx2_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
AND2x2_ASAP7_75t_L g447 ( .A(n_395), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g530 ( .A(n_395), .Y(n_530) );
BUFx2_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_396), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g448 ( .A(n_396), .Y(n_448) );
OR2x2_ASAP7_75t_L g529 ( .A(n_396), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g587 ( .A(n_396), .B(n_443), .Y(n_587) );
INVx1_ASAP7_75t_L g601 ( .A(n_396), .Y(n_601) );
OR2x6_ASAP7_75t_L g847 ( .A(n_397), .B(n_627), .Y(n_847) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g424 ( .A(n_399), .Y(n_424) );
AND2x4_ASAP7_75t_L g429 ( .A(n_399), .B(n_430), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_1353), .B1(n_1354), .B2(n_1674), .Y(n_400) );
INVx1_ASAP7_75t_L g1674 ( .A(n_401), .Y(n_1674) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_860), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_713), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_580), .B2(n_712), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_455), .C(n_507), .Y(n_408) );
OAI31xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_432), .A3(n_444), .B(n_449), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_411), .A2(n_877), .B1(n_885), .B2(n_898), .Y(n_897) );
OAI211xp5_ASAP7_75t_L g964 ( .A1(n_411), .A2(n_965), .B(n_966), .C(n_969), .Y(n_964) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g538 ( .A(n_412), .Y(n_538) );
INVx2_ASAP7_75t_L g761 ( .A(n_412), .Y(n_761) );
INVx1_ASAP7_75t_L g957 ( .A(n_412), .Y(n_957) );
INVx2_ASAP7_75t_L g1521 ( .A(n_412), .Y(n_1521) );
INVx4_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx4f_ASAP7_75t_L g532 ( .A(n_413), .Y(n_532) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_413), .Y(n_756) );
BUFx4f_ASAP7_75t_L g895 ( .A(n_413), .Y(n_895) );
BUFx4f_ASAP7_75t_L g1089 ( .A(n_413), .Y(n_1089) );
OR2x6_ASAP7_75t_L g1092 ( .A(n_413), .B(n_1093), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g1290 ( .A1(n_413), .A2(n_536), .B1(n_545), .B2(n_1291), .C(n_1292), .Y(n_1290) );
BUFx4f_ASAP7_75t_L g1370 ( .A(n_413), .Y(n_1370) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g773 ( .A(n_414), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_415), .B(n_1300), .C(n_1305), .Y(n_1299) );
NAND3xp33_ASAP7_75t_L g1594 ( .A(n_415), .B(n_1595), .C(n_1598), .Y(n_1594) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g921 ( .A(n_416), .Y(n_921) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_417), .B(n_1328), .Y(n_1401) );
BUFx3_ASAP7_75t_L g591 ( .A(n_418), .Y(n_591) );
AND2x6_ASAP7_75t_L g604 ( .A(n_418), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_418), .B(n_588), .Y(n_618) );
INVx1_ASAP7_75t_L g633 ( .A(n_418), .Y(n_633) );
BUFx6f_ASAP7_75t_L g1078 ( .A(n_418), .Y(n_1078) );
BUFx3_ASAP7_75t_L g1189 ( .A(n_418), .Y(n_1189) );
BUFx3_ASAP7_75t_L g1650 ( .A(n_418), .Y(n_1650) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g1329 ( .A(n_419), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_426), .B2(n_427), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_421), .A2(n_482), .B1(n_486), .B2(n_487), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_422), .A2(n_907), .B1(n_919), .B2(n_920), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_422), .A2(n_919), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_422), .A2(n_427), .B1(n_1531), .B2(n_1539), .Y(n_1538) );
AOI222xp33_ASAP7_75t_L g1598 ( .A1(n_422), .A2(n_591), .B1(n_843), .B2(n_1599), .C1(n_1600), .C2(n_1601), .Y(n_1598) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g1441 ( .A1(n_423), .A2(n_429), .B1(n_1442), .B2(n_1443), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_423), .A2(n_429), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OR2x2_ASAP7_75t_L g440 ( .A(n_424), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g775 ( .A(n_424), .B(n_425), .Y(n_775) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_424), .B(n_955), .Y(n_1301) );
INVx1_ASAP7_75t_L g622 ( .A(n_425), .Y(n_622) );
BUFx2_ASAP7_75t_L g959 ( .A(n_425), .Y(n_959) );
INVx1_ASAP7_75t_L g1099 ( .A(n_425), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_425), .A2(n_961), .B1(n_1147), .B2(n_1166), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_427), .A2(n_775), .B1(n_1391), .B2(n_1403), .Y(n_1402) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g778 ( .A(n_429), .Y(n_778) );
BUFx3_ASAP7_75t_L g919 ( .A(n_429), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_430), .B(n_605), .Y(n_655) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g781 ( .A(n_435), .Y(n_781) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_435), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g1405 ( .A(n_435), .Y(n_1405) );
AND2x4_ASAP7_75t_L g446 ( .A(n_436), .B(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g1303 ( .A(n_438), .Y(n_1303) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g783 ( .A(n_440), .Y(n_783) );
BUFx2_ASAP7_75t_L g915 ( .A(n_440), .Y(n_915) );
INVx8_ASAP7_75t_L g523 ( .A(n_441), .Y(n_523) );
BUFx2_ASAP7_75t_L g629 ( .A(n_441), .Y(n_629) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g768 ( .A(n_446), .Y(n_768) );
INVx3_ASAP7_75t_SL g1008 ( .A(n_446), .Y(n_1008) );
INVx2_ASAP7_75t_L g595 ( .A(n_447), .Y(n_595) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_447), .Y(n_613) );
BUFx3_ASAP7_75t_L g967 ( .A(n_447), .Y(n_967) );
OAI31xp33_ASAP7_75t_L g766 ( .A1(n_449), .A2(n_767), .A3(n_769), .B(n_780), .Y(n_766) );
OAI31xp33_ASAP7_75t_L g1397 ( .A1(n_449), .A2(n_1398), .A3(n_1399), .B(n_1404), .Y(n_1397) );
OAI31xp33_ASAP7_75t_SL g1534 ( .A1(n_449), .A2(n_1535), .A3(n_1537), .B(n_1540), .Y(n_1534) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI31xp33_ASAP7_75t_L g839 ( .A1(n_450), .A2(n_840), .A3(n_845), .B(n_846), .Y(n_839) );
BUFx2_ASAP7_75t_SL g922 ( .A(n_450), .Y(n_922) );
OAI31xp33_ASAP7_75t_L g1001 ( .A1(n_450), .A2(n_1002), .A3(n_1006), .B(n_1009), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_450), .Y(n_1311) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g654 ( .A(n_452), .B(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g663 ( .A(n_452), .Y(n_663) );
INVx1_ASAP7_75t_L g933 ( .A(n_452), .Y(n_933) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI31xp33_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_469), .A3(n_489), .B(n_500), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_459), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1447 ( .A(n_459), .Y(n_1447) );
INVx1_ASAP7_75t_L g1528 ( .A(n_459), .Y(n_1528) );
OR2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
OR2x4_ASAP7_75t_L g467 ( .A(n_460), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g557 ( .A(n_460), .Y(n_557) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_460), .Y(n_578) );
BUFx3_ASAP7_75t_L g724 ( .A(n_460), .Y(n_724) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_460), .Y(n_1128) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_461), .Y(n_476) );
AND2x4_ASAP7_75t_L g479 ( .A(n_461), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g495 ( .A(n_461), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_461), .B(n_475), .Y(n_499) );
INVx1_ASAP7_75t_L g660 ( .A(n_462), .Y(n_660) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
INVx1_ASAP7_75t_L g468 ( .A(n_464), .Y(n_468) );
AND2x4_ASAP7_75t_L g478 ( .A(n_464), .B(n_479), .Y(n_478) );
OR2x6_ASAP7_75t_L g497 ( .A(n_464), .B(n_498), .Y(n_497) );
NAND3x1_ASAP7_75t_L g572 ( .A(n_464), .B(n_573), .C(n_575), .Y(n_572) );
AND2x4_ASAP7_75t_L g661 ( .A(n_464), .B(n_662), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_464), .B(n_575), .Y(n_686) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g484 ( .A(n_465), .Y(n_484) );
NAND2xp33_ASAP7_75t_SL g554 ( .A(n_465), .B(n_503), .Y(n_554) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g795 ( .A(n_467), .Y(n_795) );
BUFx3_ASAP7_75t_L g1318 ( .A(n_467), .Y(n_1318) );
BUFx2_ASAP7_75t_L g1454 ( .A(n_467), .Y(n_1454) );
AND2x4_ASAP7_75t_L g491 ( .A(n_468), .B(n_492), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g1937 ( .A1(n_470), .A2(n_1925), .B1(n_1938), .B2(n_1940), .Y(n_1937) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g995 ( .A(n_471), .Y(n_995) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g656 ( .A(n_472), .B(n_646), .Y(n_656) );
INVx4_ASAP7_75t_L g790 ( .A(n_472), .Y(n_790) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_472), .Y(n_824) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g560 ( .A(n_473), .Y(n_560) );
BUFx2_ASAP7_75t_L g745 ( .A(n_473), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
BUFx2_ASAP7_75t_L g488 ( .A(n_474), .Y(n_488) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g480 ( .A(n_475), .Y(n_480) );
BUFx2_ASAP7_75t_L g485 ( .A(n_476), .Y(n_485) );
AND2x4_ASAP7_75t_L g677 ( .A(n_476), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g694 ( .A(n_476), .Y(n_694) );
CKINVDCx8_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
CKINVDCx8_ASAP7_75t_R g1049 ( .A(n_478), .Y(n_1049) );
OAI31xp33_ASAP7_75t_L g1239 ( .A1(n_478), .A2(n_1240), .A3(n_1250), .B(n_1251), .Y(n_1239) );
BUFx2_ASAP7_75t_L g672 ( .A(n_479), .Y(n_672) );
INVx2_ASAP7_75t_L g689 ( .A(n_479), .Y(n_689) );
BUFx2_ASAP7_75t_L g711 ( .A(n_479), .Y(n_711) );
BUFx3_ASAP7_75t_L g1113 ( .A(n_479), .Y(n_1113) );
BUFx2_ASAP7_75t_L g1122 ( .A(n_479), .Y(n_1122) );
BUFx2_ASAP7_75t_L g1237 ( .A(n_479), .Y(n_1237) );
BUFx2_ASAP7_75t_L g1630 ( .A(n_479), .Y(n_1630) );
INVx1_ASAP7_75t_L g678 ( .A(n_480), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_482), .A2(n_487), .B1(n_776), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_482), .A2(n_487), .B1(n_842), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_482), .A2(n_487), .B1(n_907), .B2(n_908), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_482), .A2(n_487), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_482), .A2(n_487), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_482), .A2(n_487), .B1(n_1463), .B2(n_1471), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_482), .A2(n_487), .B1(n_1531), .B2(n_1532), .Y(n_1530) );
AOI22xp33_ASAP7_75t_SL g1993 ( .A1(n_482), .A2(n_487), .B1(n_1986), .B2(n_1994), .Y(n_1993) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
AND2x4_ASAP7_75t_L g487 ( .A(n_483), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_483), .B(n_485), .Y(n_1052) );
A2O1A1Ixp33_ASAP7_75t_L g1240 ( .A1(n_483), .A2(n_1241), .B(n_1244), .C(n_1247), .Y(n_1240) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND3x4_ASAP7_75t_L g667 ( .A(n_484), .B(n_503), .C(n_640), .Y(n_667) );
BUFx6f_ASAP7_75t_L g1053 ( .A(n_487), .Y(n_1053) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g786 ( .A(n_491), .Y(n_786) );
INVx2_ASAP7_75t_L g850 ( .A(n_491), .Y(n_850) );
INVxp67_ASAP7_75t_L g1314 ( .A(n_491), .Y(n_1314) );
INVx1_ASAP7_75t_L g1448 ( .A(n_491), .Y(n_1448) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_492), .Y(n_674) );
INVx1_ASAP7_75t_L g728 ( .A(n_492), .Y(n_728) );
BUFx6f_ASAP7_75t_L g1132 ( .A(n_492), .Y(n_1132) );
INVx2_ASAP7_75t_L g1611 ( .A(n_492), .Y(n_1611) );
INVx2_ASAP7_75t_L g1936 ( .A(n_492), .Y(n_1936) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx8_ASAP7_75t_L g563 ( .A(n_493), .Y(n_563) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_493), .Y(n_682) );
INVx2_ASAP7_75t_L g816 ( .A(n_493), .Y(n_816) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x4_ASAP7_75t_L g659 ( .A(n_495), .B(n_660), .Y(n_659) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g797 ( .A(n_497), .Y(n_797) );
INVx2_ASAP7_75t_L g858 ( .A(n_497), .Y(n_858) );
INVx1_ASAP7_75t_L g1395 ( .A(n_497), .Y(n_1395) );
BUFx3_ASAP7_75t_L g564 ( .A(n_498), .Y(n_564) );
INVx1_ASAP7_75t_L g732 ( .A(n_498), .Y(n_732) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g569 ( .A(n_499), .Y(n_569) );
OAI31xp33_ASAP7_75t_SL g903 ( .A1(n_500), .A2(n_904), .A3(n_905), .B(n_909), .Y(n_903) );
OAI31xp33_ASAP7_75t_L g1044 ( .A1(n_500), .A2(n_1045), .A3(n_1048), .B(n_1055), .Y(n_1044) );
OAI31xp33_ASAP7_75t_L g1445 ( .A1(n_500), .A2(n_1446), .A3(n_1449), .B(n_1453), .Y(n_1445) );
OAI31xp33_ASAP7_75t_L g1525 ( .A1(n_500), .A2(n_1526), .A3(n_1529), .B(n_1533), .Y(n_1525) );
OAI21xp33_ASAP7_75t_L g1625 ( .A1(n_500), .A2(n_1626), .B(n_1632), .Y(n_1625) );
AND2x2_ASAP7_75t_SL g500 ( .A(n_501), .B(n_504), .Y(n_500) );
AND2x4_ASAP7_75t_L g798 ( .A(n_501), .B(n_504), .Y(n_798) );
AND2x2_ASAP7_75t_L g859 ( .A(n_501), .B(n_504), .Y(n_859) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_501), .B(n_504), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_501), .B(n_504), .Y(n_1396) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g662 ( .A(n_503), .Y(n_662) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
OR2x2_ASAP7_75t_L g553 ( .A(n_506), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g646 ( .A(n_506), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_SL g836 ( .A(n_506), .B(n_545), .Y(n_836) );
NOR2xp33_ASAP7_75t_SL g507 ( .A(n_508), .B(n_551), .Y(n_507) );
OAI33xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_514), .A3(n_524), .B1(n_533), .B2(n_540), .B3(n_546), .Y(n_508) );
OAI33xp33_ASAP7_75t_L g1033 ( .A1(n_509), .A2(n_540), .A3(n_1034), .B1(n_1040), .B2(n_1042), .B3(n_1043), .Y(n_1033) );
INVx1_ASAP7_75t_L g1085 ( .A(n_509), .Y(n_1085) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g749 ( .A(n_510), .Y(n_749) );
INVx4_ASAP7_75t_L g829 ( .A(n_510), .Y(n_829) );
INVx2_ASAP7_75t_L g892 ( .A(n_510), .Y(n_892) );
INVx2_ASAP7_75t_L g1479 ( .A(n_510), .Y(n_1479) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
OR2x6_ASAP7_75t_L g685 ( .A(n_511), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g1141 ( .A(n_511), .Y(n_1141) );
BUFx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g640 ( .A(n_512), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_512), .B(n_605), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_519), .B2(n_520), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_515), .A2(n_537), .B1(n_556), .B2(n_558), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_516), .A2(n_547), .B1(n_548), .B2(n_550), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_516), .A2(n_520), .B1(n_870), .B2(n_888), .Y(n_893) );
OAI22xp33_ASAP7_75t_L g1519 ( .A1(n_516), .A2(n_548), .B1(n_1505), .B2(n_1515), .Y(n_1519) );
OAI22xp33_ASAP7_75t_L g1524 ( .A1(n_516), .A2(n_548), .B1(n_1510), .B2(n_1513), .Y(n_1524) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g1429 ( .A(n_517), .Y(n_1429) );
INVx2_ASAP7_75t_L g1436 ( .A(n_517), .Y(n_1436) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g1037 ( .A(n_518), .Y(n_1037) );
INVx4_ASAP7_75t_L g1194 ( .A(n_518), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_539), .B1(n_577), .B2(n_579), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_520), .A2(n_534), .B1(n_871), .B2(n_890), .Y(n_896) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_522), .A2(n_1362), .B1(n_1363), .B2(n_1365), .Y(n_1361) );
HB1xp67_ASAP7_75t_L g1915 ( .A(n_522), .Y(n_1915) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g549 ( .A(n_523), .Y(n_549) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_523), .Y(n_752) );
INVx2_ASAP7_75t_L g765 ( .A(n_523), .Y(n_765) );
INVx4_ASAP7_75t_L g831 ( .A(n_523), .Y(n_831) );
INVx2_ASAP7_75t_L g1083 ( .A(n_523), .Y(n_1083) );
INVx2_ASAP7_75t_L g1284 ( .A(n_523), .Y(n_1284) );
INVx1_ASAP7_75t_L g1430 ( .A(n_523), .Y(n_1430) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_531), .B2(n_532), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_525), .A2(n_547), .B1(n_562), .B2(n_564), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_526), .A2(n_873), .B1(n_882), .B2(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g1368 ( .A(n_527), .Y(n_1368) );
INVx2_ASAP7_75t_L g1433 ( .A(n_527), .Y(n_1433) );
INVx4_ASAP7_75t_L g1484 ( .A(n_527), .Y(n_1484) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g536 ( .A(n_529), .Y(n_536) );
INVx1_ASAP7_75t_L g755 ( .A(n_529), .Y(n_755) );
INVx2_ASAP7_75t_L g760 ( .A(n_529), .Y(n_760) );
BUFx2_ASAP7_75t_L g833 ( .A(n_529), .Y(n_833) );
AND2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_530), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_531), .A2(n_550), .B1(n_566), .B2(n_567), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_532), .A2(n_1020), .B1(n_1025), .B2(n_1041), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_532), .A2(n_1018), .B1(n_1032), .B2(n_1041), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_537), .B1(n_538), .B2(n_539), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g1190 ( .A1(n_536), .A2(n_545), .B(n_1191), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1483 ( .A1(n_538), .A2(n_1484), .B1(n_1485), .B2(n_1486), .Y(n_1483) );
OAI22xp5_ASAP7_75t_L g1980 ( .A1(n_538), .A2(n_1484), .B1(n_1964), .B2(n_1974), .Y(n_1980) );
OAI33xp33_ASAP7_75t_L g1518 ( .A1(n_540), .A2(n_748), .A3(n_1519), .B1(n_1520), .B2(n_1522), .B3(n_1524), .Y(n_1518) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x4_ASAP7_75t_L g763 ( .A(n_543), .B(n_545), .Y(n_763) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_SL g596 ( .A(n_545), .Y(n_596) );
INVx4_ASAP7_75t_L g976 ( .A(n_545), .Y(n_976) );
INVx4_ASAP7_75t_L g1918 ( .A(n_545), .Y(n_1918) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI33xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .A3(n_561), .B1(n_565), .B2(n_570), .B3(n_576), .Y(n_551) );
BUFx4f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx8_ASAP7_75t_L g719 ( .A(n_553), .Y(n_719) );
BUFx2_ASAP7_75t_L g805 ( .A(n_553), .Y(n_805) );
BUFx4f_ASAP7_75t_L g868 ( .A(n_553), .Y(n_868) );
BUFx2_ASAP7_75t_L g1137 ( .A(n_554), .Y(n_1137) );
OR2x2_ASAP7_75t_L g702 ( .A(n_556), .B(n_703), .Y(n_702) );
OR2x6_ASAP7_75t_L g934 ( .A(n_556), .B(n_703), .Y(n_934) );
INVx2_ASAP7_75t_SL g1017 ( .A(n_556), .Y(n_1017) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_556), .A2(n_995), .B1(n_1505), .B2(n_1506), .Y(n_1504) );
OAI22xp33_ASAP7_75t_L g1514 ( .A1(n_556), .A2(n_1515), .B1(n_1516), .B2(n_1517), .Y(n_1514) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g809 ( .A(n_557), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_558), .A2(n_721), .B1(n_722), .B2(n_725), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_558), .A2(n_1016), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g1608 ( .A(n_559), .Y(n_1608) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_560), .Y(n_579) );
HB1xp67_ASAP7_75t_L g1415 ( .A(n_560), .Y(n_1415) );
HB1xp67_ASAP7_75t_L g1426 ( .A(n_560), .Y(n_1426) );
OAI22xp33_ASAP7_75t_L g1496 ( .A1(n_560), .A2(n_809), .B1(n_1478), .B2(n_1486), .Y(n_1496) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g566 ( .A(n_563), .Y(n_566) );
AND2x4_ASAP7_75t_L g706 ( .A(n_563), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g991 ( .A(n_563), .Y(n_991) );
INVx2_ASAP7_75t_SL g1495 ( .A(n_563), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g1419 ( .A1(n_564), .A2(n_1420), .B1(n_1421), .B2(n_1422), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1609 ( .A1(n_564), .A2(n_1610), .B1(n_1611), .B2(n_1612), .Y(n_1609) );
OAI221xp5_ASAP7_75t_L g1943 ( .A1(n_564), .A2(n_735), .B1(n_1916), .B2(n_1944), .C(n_1945), .Y(n_1943) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_566), .A2(n_1023), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
INVx1_ASAP7_75t_L g1348 ( .A(n_566), .Y(n_1348) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_567), .A2(n_814), .B1(n_815), .B2(n_817), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g1494 ( .A1(n_567), .A2(n_1482), .B1(n_1489), .B2(n_1495), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1934 ( .A1(n_567), .A2(n_1914), .B1(n_1935), .B2(n_1936), .Y(n_1934) );
OAI22xp5_ASAP7_75t_L g1969 ( .A1(n_567), .A2(n_1495), .B1(n_1970), .B2(n_1971), .Y(n_1969) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
CKINVDCx8_ASAP7_75t_R g737 ( .A(n_568), .Y(n_737) );
INVx3_ASAP7_75t_L g889 ( .A(n_568), .Y(n_889) );
INVx3_ASAP7_75t_L g1023 ( .A(n_568), .Y(n_1023) );
INVx1_ASAP7_75t_L g1493 ( .A(n_568), .Y(n_1493) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
OAI33xp33_ASAP7_75t_L g866 ( .A1(n_570), .A2(n_867), .A3(n_869), .B1(n_872), .B2(n_879), .B3(n_886), .Y(n_866) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_571), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_571), .A2(n_710), .B1(n_984), .B2(n_989), .C(n_996), .Y(n_983) );
INVx2_ASAP7_75t_L g1238 ( .A(n_571), .Y(n_1238) );
NAND3xp33_ASAP7_75t_L g1346 ( .A(n_571), .B(n_1347), .C(n_1350), .Y(n_1346) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g1029 ( .A(n_572), .Y(n_1029) );
OAI33xp33_ASAP7_75t_L g1379 ( .A1(n_572), .A2(n_719), .A3(n_1380), .B1(n_1382), .B2(n_1383), .B3(n_1385), .Y(n_1379) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g649 ( .A(n_574), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_574), .B(n_588), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g869 ( .A1(n_577), .A2(n_579), .B1(n_870), .B2(n_871), .Y(n_869) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_578), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_578), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
INVx1_ASAP7_75t_L g1939 ( .A(n_578), .Y(n_1939) );
OAI22xp5_ASAP7_75t_L g1569 ( .A1(n_579), .A2(n_1570), .B1(n_1571), .B2(n_1573), .Y(n_1569) );
INVx1_ASAP7_75t_L g712 ( .A(n_580), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_641), .C(n_664), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_614), .B(n_636), .Y(n_582) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_585), .A2(n_612), .B1(n_1562), .B2(n_1563), .Y(n_1561) );
INVx3_ASAP7_75t_L g1637 ( .A(n_585), .Y(n_1637) );
AND2x4_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g1277 ( .A(n_586), .Y(n_1277) );
BUFx2_ASAP7_75t_L g1339 ( .A(n_586), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1622 ( .A(n_586), .Y(n_1622) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g603 ( .A(n_587), .Y(n_603) );
BUFx3_ASAP7_75t_L g971 ( .A(n_587), .Y(n_971) );
BUFx3_ASAP7_75t_L g1173 ( .A(n_587), .Y(n_1173) );
AND2x2_ASAP7_75t_L g609 ( .A(n_588), .B(n_600), .Y(n_609) );
AND2x4_ASAP7_75t_L g612 ( .A(n_588), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g942 ( .A(n_588), .B(n_613), .Y(n_942) );
AND2x2_ASAP7_75t_L g980 ( .A(n_588), .B(n_602), .Y(n_980) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_588), .Y(n_1180) );
AOI21xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_597), .B(n_604), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g1305 ( .A1(n_591), .A2(n_775), .B1(n_843), .B2(n_1306), .C1(n_1307), .C2(n_1308), .Y(n_1305) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g1076 ( .A(n_593), .Y(n_1076) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g1333 ( .A(n_594), .Y(n_1333) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g1640 ( .A(n_595), .Y(n_1640) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g970 ( .A(n_599), .Y(n_970) );
INVx1_ASAP7_75t_L g1325 ( .A(n_599), .Y(n_1325) );
INVx2_ASAP7_75t_L g1552 ( .A(n_599), .Y(n_1552) );
INVx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_600), .B(n_605), .Y(n_650) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_600), .Y(n_955) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_602), .B(n_1071), .Y(n_1070) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g1219 ( .A(n_603), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1547 ( .A1(n_604), .A2(n_1548), .B1(n_1551), .B2(n_1553), .C(n_1554), .Y(n_1547) );
AOI21xp5_ASAP7_75t_L g1638 ( .A1(n_604), .A2(n_1639), .B(n_1641), .Y(n_1638) );
INVx1_ASAP7_75t_L g1919 ( .A(n_604), .Y(n_1919) );
INVx1_ASAP7_75t_L g623 ( .A(n_605), .Y(n_623) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_605), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_610), .B2(n_611), .Y(n_606) );
AOI221xp5_ASAP7_75t_SL g1555 ( .A1(n_608), .A2(n_1556), .B1(n_1557), .B2(n_1559), .C(n_1560), .Y(n_1555) );
AOI22xp33_ASAP7_75t_L g1642 ( .A1(n_608), .A2(n_612), .B1(n_1643), .B2(n_1644), .Y(n_1642) );
INVx1_ASAP7_75t_L g1929 ( .A(n_608), .Y(n_1929) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g932 ( .A(n_609), .B(n_933), .Y(n_932) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g1922 ( .A(n_612), .Y(n_1922) );
BUFx6f_ASAP7_75t_L g975 ( .A(n_613), .Y(n_975) );
INVx2_ASAP7_75t_L g1183 ( .A(n_613), .Y(n_1183) );
INVx1_ASAP7_75t_L g1550 ( .A(n_613), .Y(n_1550) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g981 ( .A(n_616), .Y(n_981) );
INVx4_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx3_ASAP7_75t_L g1553 ( .A(n_618), .Y(n_1553) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g1923 ( .A(n_621), .Y(n_1923) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g1224 ( .A(n_622), .Y(n_1224) );
INVx1_ASAP7_75t_L g1288 ( .A(n_623), .Y(n_1288) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .B1(n_629), .B2(n_630), .C(n_631), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_625), .A2(n_721), .B1(n_742), .B2(n_751), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_625), .A2(n_729), .B1(n_736), .B2(n_765), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g830 ( .A1(n_625), .A2(n_807), .B1(n_823), .B2(n_831), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_625), .A2(n_751), .B1(n_1377), .B2(n_1378), .Y(n_1376) );
OAI221xp5_ASAP7_75t_L g1646 ( .A1(n_625), .A2(n_1038), .B1(n_1647), .B2(n_1648), .C(n_1649), .Y(n_1646) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
BUFx3_ASAP7_75t_L g1081 ( .A(n_627), .Y(n_1081) );
BUFx6f_ASAP7_75t_L g1477 ( .A(n_627), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_629), .A2(n_817), .B1(n_821), .B2(n_838), .Y(n_837) );
OAI221xp5_ASAP7_75t_L g1924 ( .A1(n_629), .A2(n_1477), .B1(n_1925), .B2(n_1926), .C(n_1927), .Y(n_1924) );
OAI22xp5_ASAP7_75t_L g1979 ( .A1(n_629), .A2(n_838), .B1(n_1968), .B2(n_1971), .Y(n_1979) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g968 ( .A(n_635), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g1174 ( .A1(n_635), .A2(n_761), .B1(n_1175), .B2(n_1176), .C(n_1177), .Y(n_1174) );
INVx1_ASAP7_75t_L g1217 ( .A(n_635), .Y(n_1217) );
OAI221xp5_ASAP7_75t_L g1278 ( .A1(n_635), .A2(n_761), .B1(n_1041), .B2(n_1279), .C(n_1280), .Y(n_1278) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g982 ( .A(n_638), .Y(n_982) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g1169 ( .A1(n_639), .A2(n_1170), .A3(n_1178), .B(n_1188), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_639), .Y(n_1205) );
OAI31xp33_ASAP7_75t_L g1274 ( .A1(n_639), .A2(n_1275), .A3(n_1281), .B(n_1289), .Y(n_1274) );
BUFx2_ASAP7_75t_L g1564 ( .A(n_639), .Y(n_1564) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI21xp33_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_651), .B(n_652), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g1581 ( .A1(n_642), .A2(n_1582), .B(n_1583), .Y(n_1581) );
AOI21xp5_ASAP7_75t_L g1669 ( .A1(n_642), .A2(n_1670), .B(n_1671), .Y(n_1669) );
INVx8_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g1151 ( .A(n_644), .Y(n_1151) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
BUFx3_ASAP7_75t_L g820 ( .A(n_645), .Y(n_820) );
INVx1_ASAP7_75t_L g704 ( .A(n_646), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_646), .Y(n_707) );
INVx1_ASAP7_75t_L g1125 ( .A(n_647), .Y(n_1125) );
INVx1_ASAP7_75t_L g1068 ( .A(n_648), .Y(n_1068) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
AND2x4_ASAP7_75t_L g695 ( .A(n_649), .B(n_661), .Y(n_695) );
INVx2_ASAP7_75t_L g1544 ( .A(n_653), .Y(n_1544) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
AND2x4_ASAP7_75t_L g1655 ( .A(n_654), .B(n_656), .Y(n_1655) );
INVx2_ASAP7_75t_L g1146 ( .A(n_656), .Y(n_1146) );
INVx5_ASAP7_75t_L g1198 ( .A(n_657), .Y(n_1198) );
INVx3_ASAP7_75t_L g1906 ( .A(n_657), .Y(n_1906) );
OR2x6_ASAP7_75t_L g657 ( .A(n_658), .B(n_663), .Y(n_657) );
NAND2x1p5_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
BUFx3_ASAP7_75t_L g671 ( .A(n_659), .Y(n_671) );
INVx8_ASAP7_75t_L g1112 ( .A(n_659), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_659), .Y(n_1118) );
BUFx3_ASAP7_75t_L g1580 ( .A(n_659), .Y(n_1580) );
AND2x6_ASAP7_75t_L g1106 ( .A(n_661), .B(n_693), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_661), .B(n_700), .Y(n_1108) );
INVx1_ASAP7_75t_L g1115 ( .A(n_661), .Y(n_1115) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_701), .C(n_708), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_690), .Y(n_665) );
AOI33xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .A3(n_673), .B1(n_679), .B2(n_684), .B3(n_687), .Y(n_666) );
BUFx3_ASAP7_75t_L g996 ( .A(n_667), .Y(n_996) );
AOI33xp33_ASAP7_75t_L g1153 ( .A1(n_667), .A2(n_684), .A3(n_1154), .B1(n_1156), .B2(n_1157), .B3(n_1160), .Y(n_1153) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_667), .B(n_1256), .C(n_1257), .Y(n_1255) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
BUFx3_ASAP7_75t_L g1345 ( .A(n_671), .Y(n_1345) );
INVx1_ASAP7_75t_L g1384 ( .A(n_674), .Y(n_1384) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1349 ( .A(n_676), .Y(n_1349) );
INVx5_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx3_ASAP7_75t_L g683 ( .A(n_677), .Y(n_683) );
BUFx3_ASAP7_75t_L g985 ( .A(n_677), .Y(n_985) );
BUFx12f_ASAP7_75t_L g1242 ( .A(n_677), .Y(n_1242) );
INVx1_ASAP7_75t_L g700 ( .A(n_678), .Y(n_700) );
INVx2_ASAP7_75t_L g1021 ( .A(n_680), .Y(n_1021) );
INVx8_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx3_ASAP7_75t_L g735 ( .A(n_681), .Y(n_735) );
INVx5_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx3_ASAP7_75t_L g876 ( .A(n_682), .Y(n_876) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_682), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_682), .A2(n_1155), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
NAND3xp33_ASAP7_75t_L g1265 ( .A(n_684), .B(n_1266), .C(n_1267), .Y(n_1265) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI33xp33_ASAP7_75t_L g804 ( .A1(n_685), .A2(n_805), .A3(n_806), .B1(n_813), .B2(n_818), .B3(n_822), .Y(n_804) );
OAI33xp33_ASAP7_75t_L g1490 ( .A1(n_685), .A2(n_805), .A3(n_1491), .B1(n_1492), .B2(n_1494), .B3(n_1496), .Y(n_1490) );
OAI33xp33_ASAP7_75t_L g1961 ( .A1(n_685), .A2(n_805), .A3(n_1962), .B1(n_1966), .B2(n_1969), .B3(n_1972), .Y(n_1961) );
INVx3_ASAP7_75t_L g1129 ( .A(n_686), .Y(n_1129) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g1232 ( .A(n_689), .Y(n_1232) );
INVx1_ASAP7_75t_L g1258 ( .A(n_689), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_696), .B2(n_697), .Y(n_690) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
NAND2x1_ASAP7_75t_L g946 ( .A(n_693), .B(n_695), .Y(n_946) );
AND2x4_ASAP7_75t_SL g1165 ( .A(n_693), .B(n_695), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1902 ( .A(n_693), .B(n_695), .Y(n_1902) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g697 ( .A(n_695), .B(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g710 ( .A(n_695), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_SL g1167 ( .A(n_695), .B(n_698), .Y(n_1167) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_697), .A2(n_945), .B1(n_947), .B2(n_948), .C(n_949), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g1584 ( .A1(n_697), .A2(n_710), .B1(n_1165), .B2(n_1554), .C(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1659 ( .A(n_697), .Y(n_1659) );
AOI22xp33_ASAP7_75t_L g1900 ( .A1(n_697), .A2(n_1901), .B1(n_1902), .B2(n_1903), .Y(n_1900) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g938 ( .A(n_704), .B(n_939), .Y(n_938) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_706), .B(n_1162), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_706), .B(n_1260), .Y(n_1259) );
INVx2_ASAP7_75t_L g1947 ( .A(n_706), .Y(n_1947) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_707), .B(n_1149), .Y(n_1148) );
AND2x4_ASAP7_75t_L g1588 ( .A(n_707), .B(n_1149), .Y(n_1588) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
NAND5xp2_ASAP7_75t_L g1899 ( .A(n_709), .B(n_1900), .C(n_1904), .D(n_1907), .E(n_1908), .Y(n_1899) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g1164 ( .A1(n_710), .A2(n_1165), .B1(n_1166), .B2(n_1167), .C(n_1168), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_710), .A2(n_1165), .B1(n_1167), .B2(n_1270), .C(n_1271), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g1671 ( .A(n_710), .Y(n_1671) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_799), .B2(n_800), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_766), .C(n_784), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_747), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .A3(n_726), .B1(n_733), .B2(n_738), .B3(n_739), .Y(n_718) );
OAI33xp33_ASAP7_75t_L g1411 ( .A1(n_719), .A2(n_738), .A3(n_1412), .B1(n_1416), .B2(n_1419), .B3(n_1423), .Y(n_1411) );
OAI22xp33_ASAP7_75t_L g1380 ( .A1(n_722), .A2(n_1362), .B1(n_1372), .B2(n_1381), .Y(n_1380) );
OAI22xp33_ASAP7_75t_L g1385 ( .A1(n_722), .A2(n_1365), .B1(n_1375), .B2(n_1386), .Y(n_1385) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g741 ( .A(n_724), .Y(n_741) );
INVxp67_ASAP7_75t_SL g1572 ( .A(n_724), .Y(n_1572) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_725), .A2(n_746), .B1(n_758), .B2(n_761), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_727), .A2(n_734), .B1(n_754), .B2(n_756), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g1616 ( .A1(n_728), .A2(n_889), .B1(n_1617), .B2(n_1618), .Y(n_1616) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_730), .A2(n_1369), .B1(n_1378), .B2(n_1384), .Y(n_1383) );
INVx3_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g878 ( .A(n_732), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g1416 ( .A1(n_735), .A2(n_737), .B1(n_1417), .B2(n_1418), .Y(n_1416) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_735), .A2(n_737), .B1(n_1567), .B2(n_1568), .Y(n_1566) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_737), .A2(n_1131), .B1(n_1133), .B2(n_1134), .Y(n_1130) );
OAI221xp5_ASAP7_75t_L g1227 ( .A1(n_737), .A2(n_1228), .B1(n_1229), .B2(n_1230), .C(n_1231), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1233 ( .A1(n_737), .A2(n_1215), .B1(n_1234), .B2(n_1235), .C(n_1236), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_737), .A2(n_1234), .B1(n_1367), .B2(n_1377), .Y(n_1382) );
OAI33xp33_ASAP7_75t_L g1604 ( .A1(n_738), .A2(n_867), .A3(n_1605), .B1(n_1609), .B2(n_1613), .B3(n_1616), .Y(n_1604) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_742), .B1(n_743), .B2(n_746), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g1381 ( .A(n_744), .Y(n_1381) );
INVxp67_ASAP7_75t_SL g1975 ( .A(n_744), .Y(n_1975) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g812 ( .A(n_745), .Y(n_812) );
OAI33xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .A3(n_753), .B1(n_757), .B2(n_762), .B3(n_764), .Y(n_747) );
OAI33xp33_ASAP7_75t_L g1360 ( .A1(n_748), .A2(n_762), .A3(n_1361), .B1(n_1366), .B2(n_1371), .B3(n_1376), .Y(n_1360) );
OAI33xp33_ASAP7_75t_L g1427 ( .A1(n_748), .A2(n_902), .A3(n_1428), .B1(n_1431), .B2(n_1432), .B3(n_1435), .Y(n_1427) );
OAI22xp5_ASAP7_75t_L g1619 ( .A1(n_748), .A2(n_762), .B1(n_1620), .B2(n_1623), .Y(n_1619) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g1487 ( .A1(n_751), .A2(n_838), .B1(n_1488), .B2(n_1489), .Y(n_1487) );
INVx5_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx6_ASAP7_75t_L g1437 ( .A(n_752), .Y(n_1437) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_754), .A2(n_1088), .B1(n_1089), .B2(n_1090), .C(n_1091), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_754), .A2(n_1372), .B1(n_1373), .B2(n_1375), .Y(n_1371) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
HB1xp67_ASAP7_75t_L g1523 ( .A(n_756), .Y(n_1523) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_758), .A2(n_1373), .B1(n_1417), .B2(n_1420), .Y(n_1431) );
INVx4_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g1041 ( .A(n_760), .Y(n_1041) );
INVx2_ASAP7_75t_L g1177 ( .A(n_760), .Y(n_1177) );
OAI211xp5_ASAP7_75t_L g972 ( .A1(n_761), .A2(n_973), .B(n_974), .C(n_977), .Y(n_972) );
OAI21xp5_ASAP7_75t_L g1086 ( .A1(n_762), .A2(n_1087), .B(n_1092), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g902 ( .A(n_763), .Y(n_902) );
NAND3xp33_ASAP7_75t_L g1331 ( .A(n_763), .B(n_1332), .C(n_1338), .Y(n_1331) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_772), .A2(n_814), .B1(n_819), .B2(n_833), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_772), .A2(n_810), .B1(n_825), .B2(n_833), .Y(n_834) );
BUFx2_ASAP7_75t_L g917 ( .A(n_772), .Y(n_917) );
BUFx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_773), .B(n_1072), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_773), .B(n_1187), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_773), .B(n_1287), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1374 ( .A(n_773), .Y(n_1374) );
BUFx2_ASAP7_75t_SL g1434 ( .A(n_773), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B1(n_777), .B2(n_779), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_775), .A2(n_842), .B1(n_843), .B2(n_844), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1985 ( .A1(n_775), .A2(n_843), .B1(n_1986), .B2(n_1987), .Y(n_1985) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g843 ( .A(n_778), .Y(n_843) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g1011 ( .A(n_783), .Y(n_1011) );
INVx2_ASAP7_75t_L g1406 ( .A(n_783), .Y(n_1406) );
OAI31xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_787), .A3(n_793), .B(n_798), .Y(n_784) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g853 ( .A(n_790), .Y(n_853) );
INVx2_ASAP7_75t_L g988 ( .A(n_790), .Y(n_988) );
INVx1_ASAP7_75t_L g1386 ( .A(n_790), .Y(n_1386) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g1056 ( .A(n_795), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1631 ( .A1(n_795), .A2(n_858), .B1(n_1596), .B2(n_1597), .Y(n_1631) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OAI31xp33_ASAP7_75t_L g1312 ( .A1(n_798), .A2(n_1313), .A3(n_1315), .B(n_1317), .Y(n_1312) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_839), .C(n_848), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_826), .Y(n_803) );
OAI22xp5_ASAP7_75t_SL g1660 ( .A1(n_805), .A2(n_1027), .B1(n_1661), .B2(n_1665), .Y(n_1660) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_810), .B2(n_811), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_808), .A2(n_973), .B1(n_987), .B2(n_988), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1962 ( .A1(n_808), .A2(n_1963), .B1(n_1964), .B2(n_1965), .Y(n_1962) );
BUFx4f_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
OAI22xp33_ASAP7_75t_L g822 ( .A1(n_809), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g1491 ( .A1(n_809), .A2(n_995), .B1(n_1476), .B2(n_1485), .Y(n_1491) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1965 ( .A(n_812), .Y(n_1965) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_815), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_818) );
INVx2_ASAP7_75t_L g1342 ( .A(n_815), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_815), .A2(n_1481), .B1(n_1488), .B2(n_1493), .Y(n_1492) );
OAI22xp5_ASAP7_75t_L g1966 ( .A1(n_815), .A2(n_1493), .B1(n_1967), .B2(n_1968), .Y(n_1966) );
BUFx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g881 ( .A(n_816), .Y(n_881) );
INVx3_ASAP7_75t_L g939 ( .A(n_816), .Y(n_939) );
BUFx2_ASAP7_75t_L g1509 ( .A(n_816), .Y(n_1509) );
INVx1_ASAP7_75t_L g884 ( .A(n_824), .Y(n_884) );
HB1xp67_ASAP7_75t_L g1516 ( .A(n_824), .Y(n_1516) );
OAI33xp33_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_830), .A3(n_832), .B1(n_834), .B2(n_835), .B3(n_837), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_SL g1330 ( .A(n_829), .Y(n_1330) );
INVx2_ASAP7_75t_L g1039 ( .A(n_831), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_831), .A2(n_1193), .B1(n_1194), .B2(n_1195), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g1475 ( .A1(n_831), .A2(n_1476), .B1(n_1477), .B2(n_1478), .Y(n_1475) );
OAI22xp33_ASAP7_75t_L g1978 ( .A1(n_831), .A2(n_1477), .B1(n_1963), .B2(n_1973), .Y(n_1978) );
OAI22xp5_ASAP7_75t_SL g1480 ( .A1(n_833), .A2(n_957), .B1(n_1481), .B2(n_1482), .Y(n_1480) );
OAI22xp5_ASAP7_75t_L g1977 ( .A1(n_833), .A2(n_1370), .B1(n_1967), .B2(n_1970), .Y(n_1977) );
OAI33xp33_ASAP7_75t_L g1474 ( .A1(n_835), .A2(n_1475), .A3(n_1479), .B1(n_1480), .B2(n_1483), .B3(n_1487), .Y(n_1474) );
OAI33xp33_ASAP7_75t_L g1976 ( .A1(n_835), .A2(n_892), .A3(n_1977), .B1(n_1978), .B2(n_1979), .B3(n_1980), .Y(n_1976) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OAI31xp33_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_851), .A3(n_856), .B(n_859), .Y(n_848) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_853), .A2(n_1084), .B1(n_1090), .B2(n_1128), .C(n_1129), .Y(n_1127) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI31xp33_ASAP7_75t_L g1467 ( .A1(n_859), .A2(n_1468), .A3(n_1469), .B(n_1472), .Y(n_1467) );
OAI31xp33_ASAP7_75t_SL g1989 ( .A1(n_859), .A2(n_1990), .A3(n_1991), .B(n_1992), .Y(n_1989) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
XNOR2x1_ASAP7_75t_L g861 ( .A(n_862), .B(n_1059), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_923), .Y(n_862) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_903), .C(n_910), .Y(n_864) );
NOR2xp33_ASAP7_75t_SL g865 ( .A(n_866), .B(n_891), .Y(n_865) );
OAI33xp33_ASAP7_75t_L g1013 ( .A1(n_867), .A2(n_1014), .A3(n_1019), .B1(n_1024), .B2(n_1027), .B3(n_1030), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1226 ( .A1(n_867), .A2(n_1227), .B1(n_1233), .B2(n_1238), .Y(n_1226) );
OAI33xp33_ASAP7_75t_L g1503 ( .A1(n_867), .A2(n_1027), .A3(n_1504), .B1(n_1507), .B2(n_1511), .B3(n_1514), .Y(n_1503) );
BUFx3_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OAI22xp33_ASAP7_75t_SL g872 ( .A1(n_873), .A2(n_874), .B1(n_877), .B2(n_878), .Y(n_872) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_875), .A2(n_1101), .B1(n_1102), .B2(n_1118), .Y(n_1117) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_882), .B1(n_883), .B2(n_885), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1421 ( .A(n_881), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_883), .A2(n_1015), .B1(n_1016), .B2(n_1018), .Y(n_1014) );
INVx2_ASAP7_75t_SL g883 ( .A(n_884), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g1507 ( .A1(n_889), .A2(n_1508), .B1(n_1509), .B2(n_1510), .Y(n_1507) );
OAI33xp33_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .A3(n_894), .B1(n_896), .B2(n_897), .B3(n_902), .Y(n_891) );
OAI221xp5_ASAP7_75t_SL g1620 ( .A1(n_895), .A2(n_1177), .B1(n_1610), .B2(n_1617), .C(n_1621), .Y(n_1620) );
OAI221xp5_ASAP7_75t_SL g1623 ( .A1(n_895), .A2(n_1177), .B1(n_1607), .B2(n_1615), .C(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI31xp33_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_912), .A3(n_916), .B(n_922), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1595 ( .A1(n_914), .A2(n_1301), .B1(n_1596), .B2(n_1597), .Y(n_1595) );
INVx2_ASAP7_75t_SL g914 ( .A(n_915), .Y(n_914) );
OAI31xp33_ASAP7_75t_L g1438 ( .A1(n_922), .A2(n_1439), .A3(n_1440), .B(n_1444), .Y(n_1438) );
OAI31xp33_ASAP7_75t_L g1460 ( .A1(n_922), .A2(n_1461), .A3(n_1465), .B(n_1466), .Y(n_1460) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AO22x2_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_997), .B1(n_998), .B2(n_1058), .Y(n_924) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_925), .Y(n_1058) );
XNOR2x1_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
NOR2x1_ASAP7_75t_L g927 ( .A(n_928), .B(n_943), .Y(n_927) );
INVxp67_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_934), .Y(n_930) );
INVx3_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_932), .A2(n_941), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
AND2x4_ASAP7_75t_L g941 ( .A(n_933), .B(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND2x1_ASAP7_75t_L g936 ( .A(n_937), .B(n_940), .Y(n_936) );
INVx2_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_L g1234 ( .A(n_939), .Y(n_1234) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
NAND3xp33_ASAP7_75t_SL g943 ( .A(n_944), .B(n_950), .C(n_983), .Y(n_943) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_947), .A2(n_959), .B1(n_960), .B2(n_961), .Y(n_958) );
OAI21xp5_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_978), .B(n_982), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_964), .C(n_972), .Y(n_951) );
A2O1A1Ixp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B(n_956), .C(n_963), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_SL g1220 ( .A1(n_954), .A2(n_963), .B(n_1221), .C(n_1222), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx3_ASAP7_75t_L g1172 ( .A(n_955), .Y(n_1172) );
A2O1A1Ixp33_ASAP7_75t_L g1185 ( .A1(n_955), .A2(n_963), .B(n_1152), .C(n_1186), .Y(n_1185) );
A2O1A1Ixp33_ASAP7_75t_L g1285 ( .A1(n_955), .A2(n_1264), .B(n_1286), .C(n_1288), .Y(n_1285) );
NAND2xp5_ASAP7_75t_SL g956 ( .A(n_957), .B(n_958), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_959), .A2(n_961), .B1(n_1262), .B2(n_1270), .Y(n_1287) );
INVx1_ASAP7_75t_L g1225 ( .A(n_961), .Y(n_1225) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
BUFx2_ASAP7_75t_L g1322 ( .A(n_967), .Y(n_1322) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_971), .Y(n_1323) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_985), .A2(n_1120), .B1(n_1121), .B2(n_1122), .Y(n_1119) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g1511 ( .A1(n_991), .A2(n_1023), .B1(n_1512), .B2(n_1513), .Y(n_1511) );
OAI211xp5_ASAP7_75t_L g1135 ( .A1(n_995), .A2(n_1088), .B(n_1136), .C(n_1138), .Y(n_1135) );
NAND3xp33_ASAP7_75t_L g1340 ( .A(n_996), .B(n_1341), .C(n_1344), .Y(n_1340) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
NAND3xp33_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1012), .C(n_1044), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_1004), .A2(n_1051), .B1(n_1053), .B2(n_1054), .Y(n_1050) );
NOR2xp33_ASAP7_75t_SL g1012 ( .A(n_1013), .B(n_1033), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_1015), .A2(n_1031), .B1(n_1035), .B2(n_1038), .Y(n_1034) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_1022), .A2(n_1026), .B1(n_1035), .B2(n_1038), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1665 ( .A1(n_1023), .A2(n_1421), .B1(n_1666), .B2(n_1667), .C(n_1668), .Y(n_1665) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1942 ( .A(n_1029), .Y(n_1942) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_SL g1036 ( .A(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
OAI22xp33_ASAP7_75t_SL g1522 ( .A1(n_1041), .A2(n_1506), .B1(n_1517), .B2(n_1523), .Y(n_1522) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_1047), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1626 ( .A(n_1049), .B(n_1627), .C(n_1631), .Y(n_1626) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_1051), .A2(n_1053), .B1(n_1307), .B2(n_1308), .Y(n_1316) );
BUFx3_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
BUFx3_ASAP7_75t_L g1451 ( .A(n_1052), .Y(n_1451) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_1053), .A2(n_1442), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
AOI222xp33_ASAP7_75t_L g1627 ( .A1(n_1053), .A2(n_1451), .B1(n_1599), .B2(n_1600), .C1(n_1601), .C2(n_1628), .Y(n_1627) );
XNOR2x1_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1295), .Y(n_1059) );
OA22x2_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1062), .B1(n_1200), .B2(n_1294), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
XOR2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1142), .Y(n_1062) );
XNOR2x1_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
NAND4xp75_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1074), .C(n_1100), .D(n_1103), .Y(n_1065) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
AOI211x1_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1085), .B(n_1086), .C(n_1096), .Y(n_1074) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
AOI221xp5_ASAP7_75t_L g1181 ( .A1(n_1078), .A2(n_1162), .B1(n_1168), .B2(n_1182), .C(n_1184), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_1078), .A2(n_1182), .B1(n_1260), .B2(n_1271), .C(n_1283), .Y(n_1282) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1082), .B2(n_1084), .Y(n_1079) );
BUFx6f_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
OAI211xp5_ASAP7_75t_SL g1210 ( .A1(n_1089), .A2(n_1211), .B(n_1212), .C(n_1213), .Y(n_1210) );
OAI211xp5_ASAP7_75t_SL g1214 ( .A1(n_1089), .A2(n_1215), .B(n_1216), .C(n_1218), .Y(n_1214) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
NAND2x2_ASAP7_75t_L g1097 ( .A(n_1094), .B(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_1099), .Y(n_1098) );
OAI31xp67_ASAP7_75t_L g1103 ( .A1(n_1104), .A2(n_1116), .A3(n_1126), .B(n_1140), .Y(n_1103) );
INVx4_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
A2O1A1Ixp33_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1111), .B(n_1113), .C(n_1114), .Y(n_1109) );
CKINVDCx5p33_ASAP7_75t_R g1111 ( .A(n_1112), .Y(n_1111) );
INVx3_ASAP7_75t_L g1139 ( .A(n_1112), .Y(n_1139) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1112), .Y(n_1149) );
INVx8_ASAP7_75t_L g1155 ( .A(n_1112), .Y(n_1155) );
INVx2_ASAP7_75t_L g1946 ( .A(n_1112), .Y(n_1946) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_1113), .A2(n_1221), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
AOI21xp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1119), .B(n_1123), .Y(n_1116) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
OAI21xp5_ASAP7_75t_SL g1126 ( .A1(n_1127), .A2(n_1130), .B(n_1135), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_1128), .A2(n_1413), .B1(n_1414), .B2(n_1415), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g1423 ( .A1(n_1128), .A2(n_1424), .B1(n_1425), .B2(n_1426), .Y(n_1423) );
OAI22xp33_ASAP7_75t_L g1605 ( .A1(n_1128), .A2(n_1606), .B1(n_1607), .B2(n_1608), .Y(n_1605) );
OAI22xp33_ASAP7_75t_L g1613 ( .A1(n_1128), .A2(n_1516), .B1(n_1614), .B2(n_1615), .Y(n_1613) );
OAI22xp33_ASAP7_75t_L g1972 ( .A1(n_1128), .A2(n_1973), .B1(n_1974), .B2(n_1975), .Y(n_1972) );
OAI221xp5_ASAP7_75t_L g1574 ( .A1(n_1131), .A2(n_1493), .B1(n_1575), .B2(n_1576), .C(n_1577), .Y(n_1574) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1228 ( .A(n_1132), .Y(n_1228) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1140), .Y(n_1651) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1141), .Y(n_1930) );
XNOR2x1_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1199), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1163), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1153), .C(n_1161), .Y(n_1144) );
AOI222xp33_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1147), .B1(n_1148), .B2(n_1150), .C1(n_1151), .C2(n_1152), .Y(n_1145) );
AOI222xp33_ASAP7_75t_L g1261 ( .A1(n_1146), .A2(n_1148), .B1(n_1151), .B2(n_1262), .C1(n_1263), .C2(n_1264), .Y(n_1261) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
NAND3xp33_ASAP7_75t_SL g1163 ( .A(n_1164), .B(n_1169), .C(n_1196), .Y(n_1163) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1558 ( .A(n_1172), .Y(n_1558) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_1177), .A2(n_1508), .B1(n_1512), .B2(n_1521), .Y(n_1520) );
OAI21xp33_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1181), .B(n_1185), .Y(n_1178) );
OAI21xp5_ASAP7_75t_SL g1281 ( .A1(n_1179), .A2(n_1282), .B(n_1285), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
OAI21xp5_ASAP7_75t_L g1207 ( .A1(n_1180), .A2(n_1208), .B(n_1209), .Y(n_1207) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1198), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1198), .B(n_1273), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1198), .B(n_1563), .Y(n_1586) );
XNOR2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1252), .Y(n_1200) );
XOR2xp5_ASAP7_75t_L g1294 ( .A(n_1201), .B(n_1252), .Y(n_1294) );
XNOR2x1_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1239), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1206), .B(n_1226), .Y(n_1204) );
NAND4xp25_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1210), .C(n_1214), .D(n_1220), .Y(n_1206) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
HB1xp67_ASAP7_75t_L g1343 ( .A(n_1237), .Y(n_1343) );
XNOR2x1_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1293), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1268), .Y(n_1253) );
NAND4xp25_ASAP7_75t_SL g1254 ( .A(n_1255), .B(n_1259), .C(n_1261), .D(n_1265), .Y(n_1254) );
NAND3xp33_ASAP7_75t_SL g1268 ( .A(n_1269), .B(n_1272), .C(n_1274), .Y(n_1268) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1297), .Y(n_1351) );
NAND3xp33_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1312), .C(n_1319), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1309), .B(n_1311), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B1(n_1303), .B2(n_1304), .Y(n_1300) );
OAI21xp5_ASAP7_75t_L g1593 ( .A1(n_1311), .A2(n_1594), .B(n_1602), .Y(n_1593) );
OAI31xp33_ASAP7_75t_L g1981 ( .A1(n_1311), .A2(n_1982), .A3(n_1983), .B(n_1988), .Y(n_1981) );
AND4x1_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1331), .C(n_1340), .D(n_1346), .Y(n_1319) );
NAND3xp33_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1324), .C(n_1330), .Y(n_1320) );
INVx2_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
BUFx2_ASAP7_75t_L g1337 ( .A(n_1329), .Y(n_1337) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
XNOR2xp5_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1456), .Y(n_1354) );
OAI22xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B1(n_1407), .B2(n_1455), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND3xp33_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1387), .C(n_1397), .Y(n_1358) );
NOR2xp33_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1379), .Y(n_1359) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_1367), .A2(n_1368), .B1(n_1369), .B2(n_1370), .Y(n_1366) );
INVx5_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
OAI31xp33_ASAP7_75t_L g1387 ( .A1(n_1388), .A2(n_1389), .A3(n_1393), .B(n_1396), .Y(n_1387) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx2_ASAP7_75t_L g1984 ( .A(n_1401), .Y(n_1984) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1407), .Y(n_1455) );
BUFx2_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
AND3x1_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1438), .C(n_1445), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1427), .Y(n_1410) );
OAI22xp33_ASAP7_75t_L g1428 ( .A1(n_1413), .A2(n_1424), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_1414), .A2(n_1425), .B1(n_1433), .B2(n_1434), .Y(n_1432) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_1418), .A2(n_1422), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
AOI22xp5_ASAP7_75t_L g1456 ( .A1(n_1457), .A2(n_1458), .B1(n_1497), .B2(n_1498), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
NAND3xp33_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1467), .C(n_1473), .Y(n_1459) );
NOR2xp33_ASAP7_75t_SL g1473 ( .A(n_1474), .B(n_1490), .Y(n_1473) );
OAI221xp5_ASAP7_75t_L g1913 ( .A1(n_1477), .A2(n_1914), .B1(n_1915), .B2(n_1916), .C(n_1917), .Y(n_1913) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
AO22x2_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1590), .B1(n_1672), .B2(n_1673), .Y(n_1498) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1499), .Y(n_1672) );
XNOR2xp5_ASAP7_75t_L g1499 ( .A(n_1500), .B(n_1541), .Y(n_1499) );
NAND3xp33_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1525), .C(n_1534), .Y(n_1501) );
NOR2xp33_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1518), .Y(n_1502) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
XNOR2xp5_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1589), .Y(n_1541) );
NAND2xp5_ASAP7_75t_SL g1542 ( .A(n_1543), .B(n_1581), .Y(n_1542) );
AOI221xp5_ASAP7_75t_L g1543 ( .A1(n_1544), .A2(n_1545), .B1(n_1546), .B2(n_1564), .C(n_1565), .Y(n_1543) );
AOI21xp5_ASAP7_75t_SL g1931 ( .A1(n_1544), .A2(n_1932), .B(n_1933), .Y(n_1931) );
NAND3xp33_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1555), .C(n_1561), .Y(n_1546) );
INVx2_ASAP7_75t_SL g1549 ( .A(n_1550), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1559), .B(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
BUFx2_ASAP7_75t_L g1663 ( .A(n_1580), .Y(n_1663) );
NAND3xp33_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1586), .C(n_1587), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1908 ( .A(n_1588), .B(n_1909), .Y(n_1908) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1590), .Y(n_1673) );
XNOR2x1_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1634), .Y(n_1590) );
XOR2x2_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1633), .Y(n_1591) );
NAND3x1_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1603), .C(n_1625), .Y(n_1592) );
NOR2x1_ASAP7_75t_L g1603 ( .A(n_1604), .B(n_1619), .Y(n_1603) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
O2A1O1Ixp5_ASAP7_75t_L g1635 ( .A1(n_1636), .A2(n_1645), .B(n_1651), .C(n_1652), .Y(n_1635) );
OAI21xp5_ASAP7_75t_L g1661 ( .A1(n_1647), .A2(n_1662), .B(n_1664), .Y(n_1661) );
NAND3xp33_ASAP7_75t_L g1652 ( .A(n_1653), .B(n_1657), .C(n_1669), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1653 ( .A(n_1654), .B(n_1656), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1660), .Y(n_1657) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
OAI221xp5_ASAP7_75t_L g1675 ( .A1(n_1676), .A2(n_1893), .B1(n_1896), .B2(n_1949), .C(n_1952), .Y(n_1675) );
AOI211xp5_ASAP7_75t_L g1676 ( .A1(n_1677), .A2(n_1693), .B(n_1775), .C(n_1887), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1827 ( .A(n_1677), .B(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1677), .Y(n_1878) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
NAND3xp33_ASAP7_75t_L g1869 ( .A(n_1678), .B(n_1731), .C(n_1813), .Y(n_1869) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_1678), .B(n_1829), .Y(n_1886) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
AOI32xp33_ASAP7_75t_L g1795 ( .A1(n_1679), .A2(n_1723), .A3(n_1765), .B1(n_1796), .B2(n_1798), .Y(n_1795) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1679), .Y(n_1799) );
NOR2xp33_ASAP7_75t_L g1810 ( .A(n_1679), .B(n_1705), .Y(n_1810) );
AOI211xp5_ASAP7_75t_L g1811 ( .A1(n_1679), .A2(n_1812), .B(n_1813), .C(n_1817), .Y(n_1811) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1687), .Y(n_1679) );
INVx2_ASAP7_75t_L g1895 ( .A(n_1681), .Y(n_1895) );
AND2x6_ASAP7_75t_L g1681 ( .A(n_1682), .B(n_1683), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1682), .B(n_1686), .Y(n_1685) );
AND2x4_ASAP7_75t_L g1688 ( .A(n_1682), .B(n_1689), .Y(n_1688) );
AND2x6_ASAP7_75t_L g1691 ( .A(n_1682), .B(n_1692), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1682), .B(n_1686), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1682), .B(n_1686), .Y(n_1721) );
OAI21xp5_ASAP7_75t_L g1996 ( .A1(n_1683), .A2(n_1997), .B(n_1998), .Y(n_1996) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1684), .B(n_1690), .Y(n_1689) );
NAND5xp2_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1753), .C(n_1763), .D(n_1768), .E(n_1771), .Y(n_1693) );
AOI221xp5_ASAP7_75t_SL g1694 ( .A1(n_1695), .A2(n_1709), .B1(n_1716), .B2(n_1731), .C(n_1733), .Y(n_1694) );
O2A1O1Ixp33_ASAP7_75t_L g1854 ( .A1(n_1695), .A2(n_1797), .B(n_1855), .C(n_1857), .Y(n_1854) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
OR2x2_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1701), .Y(n_1696) );
NOR3xp33_ASAP7_75t_L g1838 ( .A(n_1697), .B(n_1805), .C(n_1839), .Y(n_1838) );
AND2x2_ASAP7_75t_L g1842 ( .A(n_1697), .B(n_1705), .Y(n_1842) );
OAI31xp33_ASAP7_75t_L g1873 ( .A1(n_1697), .A2(n_1752), .A3(n_1874), .B(n_1876), .Y(n_1873) );
INVx3_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1698), .B(n_1705), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1698), .B(n_1736), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1698), .B(n_1743), .Y(n_1742) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1698), .B(n_1755), .Y(n_1754) );
INVx3_ASAP7_75t_L g1829 ( .A(n_1698), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1835 ( .A(n_1698), .B(n_1817), .Y(n_1835) );
OR2x2_ASAP7_75t_L g1847 ( .A(n_1698), .B(n_1705), .Y(n_1847) );
AND2x2_ASAP7_75t_L g1850 ( .A(n_1698), .B(n_1799), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1872 ( .A(n_1698), .B(n_1860), .Y(n_1872) );
AND2x4_ASAP7_75t_SL g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1701), .Y(n_1787) );
OR2x2_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1705), .Y(n_1701) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1702), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1702), .B(n_1705), .Y(n_1743) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1702), .Y(n_1757) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1702), .Y(n_1812) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1704), .Y(n_1702) );
OR2x2_ASAP7_75t_L g1756 ( .A(n_1705), .B(n_1757), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1708), .Y(n_1705) );
AND2x4_ASAP7_75t_L g1765 ( .A(n_1706), .B(n_1708), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1709), .B(n_1719), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1709), .B(n_1770), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1709), .B(n_1718), .Y(n_1783) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1709), .Y(n_1875) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1713), .Y(n_1709) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1710), .Y(n_1726) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1710), .Y(n_1866) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1712), .Y(n_1710) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1713), .B(n_1726), .Y(n_1725) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1713), .Y(n_1740) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1713), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1713), .B(n_1726), .Y(n_1761) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1714), .B(n_1715), .Y(n_1713) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
AOI221xp5_ASAP7_75t_SL g1887 ( .A1(n_1717), .A2(n_1764), .B1(n_1787), .B2(n_1888), .C(n_1892), .Y(n_1887) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1718), .B(n_1723), .Y(n_1717) );
AND2x2_ASAP7_75t_L g1797 ( .A(n_1718), .B(n_1724), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1802 ( .A(n_1718), .B(n_1758), .Y(n_1802) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1718), .B(n_1816), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1821 ( .A(n_1718), .B(n_1748), .Y(n_1821) );
AND2x2_ASAP7_75t_L g1882 ( .A(n_1718), .B(n_1866), .Y(n_1882) );
CKINVDCx5p33_ASAP7_75t_R g1718 ( .A(n_1719), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1719), .B(n_1739), .Y(n_1738) );
NOR2xp33_ASAP7_75t_L g1767 ( .A(n_1719), .B(n_1728), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1770 ( .A(n_1719), .B(n_1728), .Y(n_1770) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1719), .B(n_1749), .Y(n_1772) );
OR2x2_ASAP7_75t_L g1856 ( .A(n_1719), .B(n_1740), .Y(n_1856) );
NAND2xp5_ASAP7_75t_L g1865 ( .A(n_1719), .B(n_1866), .Y(n_1865) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1720), .B(n_1722), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1720), .B(n_1722), .Y(n_1786) );
NAND2xp5_ASAP7_75t_SL g1723 ( .A(n_1724), .B(n_1727), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1724), .B(n_1786), .Y(n_1785) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
NOR2xp33_ASAP7_75t_L g1758 ( .A(n_1725), .B(n_1747), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1726), .B(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1726), .Y(n_1816) );
OAI322xp33_ASAP7_75t_L g1733 ( .A1(n_1727), .A2(n_1734), .A3(n_1737), .B1(n_1741), .B2(n_1744), .C1(n_1750), .C2(n_1752), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1750 ( .A(n_1727), .B(n_1751), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1781 ( .A(n_1727), .B(n_1782), .Y(n_1781) );
INVx2_ASAP7_75t_L g1826 ( .A(n_1727), .Y(n_1826) );
NAND2xp5_ASAP7_75t_L g1837 ( .A(n_1727), .B(n_1772), .Y(n_1837) );
INVx2_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx3_ASAP7_75t_L g1747 ( .A(n_1728), .Y(n_1747) );
OR2x2_ASAP7_75t_L g1805 ( .A(n_1728), .B(n_1757), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1730), .Y(n_1728) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
NOR2xp33_ASAP7_75t_L g1857 ( .A(n_1732), .B(n_1858), .Y(n_1857) );
A2O1A1Ixp33_ASAP7_75t_SL g1830 ( .A1(n_1734), .A2(n_1831), .B(n_1832), .C(n_1834), .Y(n_1830) );
OAI221xp5_ASAP7_75t_L g1870 ( .A1(n_1734), .A2(n_1766), .B1(n_1852), .B2(n_1871), .C(n_1873), .Y(n_1870) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1736), .Y(n_1779) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1736), .B(n_1766), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1801 ( .A(n_1736), .B(n_1802), .Y(n_1801) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1736), .Y(n_1824) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
OAI22xp5_ASAP7_75t_SL g1848 ( .A1(n_1739), .A2(n_1849), .B1(n_1851), .B2(n_1853), .Y(n_1848) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
CKINVDCx14_ASAP7_75t_R g1752 ( .A(n_1743), .Y(n_1752) );
AOI22xp5_ASAP7_75t_L g1818 ( .A1(n_1743), .A2(n_1819), .B1(n_1824), .B2(n_1825), .Y(n_1818) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
AOI321xp33_ASAP7_75t_L g1877 ( .A1(n_1745), .A2(n_1751), .A3(n_1846), .B1(n_1878), .B2(n_1879), .C(n_1880), .Y(n_1877) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1746), .B(n_1748), .Y(n_1745) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1746), .B(n_1761), .Y(n_1808) );
AOI21xp33_ASAP7_75t_L g1879 ( .A1(n_1746), .A2(n_1756), .B(n_1828), .Y(n_1879) );
AND2x2_ASAP7_75t_L g1884 ( .A(n_1746), .B(n_1779), .Y(n_1884) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
NAND2xp5_ASAP7_75t_L g1762 ( .A(n_1747), .B(n_1755), .Y(n_1762) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1747), .B(n_1757), .Y(n_1774) );
NAND2xp5_ASAP7_75t_L g1814 ( .A(n_1747), .B(n_1815), .Y(n_1814) );
AND2x2_ASAP7_75t_L g1823 ( .A(n_1747), .B(n_1761), .Y(n_1823) );
NOR2xp33_ASAP7_75t_L g1855 ( .A(n_1747), .B(n_1856), .Y(n_1855) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1748), .B(n_1786), .Y(n_1794) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1748), .Y(n_1839) );
AND2x2_ASAP7_75t_L g1852 ( .A(n_1748), .B(n_1767), .Y(n_1852) );
AOI211xp5_ASAP7_75t_L g1803 ( .A1(n_1751), .A2(n_1804), .B(n_1806), .C(n_1809), .Y(n_1803) );
NAND2xp5_ASAP7_75t_L g1892 ( .A(n_1751), .B(n_1886), .Y(n_1892) );
AOI21xp5_ASAP7_75t_L g1753 ( .A1(n_1754), .A2(n_1758), .B(n_1759), .Y(n_1753) );
INVx2_ASAP7_75t_SL g1755 ( .A(n_1756), .Y(n_1755) );
OAI22xp5_ASAP7_75t_L g1888 ( .A1(n_1756), .A2(n_1817), .B1(n_1889), .B2(n_1891), .Y(n_1888) );
AND2x2_ASAP7_75t_L g1764 ( .A(n_1757), .B(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1758), .Y(n_1831) );
NOR2xp33_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1762), .Y(n_1759) );
OR2x2_ASAP7_75t_L g1792 ( .A(n_1760), .B(n_1786), .Y(n_1792) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1761), .B(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1845 ( .A(n_1761), .B(n_1770), .Y(n_1845) );
AOI211xp5_ASAP7_75t_L g1864 ( .A1(n_1762), .A2(n_1828), .B(n_1865), .C(n_1867), .Y(n_1864) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1764), .B(n_1766), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1768 ( .A(n_1764), .B(n_1769), .Y(n_1768) );
AOI21xp5_ASAP7_75t_L g1790 ( .A1(n_1764), .A2(n_1791), .B(n_1795), .Y(n_1790) );
NAND3xp33_ASAP7_75t_L g1849 ( .A(n_1764), .B(n_1826), .C(n_1850), .Y(n_1849) );
NOR2xp33_ASAP7_75t_L g1798 ( .A(n_1765), .B(n_1799), .Y(n_1798) );
INVx2_ASAP7_75t_L g1817 ( .A(n_1765), .Y(n_1817) );
NAND2xp5_ASAP7_75t_L g1858 ( .A(n_1769), .B(n_1859), .Y(n_1858) );
CKINVDCx14_ASAP7_75t_R g1876 ( .A(n_1770), .Y(n_1876) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_1772), .B(n_1773), .Y(n_1771) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
NAND5xp2_ASAP7_75t_L g1775 ( .A(n_1776), .B(n_1854), .C(n_1861), .D(n_1870), .E(n_1877), .Y(n_1775) );
AOI321xp33_ASAP7_75t_SL g1776 ( .A1(n_1777), .A2(n_1799), .A3(n_1800), .B1(n_1827), .B2(n_1830), .C(n_1840), .Y(n_1776) );
NAND3xp33_ASAP7_75t_SL g1777 ( .A(n_1778), .B(n_1784), .C(n_1790), .Y(n_1777) );
INVxp67_ASAP7_75t_L g1891 ( .A(n_1778), .Y(n_1891) );
NAND2xp5_ASAP7_75t_L g1778 ( .A(n_1779), .B(n_1780), .Y(n_1778) );
NAND2xp5_ASAP7_75t_L g1890 ( .A(n_1779), .B(n_1806), .Y(n_1890) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
A2O1A1Ixp33_ASAP7_75t_L g1840 ( .A1(n_1781), .A2(n_1789), .B(n_1841), .C(n_1843), .Y(n_1840) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
AOI21xp5_ASAP7_75t_L g1784 ( .A1(n_1785), .A2(n_1787), .B(n_1788), .Y(n_1784) );
OR2x2_ASAP7_75t_L g1807 ( .A(n_1786), .B(n_1808), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1833 ( .A(n_1786), .B(n_1823), .Y(n_1833) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1792), .B(n_1793), .Y(n_1791) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1792), .Y(n_1862) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
A2O1A1Ixp33_ASAP7_75t_L g1800 ( .A1(n_1801), .A2(n_1803), .B(n_1811), .C(n_1818), .Y(n_1800) );
CKINVDCx14_ASAP7_75t_R g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
AND2x2_ASAP7_75t_L g1844 ( .A(n_1812), .B(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1812), .Y(n_1860) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1815), .Y(n_1867) );
NAND2xp5_ASAP7_75t_L g1819 ( .A(n_1820), .B(n_1822), .Y(n_1819) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
AND2x2_ASAP7_75t_L g1825 ( .A(n_1821), .B(n_1826), .Y(n_1825) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
AOI311xp33_ASAP7_75t_L g1861 ( .A1(n_1824), .A2(n_1862), .A3(n_1863), .B(n_1864), .C(n_1868), .Y(n_1861) );
INVxp67_ASAP7_75t_SL g1863 ( .A(n_1827), .Y(n_1863) );
INVx2_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
CKINVDCx14_ASAP7_75t_R g1832 ( .A(n_1833), .Y(n_1832) );
AOI21xp5_ASAP7_75t_L g1834 ( .A1(n_1835), .A2(n_1836), .B(n_1838), .Y(n_1834) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1835), .Y(n_1853) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
NAND2xp5_ASAP7_75t_L g1874 ( .A(n_1839), .B(n_1875), .Y(n_1874) );
AOI211xp5_ASAP7_75t_L g1880 ( .A1(n_1839), .A2(n_1881), .B(n_1883), .C(n_1885), .Y(n_1880) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
AOI21xp5_ASAP7_75t_L g1843 ( .A1(n_1844), .A2(n_1846), .B(n_1848), .Y(n_1843) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
INVxp67_ASAP7_75t_SL g1868 ( .A(n_1869), .Y(n_1868) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
INVxp67_ASAP7_75t_L g1883 ( .A(n_1884), .Y(n_1883) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
INVxp67_ASAP7_75t_L g1889 ( .A(n_1890), .Y(n_1889) );
CKINVDCx20_ASAP7_75t_R g1893 ( .A(n_1894), .Y(n_1893) );
CKINVDCx20_ASAP7_75t_R g1894 ( .A(n_1895), .Y(n_1894) );
INVx2_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
XNOR2x1_ASAP7_75t_L g1897 ( .A(n_1898), .B(n_1948), .Y(n_1897) );
NOR2x1_ASAP7_75t_L g1898 ( .A(n_1899), .B(n_1910), .Y(n_1898) );
NAND2xp5_ASAP7_75t_L g1904 ( .A(n_1905), .B(n_1906), .Y(n_1904) );
NAND2xp5_ASAP7_75t_L g1910 ( .A(n_1911), .B(n_1931), .Y(n_1910) );
OAI31xp33_ASAP7_75t_L g1911 ( .A1(n_1912), .A2(n_1920), .A3(n_1928), .B(n_1930), .Y(n_1911) );
INVxp67_ASAP7_75t_SL g1921 ( .A(n_1922), .Y(n_1921) );
INVx2_ASAP7_75t_L g1938 ( .A(n_1939), .Y(n_1938) );
INVx1_ASAP7_75t_L g1941 ( .A(n_1942), .Y(n_1941) );
INVx3_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
HB1xp67_ASAP7_75t_L g1953 ( .A(n_1954), .Y(n_1953) );
BUFx3_ASAP7_75t_L g1954 ( .A(n_1955), .Y(n_1954) );
INVxp33_ASAP7_75t_SL g1956 ( .A(n_1957), .Y(n_1956) );
HB1xp67_ASAP7_75t_L g1958 ( .A(n_1959), .Y(n_1958) );
AND3x1_ASAP7_75t_L g1959 ( .A(n_1960), .B(n_1981), .C(n_1989), .Y(n_1959) );
NOR2xp33_ASAP7_75t_SL g1960 ( .A(n_1961), .B(n_1976), .Y(n_1960) );
HB1xp67_ASAP7_75t_L g1995 ( .A(n_1996), .Y(n_1995) );
INVx1_ASAP7_75t_L g1998 ( .A(n_1999), .Y(n_1998) );
endmodule