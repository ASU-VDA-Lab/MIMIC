module real_aes_5231_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_987;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_983;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_961;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_106;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_984;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_962;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_960;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_973;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_756;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_928;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_922;
wire n_633;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_982;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_0), .A2(n_126), .B1(n_127), .B2(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_1), .B(n_305), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_2), .Y(n_628) );
INVx1_ASAP7_75t_L g268 ( .A(n_3), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_SL g661 ( .A1(n_4), .A2(n_185), .B(n_662), .C(n_663), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_5), .A2(n_94), .B1(n_961), .B2(n_962), .Y(n_960) );
INVx1_ASAP7_75t_L g962 ( .A(n_5), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_6), .A2(n_83), .B1(n_156), .B2(n_177), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_7), .B(n_155), .Y(n_226) );
INVxp67_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
BUFx2_ASAP7_75t_L g969 ( .A(n_8), .Y(n_969) );
INVx1_ASAP7_75t_L g980 ( .A(n_8), .Y(n_980) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_9), .B(n_228), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_10), .A2(n_38), .B1(n_154), .B2(n_161), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_11), .A2(n_43), .B1(n_198), .B2(n_202), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_12), .A2(n_65), .B1(n_206), .B2(n_276), .Y(n_283) );
INVx1_ASAP7_75t_L g262 ( .A(n_13), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_14), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_15), .A2(n_73), .B1(n_177), .B2(n_200), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_16), .B(n_579), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_17), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_18), .B(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g266 ( .A(n_19), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_20), .A2(n_63), .B1(n_156), .B2(n_181), .Y(n_679) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_21), .A2(n_72), .B(n_145), .Y(n_144) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_21), .A2(n_72), .B(n_145), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_22), .A2(n_69), .B1(n_206), .B2(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g259 ( .A(n_23), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_24), .Y(n_641) );
BUFx3_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
BUFx8_ASAP7_75t_SL g989 ( .A(n_25), .Y(n_989) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_26), .A2(n_282), .B(n_668), .C(n_669), .Y(n_667) );
OAI22xp33_ASAP7_75t_SL g617 ( .A1(n_27), .A2(n_47), .B1(n_152), .B2(n_156), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_28), .A2(n_36), .B1(n_152), .B2(n_224), .Y(n_607) );
AO22x1_ASAP7_75t_L g221 ( .A1(n_29), .A2(n_79), .B1(n_183), .B2(n_222), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_30), .Y(n_173) );
AND2x2_ASAP7_75t_L g293 ( .A(n_31), .B(n_202), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_32), .B(n_183), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_L g688 ( .A1(n_33), .A2(n_185), .B(n_689), .C(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g123 ( .A(n_34), .Y(n_123) );
AOI22x1_ASAP7_75t_L g205 ( .A1(n_35), .A2(n_98), .B1(n_150), .B2(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_37), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g108 ( .A(n_39), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_40), .B(n_611), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_41), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_42), .B(n_240), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_44), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_45), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_46), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g145 ( .A(n_48), .Y(n_145) );
AND2x4_ASAP7_75t_L g147 ( .A(n_49), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g605 ( .A(n_49), .B(n_148), .Y(n_605) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_50), .Y(n_142) );
INVx2_ASAP7_75t_L g278 ( .A(n_51), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_52), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_53), .A2(n_185), .B(n_644), .C(n_645), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_54), .Y(n_696) );
INVx2_ASAP7_75t_L g712 ( .A(n_55), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_56), .Y(n_625) );
INVx1_ASAP7_75t_L g573 ( .A(n_57), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_57), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_58), .A2(n_75), .B1(n_150), .B2(n_154), .Y(n_149) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_59), .Y(n_231) );
AND2x2_ASAP7_75t_L g298 ( .A(n_60), .B(n_183), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_61), .B(n_235), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_62), .A2(n_81), .B1(n_199), .B2(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_64), .B(n_246), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_66), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_67), .B(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_68), .A2(n_960), .B1(n_963), .B2(n_964), .Y(n_959) );
BUFx4f_ASAP7_75t_SL g965 ( .A(n_68), .Y(n_965) );
NAND2xp33_ASAP7_75t_R g682 ( .A(n_70), .B(n_144), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_70), .A2(n_101), .B1(n_254), .B2(n_611), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_71), .B(n_192), .Y(n_301) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_74), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_76), .B(n_155), .Y(n_241) );
OR2x6_ASAP7_75t_L g120 ( .A(n_77), .B(n_121), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_78), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_80), .Y(n_708) );
INVx1_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
INVx1_ASAP7_75t_L g109 ( .A(n_84), .Y(n_109) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
BUFx5_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g201 ( .A(n_85), .Y(n_201) );
INVxp33_ASAP7_75t_SL g572 ( .A(n_86), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_86), .Y(n_574) );
INVx2_ASAP7_75t_L g674 ( .A(n_87), .Y(n_674) );
INVx2_ASAP7_75t_L g270 ( .A(n_88), .Y(n_270) );
INVx2_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_90), .Y(n_670) );
XOR2x2_ASAP7_75t_SL g958 ( .A(n_91), .B(n_959), .Y(n_958) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_92), .B(n_151), .Y(n_295) );
INVx2_ASAP7_75t_SL g148 ( .A(n_93), .Y(n_148) );
INVx1_ASAP7_75t_L g961 ( .A(n_94), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_95), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_96), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g694 ( .A(n_97), .Y(n_694) );
INVx2_ASAP7_75t_L g699 ( .A(n_99), .Y(n_699) );
OAI21xp33_ASAP7_75t_SL g639 ( .A1(n_100), .A2(n_156), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_101), .B(n_611), .Y(n_702) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_101), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_102), .B(n_190), .Y(n_189) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_113), .B1(n_581), .B2(n_588), .C(n_985), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_110), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_107), .B(n_587), .Y(n_586) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_108), .A2(n_988), .B(n_990), .Y(n_987) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx6p67_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_112), .Y(n_587) );
OAI21x1_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_124), .B(n_578), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
BUFx8_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx12f_ASAP7_75t_L g580 ( .A(n_116), .Y(n_580) );
INVx2_ASAP7_75t_SL g584 ( .A(n_116), .Y(n_584) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_116), .Y(n_992) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx1_ASAP7_75t_L g966 ( .A(n_119), .Y(n_966) );
INVx8_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x6_ASAP7_75t_L g979 ( .A(n_120), .B(n_980), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B1(n_130), .B2(n_577), .Y(n_124) );
INVx1_ASAP7_75t_SL g577 ( .A(n_125), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_126), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_126), .B(n_236), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_128), .Y(n_986) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
XNOR2x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_570), .Y(n_130) );
INVx2_ASAP7_75t_L g970 ( .A(n_131), .Y(n_970) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_463), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_375), .C(n_411), .Y(n_132) );
NAND3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_308), .C(n_353), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_212), .B1(n_284), .B2(n_287), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g566 ( .A(n_136), .Y(n_566) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_167), .Y(n_136) );
INVx2_ASAP7_75t_L g328 ( .A(n_137), .Y(n_328) );
INVx2_ASAP7_75t_L g455 ( .A(n_137), .Y(n_455) );
INVx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g307 ( .A(n_138), .B(n_168), .Y(n_307) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_157), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_139), .B(n_157), .Y(n_323) );
OR2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_149), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_141), .A2(n_154), .B1(n_171), .B2(n_175), .Y(n_170) );
INVx4_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_141), .A2(n_239), .B(n_241), .Y(n_238) );
OA22x2_ASAP7_75t_L g606 ( .A1(n_141), .A2(n_159), .B1(n_607), .B2(n_608), .Y(n_606) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g159 ( .A(n_142), .Y(n_159) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_142), .B(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_142), .B(n_262), .Y(n_261) );
INVx4_ASAP7_75t_L g265 ( .A(n_142), .Y(n_265) );
INVx3_ASAP7_75t_L g282 ( .A(n_142), .Y(n_282) );
INVxp67_ASAP7_75t_L g296 ( .A(n_142), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_142), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_142), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_143), .B(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_L g255 ( .A(n_144), .Y(n_255) );
BUFx3_ASAP7_75t_L g604 ( .A(n_144), .Y(n_604) );
INVx1_ASAP7_75t_L g637 ( .A(n_144), .Y(n_637) );
INVx1_ASAP7_75t_L g700 ( .A(n_144), .Y(n_700) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
INVx1_ASAP7_75t_L g218 ( .A(n_147), .Y(n_218) );
INVx3_ASAP7_75t_L g249 ( .A(n_147), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_147), .B(n_193), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_147), .A2(n_185), .B1(n_282), .B2(n_624), .C(n_627), .Y(n_623) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx1_ASAP7_75t_L g240 ( .A(n_152), .Y(n_240) );
INVx2_ASAP7_75t_SL g609 ( .A(n_152), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_152), .A2(n_156), .B1(n_625), .B2(n_626), .Y(n_624) );
INVx2_ASAP7_75t_L g664 ( .A(n_152), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_152), .A2(n_156), .B1(n_707), .B2(n_708), .Y(n_706) );
INVx6_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g163 ( .A(n_153), .Y(n_163) );
INVx2_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
INVx2_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
INVx2_ASAP7_75t_L g207 ( .A(n_156), .Y(n_207) );
INVx2_ASAP7_75t_L g246 ( .A(n_156), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_156), .A2(n_181), .B1(n_628), .B2(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_156), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_156), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_156), .B(n_696), .Y(n_695) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_164), .Y(n_157) );
INVx1_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g276 ( .A(n_162), .Y(n_276) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g228 ( .A(n_163), .Y(n_228) );
INVx2_ASAP7_75t_L g244 ( .A(n_163), .Y(n_244) );
INVx1_ASAP7_75t_L g644 ( .A(n_163), .Y(n_644) );
INVx1_ASAP7_75t_L g689 ( .A(n_163), .Y(n_689) );
INVx1_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OR2x2_ASAP7_75t_L g403 ( .A(n_167), .B(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_167), .Y(n_551) );
NAND2x1_ASAP7_75t_L g167 ( .A(n_168), .B(n_194), .Y(n_167) );
AND2x2_ASAP7_75t_L g349 ( .A(n_168), .B(n_323), .Y(n_349) );
AND2x2_ASAP7_75t_L g495 ( .A(n_168), .B(n_331), .Y(n_495) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_187), .B(n_189), .Y(n_168) );
OA21x2_ASAP7_75t_L g325 ( .A1(n_169), .A2(n_187), .B(n_189), .Y(n_325) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_178), .B(n_186), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI22x1_ASAP7_75t_L g196 ( .A1(n_174), .A2(n_197), .B1(n_204), .B2(n_205), .Y(n_196) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_184), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_180), .B(n_261), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_180), .A2(n_183), .B1(n_264), .B2(n_267), .Y(n_263) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g668 ( .A(n_181), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_181), .A2(n_224), .B1(n_711), .B2(n_712), .Y(n_710) );
INVxp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g220 ( .A(n_185), .Y(n_220) );
INVx2_ASAP7_75t_SL g229 ( .A(n_185), .Y(n_229) );
INVx1_ASAP7_75t_L g247 ( .A(n_185), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_185), .A2(n_265), .B1(n_679), .B2(n_680), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_185), .A2(n_265), .B1(n_706), .B2(n_710), .Y(n_736) );
AO31x2_ASAP7_75t_L g195 ( .A1(n_186), .A2(n_196), .A3(n_208), .B(n_209), .Y(n_195) );
AO31x2_ASAP7_75t_L g289 ( .A1(n_186), .A2(n_196), .A3(n_208), .B(n_209), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_186), .B(n_603), .Y(n_735) );
INVx3_ASAP7_75t_L g211 ( .A(n_187), .Y(n_211) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx4_ASAP7_75t_L g193 ( .A(n_188), .Y(n_193) );
INVx2_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
OR2x2_ASAP7_75t_L g217 ( .A(n_190), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g277 ( .A(n_191), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g305 ( .A(n_193), .Y(n_305) );
INVx2_ASAP7_75t_L g611 ( .A(n_193), .Y(n_611) );
NOR2xp33_ASAP7_75t_SL g673 ( .A(n_193), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g321 ( .A(n_194), .Y(n_321) );
INVx1_ASAP7_75t_L g340 ( .A(n_194), .Y(n_340) );
AND2x2_ASAP7_75t_L g348 ( .A(n_194), .B(n_291), .Y(n_348) );
AND2x2_ASAP7_75t_L g484 ( .A(n_194), .B(n_364), .Y(n_484) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g356 ( .A(n_195), .B(n_324), .Y(n_356) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g662 ( .A(n_199), .Y(n_662) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g224 ( .A(n_201), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_202), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp67_ASAP7_75t_SL g209 ( .A(n_210), .B(n_211), .Y(n_209) );
OR2x2_ASAP7_75t_L g230 ( .A(n_211), .B(n_231), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_211), .A2(n_718), .B(n_719), .Y(n_717) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g560 ( .A(n_213), .Y(n_560) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_250), .Y(n_213) );
OR2x2_ASAP7_75t_L g414 ( .A(n_214), .B(n_334), .Y(n_414) );
OR2x2_ASAP7_75t_SL g524 ( .A(n_214), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g284 ( .A(n_215), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g468 ( .A(n_215), .B(n_427), .Y(n_468) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_232), .Y(n_215) );
INVx2_ASAP7_75t_SL g346 ( .A(n_216), .Y(n_346) );
AND2x2_ASAP7_75t_L g352 ( .A(n_216), .B(n_233), .Y(n_352) );
OAI21x1_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_219), .B(n_230), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_217), .A2(n_219), .B(n_230), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_218), .B(n_254), .Y(n_253) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_218), .B(n_235), .Y(n_681) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_225), .Y(n_219) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_224), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_224), .B(n_670), .Y(n_669) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_229), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_228), .A2(n_265), .B1(n_693), .B2(n_695), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_229), .B(n_301), .Y(n_302) );
INVx1_ASAP7_75t_L g390 ( .A(n_232), .Y(n_390) );
AND2x2_ASAP7_75t_L g474 ( .A(n_232), .B(n_271), .Y(n_474) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g312 ( .A(n_233), .Y(n_312) );
AND2x2_ASAP7_75t_L g345 ( .A(n_233), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
NOR2x1_ASAP7_75t_L g248 ( .A(n_235), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_236), .B(n_270), .Y(n_269) );
BUFx3_ASAP7_75t_L g697 ( .A(n_236), .Y(n_697) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_242), .B(n_248), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_245), .B(n_247), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_247), .A2(n_642), .B1(n_672), .B2(n_705), .C(n_709), .Y(n_704) );
INVx2_ASAP7_75t_L g274 ( .A(n_249), .Y(n_274) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g351 ( .A(n_251), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_251), .B(n_452), .Y(n_451) );
NAND2x1_ASAP7_75t_SL g489 ( .A(n_251), .B(n_345), .Y(n_489) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_251), .Y(n_500) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_271), .Y(n_251) );
INVx1_ASAP7_75t_L g286 ( .A(n_252), .Y(n_286) );
INVxp67_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
OR2x2_ASAP7_75t_L g336 ( .A(n_252), .B(n_315), .Y(n_336) );
INVx1_ASAP7_75t_L g398 ( .A(n_252), .Y(n_398) );
INVx1_ASAP7_75t_L g410 ( .A(n_252), .Y(n_410) );
AND2x2_ASAP7_75t_L g445 ( .A(n_252), .B(n_346), .Y(n_445) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .B(n_269), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND3xp33_ASAP7_75t_SL g273 ( .A(n_255), .B(n_265), .C(n_274), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_255), .B(n_274), .C(n_281), .Y(n_280) );
NAND3xp33_ASAP7_75t_SL g256 ( .A(n_257), .B(n_260), .C(n_263), .Y(n_256) );
NOR2xp33_ASAP7_75t_SL g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_265), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g642 ( .A(n_265), .Y(n_642) );
AND2x2_ASAP7_75t_L g285 ( .A(n_271), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
INVx1_ASAP7_75t_L g334 ( .A(n_271), .Y(n_334) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_271), .Y(n_379) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_271), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g428 ( .A(n_271), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_271), .Y(n_431) );
OR2x6_ASAP7_75t_L g271 ( .A(n_272), .B(n_279), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B(n_277), .Y(n_272) );
AOI21xp33_ASAP7_75t_SL g303 ( .A1(n_274), .A2(n_304), .B(n_306), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_282), .A2(n_619), .B(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g427 ( .A(n_286), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_307), .Y(n_287) );
BUFx3_ASAP7_75t_L g358 ( .A(n_288), .Y(n_358) );
INVx3_ASAP7_75t_L g456 ( .A(n_288), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_288), .B(n_362), .Y(n_556) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OR2x2_ASAP7_75t_L g330 ( .A(n_289), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g374 ( .A(n_289), .B(n_331), .Y(n_374) );
INVx1_ASAP7_75t_L g460 ( .A(n_289), .Y(n_460) );
INVx1_ASAP7_75t_L g450 ( .A(n_290), .Y(n_450) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_L g361 ( .A(n_291), .Y(n_361) );
INVx1_ASAP7_75t_L g442 ( .A(n_291), .Y(n_442) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_297), .B(n_303), .Y(n_291) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_292), .A2(n_297), .B(n_303), .Y(n_331) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21x1_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_299), .B(n_302), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g306 ( .A(n_301), .Y(n_306) );
INVx2_ASAP7_75t_L g622 ( .A(n_304), .Y(n_622) );
OR2x2_ASAP7_75t_L g737 ( .A(n_304), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_SL g671 ( .A(n_305), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g367 ( .A(n_307), .Y(n_367) );
AND2x2_ASAP7_75t_L g480 ( .A(n_307), .B(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_307), .Y(n_513) );
NOR2xp67_ASAP7_75t_SL g518 ( .A(n_307), .B(n_456), .Y(n_518) );
INVx1_ASAP7_75t_L g546 ( .A(n_307), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_317), .B1(n_326), .B2(n_332), .C(n_337), .Y(n_308) );
INVx2_ASAP7_75t_L g488 ( .A(n_309), .Y(n_488) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_311), .Y(n_400) );
AND2x2_ASAP7_75t_L g333 ( .A(n_312), .B(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
INVx2_ASAP7_75t_L g452 ( .A(n_312), .Y(n_452) );
OR2x2_ASAP7_75t_L g469 ( .A(n_312), .B(n_336), .Y(n_469) );
AND2x2_ASAP7_75t_L g552 ( .A(n_313), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_316), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_316), .B(n_445), .Y(n_569) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g386 ( .A(n_320), .B(n_341), .Y(n_386) );
INVx1_ASAP7_75t_L g492 ( .A(n_320), .Y(n_492) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g521 ( .A(n_321), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_322), .Y(n_522) );
INVx2_ASAP7_75t_L g564 ( .A(n_322), .Y(n_564) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g364 ( .A(n_323), .Y(n_364) );
INVx1_ASAP7_75t_L g385 ( .A(n_323), .Y(n_385) );
INVx1_ASAP7_75t_L g419 ( .A(n_323), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_323), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_324), .B(n_364), .Y(n_508) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g342 ( .A(n_325), .Y(n_342) );
OAI31xp33_ASAP7_75t_L g548 ( .A1(n_326), .A2(n_549), .A3(n_550), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND3x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_361), .C(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g373 ( .A(n_328), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g381 ( .A(n_330), .B(n_362), .Y(n_381) );
INVx2_ASAP7_75t_L g481 ( .A(n_330), .Y(n_481) );
AND2x4_ASAP7_75t_L g341 ( .A(n_331), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NAND2x2_ASAP7_75t_L g443 ( .A(n_333), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g344 ( .A(n_334), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g370 ( .A(n_335), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .B1(n_347), .B2(n_350), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
NAND2xp67_ASAP7_75t_L g416 ( .A(n_339), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_339), .Y(n_422) );
AND2x4_ASAP7_75t_SL g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g437 ( .A(n_340), .Y(n_437) );
AND2x2_ASAP7_75t_L g543 ( .A(n_340), .B(n_349), .Y(n_543) );
AND2x2_ASAP7_75t_L g363 ( .A(n_341), .B(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g397 ( .A(n_341), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_341), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_342), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_344), .A2(n_363), .B1(n_466), .B2(n_470), .C(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
INVx1_ASAP7_75t_L g531 ( .A(n_346), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g432 ( .A(n_349), .B(n_361), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_349), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_351), .Y(n_365) );
INVx2_ASAP7_75t_L g406 ( .A(n_352), .Y(n_406) );
AND2x2_ASAP7_75t_L g502 ( .A(n_352), .B(n_503), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_363), .B(n_365), .C(n_366), .Y(n_353) );
NAND3xp33_ASAP7_75t_SL g354 ( .A(n_355), .B(n_357), .C(n_359), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_356), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_361), .Y(n_515) );
OR2x2_ASAP7_75t_L g511 ( .A(n_362), .B(n_441), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_369), .B2(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g529 ( .A(n_371), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g558 ( .A(n_374), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_381), .B1(n_382), .B2(n_387), .C(n_392), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AND2x2_ASAP7_75t_L g430 ( .A(n_380), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g475 ( .A(n_380), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g526 ( .A1(n_381), .A2(n_527), .B(n_528), .Y(n_526) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AND2x2_ASAP7_75t_L g393 ( .A(n_384), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_384), .B(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_384), .A2(n_455), .B1(n_467), .B2(n_469), .Y(n_466) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g498 ( .A(n_388), .Y(n_498) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp67_ASAP7_75t_SL g434 ( .A(n_389), .B(n_398), .Y(n_434) );
OR2x2_ASAP7_75t_L g461 ( .A(n_389), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_390), .Y(n_394) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_391), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_398), .C(n_399), .Y(n_392) );
INVx1_ASAP7_75t_L g540 ( .A(n_394), .Y(n_540) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_396), .B(n_472), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_396), .A2(n_443), .B1(n_501), .B2(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g479 ( .A(n_398), .Y(n_479) );
AND2x2_ASAP7_75t_L g530 ( .A(n_398), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g553 ( .A(n_398), .B(n_452), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_407), .Y(n_399) );
INVx1_ASAP7_75t_L g503 ( .A(n_400), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_402), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_406), .A2(n_477), .B1(n_482), .B2(n_485), .C(n_487), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_407), .B(n_452), .Y(n_542) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g486 ( .A(n_408), .B(n_452), .Y(n_486) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_420), .C(n_433), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_417), .B(n_447), .Y(n_534) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21x1_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_429), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_430), .A2(n_555), .B1(n_557), .B2(n_560), .C(n_561), .Y(n_554) );
INVx2_ASAP7_75t_L g525 ( .A(n_431), .Y(n_525) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_438), .C(n_453), .Y(n_433) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_443), .B1(n_446), .B2(n_451), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g547 ( .A(n_445), .B(n_474), .Y(n_547) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B(n_457), .C(n_461), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g527 ( .A(n_455), .B(n_494), .Y(n_527) );
AND2x2_ASAP7_75t_L g549 ( .A(n_455), .B(n_495), .Y(n_549) );
INVx1_ASAP7_75t_L g470 ( .A(n_457), .Y(n_470) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g463 ( .A(n_464), .B(n_516), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .C(n_496), .Y(n_464) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_481), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_488), .B(n_513), .C(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_510), .C(n_512), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_501), .C(n_504), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND4xp25_ASAP7_75t_SL g516 ( .A(n_517), .B(n_532), .C(n_548), .D(n_554), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_519), .B(n_523), .C(n_526), .Y(n_517) );
INVxp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
OR2x2_ASAP7_75t_L g545 ( .A(n_521), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g538 ( .A(n_525), .Y(n_538) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B1(n_541), .B2(n_543), .C1(n_544), .C2(n_547), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g559 ( .A(n_543), .Y(n_559) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B(n_567), .Y(n_561) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_576), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_981), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_967), .B(n_971), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_957), .Y(n_590) );
INVx1_ASAP7_75t_L g972 ( .A(n_591), .Y(n_972) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND4xp75_ASAP7_75t_L g593 ( .A(n_594), .B(n_802), .C(n_897), .D(n_922), .Y(n_593) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_756), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_713), .Y(n_595) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_631), .B(n_656), .Y(n_596) );
INVx1_ASAP7_75t_L g906 ( .A(n_597), .Y(n_906) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_612), .Y(n_598) );
AND2x2_ASAP7_75t_L g769 ( .A(n_599), .B(n_770), .Y(n_769) );
INVx3_ASAP7_75t_L g813 ( .A(n_599), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_599), .B(n_653), .Y(n_863) );
AND2x4_ASAP7_75t_L g889 ( .A(n_599), .B(n_752), .Y(n_889) );
INVx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g761 ( .A(n_600), .B(n_648), .Y(n_761) );
INVx1_ASAP7_75t_L g773 ( .A(n_600), .Y(n_773) );
AND2x2_ASAP7_75t_L g800 ( .A(n_600), .B(n_621), .Y(n_800) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g655 ( .A(n_601), .Y(n_655) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_606), .B(n_610), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g636 ( .A(n_605), .B(n_637), .Y(n_636) );
INVx4_ASAP7_75t_L g672 ( .A(n_605), .Y(n_672) );
INVx1_ASAP7_75t_L g718 ( .A(n_606), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_610), .Y(n_719) );
AND2x2_ASAP7_75t_L g883 ( .A(n_612), .B(n_760), .Y(n_883) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_621), .Y(n_612) );
INVx2_ASAP7_75t_L g648 ( .A(n_613), .Y(n_648) );
INVx3_ASAP7_75t_L g654 ( .A(n_613), .Y(n_654) );
AND2x2_ASAP7_75t_L g770 ( .A(n_613), .B(n_634), .Y(n_770) );
INVx1_ASAP7_75t_L g792 ( .A(n_613), .Y(n_792) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_613), .Y(n_796) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
OR2x2_ASAP7_75t_L g749 ( .A(n_621), .B(n_717), .Y(n_749) );
AND2x4_ASAP7_75t_L g752 ( .A(n_621), .B(n_654), .Y(n_752) );
AND2x2_ASAP7_75t_L g772 ( .A(n_621), .B(n_773), .Y(n_772) );
OA21x2_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B(n_630), .Y(n_621) );
OA21x2_ASAP7_75t_L g651 ( .A1(n_622), .A2(n_623), .B(n_630), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_649), .B(n_652), .Y(n_631) );
AND2x2_ASAP7_75t_L g896 ( .A(n_632), .B(n_748), .Y(n_896) );
AND2x2_ASAP7_75t_L g941 ( .A(n_632), .B(n_716), .Y(n_941) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g812 ( .A(n_633), .B(n_813), .Y(n_812) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_633), .Y(n_860) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_648), .Y(n_633) );
AND2x2_ASAP7_75t_L g653 ( .A(n_634), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g729 ( .A(n_634), .B(n_650), .Y(n_729) );
INVx2_ASAP7_75t_L g760 ( .A(n_634), .Y(n_760) );
INVx1_ASAP7_75t_L g780 ( .A(n_634), .Y(n_780) );
BUFx2_ASAP7_75t_L g810 ( .A(n_634), .Y(n_810) );
INVx2_ASAP7_75t_L g845 ( .A(n_634), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_634), .B(n_651), .Y(n_912) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI21x1_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_647), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B(n_643), .Y(n_638) );
AND2x4_ASAP7_75t_L g819 ( .A(n_648), .B(n_720), .Y(n_819) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_650), .B(n_780), .Y(n_797) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g720 ( .A(n_651), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx2_ASAP7_75t_L g945 ( .A(n_653), .Y(n_945) );
INVx1_ASAP7_75t_L g715 ( .A(n_654), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_654), .B(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g793 ( .A(n_655), .Y(n_793) );
OR2x2_ASAP7_75t_L g843 ( .A(n_655), .B(n_844), .Y(n_843) );
AND2x2_ASAP7_75t_L g855 ( .A(n_655), .B(n_760), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_655), .B(n_796), .Y(n_881) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_683), .Y(n_656) );
AND2x2_ASAP7_75t_L g884 ( .A(n_657), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_675), .Y(n_657) );
AND2x2_ASAP7_75t_L g732 ( .A(n_658), .B(n_686), .Y(n_732) );
INVx1_ASAP7_75t_L g892 ( .A(n_658), .Y(n_892) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_659), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_659), .B(n_686), .Y(n_755) );
AND2x4_ASAP7_75t_L g764 ( .A(n_659), .B(n_734), .Y(n_764) );
INVx1_ASAP7_75t_L g809 ( .A(n_659), .Y(n_809) );
INVx1_ASAP7_75t_L g832 ( .A(n_659), .Y(n_832) );
OR2x2_ASAP7_75t_L g853 ( .A(n_659), .B(n_701), .Y(n_853) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_659), .Y(n_868) );
AND2x2_ASAP7_75t_L g895 ( .A(n_659), .B(n_701), .Y(n_895) );
AO31x2_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_666), .A3(n_671), .B(n_673), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_672), .B(n_688), .C(n_692), .Y(n_687) );
AND2x4_ASAP7_75t_L g724 ( .A(n_675), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g838 ( .A(n_675), .Y(n_838) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g733 ( .A(n_676), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g766 ( .A(n_676), .Y(n_766) );
AND2x2_ASAP7_75t_L g893 ( .A(n_676), .B(n_685), .Y(n_893) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_676), .Y(n_929) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_682), .Y(n_676) );
AND2x2_ASAP7_75t_L g743 ( .A(n_677), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_681), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_701), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_684), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g758 ( .A(n_685), .B(n_742), .Y(n_758) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_685), .Y(n_827) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g725 ( .A(n_686), .Y(n_725) );
AND2x2_ASAP7_75t_L g765 ( .A(n_686), .B(n_766), .Y(n_765) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_686), .Y(n_823) );
BUFx2_ASAP7_75t_R g872 ( .A(n_686), .Y(n_872) );
AO21x2_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_697), .B(n_698), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_697), .B(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_701), .Y(n_723) );
AND2x2_ASAP7_75t_L g808 ( .A(n_701), .B(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_701), .B(n_725), .Y(n_886) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
AND2x2_ASAP7_75t_L g742 ( .A(n_703), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_721), .B(n_726), .C(n_750), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
AND2x2_ASAP7_75t_L g747 ( .A(n_715), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g781 ( .A(n_716), .Y(n_781) );
INVx2_ASAP7_75t_SL g943 ( .A(n_716), .Y(n_943) );
AND2x4_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g900 ( .A(n_723), .Y(n_900) );
AND2x2_ASAP7_75t_L g801 ( .A(n_724), .B(n_764), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_724), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g940 ( .A(n_724), .Y(n_940) );
OR2x2_ASAP7_75t_L g877 ( .A(n_725), .B(n_845), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B1(n_739), .B2(n_746), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g932 ( .A(n_729), .B(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g762 ( .A1(n_731), .A2(n_752), .B1(n_763), .B2(n_767), .C1(n_774), .C2(n_777), .Y(n_762) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g776 ( .A(n_732), .Y(n_776) );
AND2x4_ASAP7_75t_L g815 ( .A(n_733), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g935 ( .A(n_733), .B(n_809), .Y(n_935) );
INVx1_ASAP7_75t_L g842 ( .A(n_734), .Y(n_842) );
OAI21x1_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B(n_737), .Y(n_734) );
HB1xp67_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g931 ( .A(n_740), .Y(n_931) );
OR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .Y(n_740) );
OR2x2_ASAP7_75t_L g951 ( .A(n_741), .B(n_809), .Y(n_951) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g754 ( .A(n_742), .Y(n_754) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g918 ( .A(n_748), .B(n_830), .Y(n_918) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g785 ( .A(n_749), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .Y(n_750) );
OR2x2_ASAP7_75t_L g786 ( .A(n_751), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g854 ( .A(n_752), .B(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_752), .B(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g904 ( .A(n_752), .B(n_813), .Y(n_904) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
OR2x2_ASAP7_75t_L g775 ( .A(n_754), .B(n_776), .Y(n_775) );
OR2x2_ASAP7_75t_L g848 ( .A(n_754), .B(n_827), .Y(n_848) );
INVx1_ASAP7_75t_L g816 ( .A(n_755), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_762), .C(n_782), .Y(n_756) );
NAND2xp33_ASAP7_75t_R g757 ( .A(n_758), .B(n_759), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g917 ( .A1(n_759), .A2(n_918), .B(n_919), .Y(n_917) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g789 ( .A(n_760), .Y(n_789) );
INVx1_ASAP7_75t_L g830 ( .A(n_760), .Y(n_830) );
OAI21xp5_ASAP7_75t_L g934 ( .A1(n_763), .A2(n_935), .B(n_936), .Y(n_934) );
AND2x4_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AND2x2_ASAP7_75t_L g821 ( .A(n_764), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_SL g839 ( .A(n_764), .Y(n_839) );
NAND2xp33_ASAP7_75t_L g807 ( .A(n_765), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_SL g865 ( .A(n_765), .Y(n_865) );
AND2x2_ASAP7_75t_L g894 ( .A(n_765), .B(n_895), .Y(n_894) );
NAND2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g874 ( .A(n_769), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_770), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g902 ( .A(n_770), .B(n_813), .Y(n_902) );
INVx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g849 ( .A(n_772), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI21xp5_ASAP7_75t_SL g887 ( .A1(n_775), .A2(n_860), .B(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND3xp33_ASAP7_75t_SL g879 ( .A(n_778), .B(n_880), .C(n_882), .Y(n_879) );
OR2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI31xp33_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_790), .A3(n_798), .B(n_801), .Y(n_782) );
NAND2xp33_ASAP7_75t_SL g783 ( .A(n_784), .B(n_786), .Y(n_783) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_785), .B(n_860), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g905 ( .A1(n_786), .A2(n_831), .B1(n_839), .B2(n_906), .Y(n_905) );
OR2x2_ASAP7_75t_L g937 ( .A(n_787), .B(n_881), .Y(n_937) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
NOR2xp67_ASAP7_75t_L g911 ( .A(n_792), .B(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g933 ( .A(n_792), .Y(n_933) );
AND2x4_ASAP7_75t_L g818 ( .A(n_793), .B(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
INVxp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NOR2x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_856), .Y(n_802) );
NAND4xp75_ASAP7_75t_L g803 ( .A(n_804), .B(n_824), .C(n_833), .D(n_846), .Y(n_803) );
NOR2x1_ASAP7_75t_SL g804 ( .A(n_805), .B(n_811), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g927 ( .A(n_808), .B(n_928), .Y(n_927) );
NAND2x1p5_ASAP7_75t_L g948 ( .A(n_810), .B(n_819), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_814), .B1(n_817), .B2(n_820), .Y(n_811) );
AND2x2_ASAP7_75t_L g914 ( .A(n_813), .B(n_819), .Y(n_914) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g828 ( .A(n_818), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OR2x2_ASAP7_75t_L g852 ( .A(n_822), .B(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .C(n_831), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_829), .B(n_889), .Y(n_956) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_830), .B(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g921 ( .A(n_832), .Y(n_921) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_839), .B(n_840), .C(n_843), .Y(n_834) );
AOI221x1_ASAP7_75t_L g897 ( .A1(n_835), .A2(n_898), .B1(n_905), .B2(n_907), .C(n_908), .Y(n_897) );
BUFx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_836), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_839), .A2(n_870), .B1(n_874), .B2(n_875), .Y(n_869) );
INVx1_ASAP7_75t_L g949 ( .A(n_840), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_841), .B(n_865), .Y(n_916) );
AOI33xp33_ASAP7_75t_L g939 ( .A1(n_841), .A2(n_935), .A3(n_940), .B1(n_941), .B2(n_942), .B3(n_944), .Y(n_939) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx2_ASAP7_75t_L g850 ( .A(n_845), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_849), .B1(n_851), .B2(n_854), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g873 ( .A(n_853), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_878), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_861), .B(n_864), .C(n_869), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVxp67_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
BUFx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
OR2x2_ASAP7_75t_L g954 ( .A(n_865), .B(n_891), .Y(n_954) );
INVxp67_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_873), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_884), .B(n_887), .Y(n_878) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B1(n_894), .B2(n_896), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_889), .B(n_927), .Y(n_926) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
BUFx2_ASAP7_75t_L g907 ( .A(n_893), .Y(n_907) );
OAI21xp33_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_901), .B(n_903), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVxp33_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_913), .B(n_915), .C(n_917), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
BUFx2_ASAP7_75t_SL g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_914), .A2(n_947), .B1(n_949), .B2(n_950), .Y(n_946) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NOR2xp67_ASAP7_75t_L g922 ( .A(n_923), .B(n_938), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_934), .Y(n_923) );
INVxp67_ASAP7_75t_SL g924 ( .A(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_930), .Y(n_925) );
INVx2_ASAP7_75t_SL g928 ( .A(n_929), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_946), .C(n_952), .Y(n_938) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx2_ASAP7_75t_SL g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_955), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_957), .B(n_976), .Y(n_982) );
NAND2xp5_ASAP7_75t_SL g957 ( .A(n_958), .B(n_966), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_958), .Y(n_974) );
INVx1_ASAP7_75t_L g963 ( .A(n_960), .Y(n_963) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_965), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_966), .B(n_974), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_967), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_981) );
INVx1_ASAP7_75t_L g984 ( .A(n_967), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_968), .B(n_970), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_969), .Y(n_968) );
BUFx8_ASAP7_75t_L g976 ( .A(n_969), .Y(n_976) );
OAI31xp33_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .A3(n_975), .B(n_977), .Y(n_971) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_973), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_987), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx5_ASAP7_75t_SL g991 ( .A(n_992), .Y(n_991) );
endmodule