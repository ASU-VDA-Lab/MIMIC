module fake_aes_7453_n_871 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_871);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_871;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_58), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_75), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_95), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_52), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
BUFx5_ASAP7_75t_L g116 ( .A(n_94), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_87), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_40), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_53), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_7), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_107), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_7), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_42), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_91), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_101), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_10), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_97), .Y(n_127) );
BUFx10_ASAP7_75t_L g128 ( .A(n_11), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_30), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_83), .Y(n_130) );
BUFx10_ASAP7_75t_L g131 ( .A(n_33), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_60), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_23), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_4), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_102), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_106), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_16), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_38), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_74), .Y(n_139) );
INVx2_ASAP7_75t_SL g140 ( .A(n_84), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_86), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_68), .Y(n_142) );
BUFx10_ASAP7_75t_L g143 ( .A(n_45), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_41), .Y(n_145) );
BUFx10_ASAP7_75t_L g146 ( .A(n_17), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_108), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_66), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_31), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_70), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_33), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_48), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
INVx5_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_140), .B(n_0), .Y(n_155) );
BUFx12f_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_123), .B(n_0), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_115), .B(n_1), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_111), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_141), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_137), .B(n_1), .Y(n_164) );
NOR2xp33_ASAP7_75t_SL g165 ( .A(n_138), .B(n_37), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_128), .B(n_2), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_149), .B(n_2), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_114), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_109), .B(n_3), .Y(n_170) );
BUFx12f_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx5_ASAP7_75t_L g172 ( .A(n_109), .Y(n_172) );
BUFx8_ASAP7_75t_SL g173 ( .A(n_151), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_117), .B(n_3), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_121), .B(n_4), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_161), .A2(n_151), .B1(n_111), .B2(n_119), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_157), .A2(n_119), .B1(n_135), .B2(n_136), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_169), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_159), .A2(n_136), .B1(n_135), .B2(n_133), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_161), .A2(n_129), .B1(n_122), .B2(n_134), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_156), .B(n_124), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_156), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_159), .A2(n_126), .B1(n_144), .B2(n_148), .Y(n_187) );
BUFx10_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_157), .A2(n_131), .B1(n_128), .B2(n_146), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_170), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_157), .A2(n_131), .B1(n_128), .B2(n_146), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_170), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_169), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_157), .A2(n_131), .B1(n_146), .B2(n_145), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
OAI22xp33_ASAP7_75t_SL g197 ( .A1(n_161), .A2(n_152), .B1(n_150), .B2(n_147), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_156), .A2(n_127), .B1(n_142), .B2(n_139), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_166), .B(n_143), .Y(n_200) );
XNOR2xp5_ASAP7_75t_L g201 ( .A(n_166), .B(n_5), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
OR2x6_ASAP7_75t_L g203 ( .A(n_171), .B(n_5), .Y(n_203) );
OR2x6_ASAP7_75t_L g204 ( .A(n_171), .B(n_6), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_166), .B(n_116), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_171), .B(n_116), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_163), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_171), .B(n_116), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_174), .A2(n_132), .B1(n_130), .B2(n_125), .Y(n_210) );
NAND2xp33_ASAP7_75t_SL g211 ( .A(n_160), .B(n_112), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_173), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g214 ( .A1(n_160), .A2(n_118), .B1(n_113), .B2(n_10), .Y(n_214) );
OAI22xp33_ASAP7_75t_SL g215 ( .A1(n_164), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_174), .A2(n_116), .B1(n_13), .B2(n_14), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_168), .B(n_116), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_168), .B(n_116), .Y(n_218) );
BUFx6f_ASAP7_75t_SL g219 ( .A(n_168), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_175), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_12), .B1(n_16), .B2(n_17), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g222 ( .A1(n_167), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_188), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_188), .Y(n_224) );
XNOR2xp5_ASAP7_75t_L g225 ( .A(n_179), .B(n_173), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_207), .Y(n_227) );
XOR2xp5_ASAP7_75t_L g228 ( .A(n_181), .B(n_167), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_176), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_190), .B(n_175), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_192), .B(n_172), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
XNOR2xp5_ASAP7_75t_L g233 ( .A(n_178), .B(n_18), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_177), .B(n_172), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_217), .Y(n_236) );
XNOR2x2_ASAP7_75t_L g237 ( .A(n_208), .B(n_19), .Y(n_237) );
INVxp67_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_184), .B(n_200), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_218), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_196), .B(n_165), .Y(n_241) );
INVx4_ASAP7_75t_SL g242 ( .A(n_219), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_205), .Y(n_243) );
XOR2xp5_ASAP7_75t_L g244 ( .A(n_201), .B(n_20), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_198), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_219), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_219), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_203), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_198), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_186), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_212), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_185), .A2(n_172), .B(n_154), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_203), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_186), .B(n_172), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_183), .B(n_206), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_206), .A2(n_172), .B(n_165), .Y(n_260) );
XOR2xp5_ASAP7_75t_L g261 ( .A(n_201), .B(n_182), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_183), .B(n_172), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_185), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_204), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
NAND2xp33_ASAP7_75t_R g267 ( .A(n_204), .B(n_21), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_209), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_204), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
INVxp33_ASAP7_75t_L g271 ( .A(n_187), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_183), .B(n_172), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_216), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_193), .Y(n_274) );
INVx4_ASAP7_75t_SL g275 ( .A(n_183), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
XOR2xp5_ASAP7_75t_L g277 ( .A(n_189), .B(n_21), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_210), .B(n_165), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_191), .B(n_172), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_208), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_208), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_194), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_211), .B(n_172), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_223), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_242), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_239), .B(n_195), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_239), .B(n_199), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_243), .B(n_214), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_275), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_275), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_243), .B(n_197), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_245), .B(n_211), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_229), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_245), .B(n_215), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_223), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_249), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_275), .B(n_172), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_250), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_22), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_240), .B(n_221), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_249), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_238), .B(n_22), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_235), .B(n_23), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_240), .A2(n_222), .B(n_213), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_232), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_232), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_227), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_264), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_230), .B(n_24), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_230), .B(n_24), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_227), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_273), .B(n_213), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_252), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_264), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_250), .B(n_25), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_254), .Y(n_320) );
INVx8_ASAP7_75t_L g321 ( .A(n_262), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_281), .A2(n_202), .B1(n_194), .B2(n_162), .Y(n_322) );
AND2x2_ASAP7_75t_SL g323 ( .A(n_281), .B(n_162), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_252), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_242), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_234), .B(n_202), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_242), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_234), .B(n_25), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_274), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_278), .B(n_26), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_276), .Y(n_332) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_282), .B(n_162), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_224), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_235), .B(n_26), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_311), .B(n_236), .Y(n_336) );
INVx4_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_311), .B(n_236), .Y(n_338) );
AND2x6_ASAP7_75t_L g339 ( .A(n_302), .B(n_282), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_296), .B(n_259), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_296), .B(n_259), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_311), .B(n_270), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_291), .B(n_247), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_330), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_296), .B(n_262), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_313), .B(n_268), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_313), .B(n_268), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_313), .B(n_263), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_296), .B(n_272), .Y(n_349) );
NAND2x1_ASAP7_75t_SL g350 ( .A(n_291), .B(n_237), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_330), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_291), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_291), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_313), .B(n_272), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_296), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_294), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_314), .B(n_228), .Y(n_357) );
NOR2xp67_ASAP7_75t_L g358 ( .A(n_291), .B(n_247), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_315), .B(n_228), .Y(n_359) );
NOR2xp33_ASAP7_75t_SL g360 ( .A(n_291), .B(n_248), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_330), .Y(n_361) );
INVx5_ASAP7_75t_L g362 ( .A(n_299), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_330), .B(n_256), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_299), .Y(n_364) );
BUFx4f_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_302), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_337), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_361), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_344), .B(n_315), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_361), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_344), .B(n_315), .Y(n_372) );
INVx3_ASAP7_75t_SL g373 ( .A(n_362), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_366), .Y(n_374) );
INVx5_ASAP7_75t_L g375 ( .A(n_362), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_361), .B(n_298), .Y(n_376) );
INVx6_ASAP7_75t_SL g377 ( .A(n_345), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_366), .A2(n_307), .B1(n_314), .B2(n_331), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_356), .Y(n_379) );
INVx8_ASAP7_75t_L g380 ( .A(n_362), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_366), .B(n_314), .Y(n_382) );
BUFx8_ASAP7_75t_L g383 ( .A(n_355), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_362), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
BUFx4_ASAP7_75t_SL g391 ( .A(n_351), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_362), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_357), .A2(n_237), .B1(n_331), .B2(n_314), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_337), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_391), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_393), .A2(n_357), .B1(n_359), .B2(n_339), .Y(n_399) );
BUFx4f_ASAP7_75t_SL g400 ( .A(n_391), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_357), .B1(n_351), .B2(n_367), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_385), .B(n_357), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_385), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_385), .B(n_351), .Y(n_404) );
CKINVDCx6p67_ASAP7_75t_R g405 ( .A(n_375), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_393), .A2(n_359), .B1(n_339), .B2(n_331), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_370), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_374), .A2(n_300), .B1(n_320), .B2(n_365), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_378), .A2(n_339), .B1(n_331), .B2(n_319), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_378), .A2(n_339), .B1(n_233), .B2(n_300), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_378), .A2(n_339), .B1(n_233), .B2(n_340), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_372), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_374), .A2(n_339), .B1(n_340), .B2(n_341), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
CKINVDCx8_ASAP7_75t_R g421 ( .A(n_375), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
BUFx4f_ASAP7_75t_SL g423 ( .A(n_377), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_369), .Y(n_426) );
INVx6_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_383), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_371), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_371), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_371), .Y(n_431) );
BUFx4f_ASAP7_75t_SL g432 ( .A(n_377), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_382), .A2(n_320), .B1(n_365), .B2(n_301), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_371), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_375), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_394), .B(n_367), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_394), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_379), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_414), .A2(n_382), .B1(n_244), .B2(n_384), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_403), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_403), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_404), .B(n_367), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_402), .B(n_382), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_399), .A2(n_383), .B1(n_339), .B2(n_380), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_414), .A2(n_383), .B1(n_339), .B2(n_380), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_424), .Y(n_449) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_400), .A2(n_244), .B1(n_384), .B2(n_261), .C1(n_225), .C2(n_387), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_417), .A2(n_384), .B1(n_387), .B2(n_375), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_424), .Y(n_452) );
BUFx4f_ASAP7_75t_SL g453 ( .A(n_412), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_416), .A2(n_384), .B1(n_387), .B2(n_375), .Y(n_454) );
BUFx4f_ASAP7_75t_SL g455 ( .A(n_412), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_406), .A2(n_383), .B1(n_339), .B2(n_380), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_401), .A2(n_383), .B1(n_339), .B2(n_380), .Y(n_457) );
INVxp33_ASAP7_75t_SL g458 ( .A(n_435), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_398), .A2(n_261), .B1(n_225), .B2(n_254), .Y(n_462) );
BUFx4f_ASAP7_75t_SL g463 ( .A(n_412), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_402), .B(n_367), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_401), .A2(n_339), .B1(n_380), .B2(n_377), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_398), .A2(n_384), .B1(n_375), .B2(n_392), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_420), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_428), .A2(n_375), .B1(n_392), .B2(n_376), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_433), .A2(n_339), .B1(n_380), .B2(n_377), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_397), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_436), .A2(n_350), .B(n_280), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_405), .A2(n_277), .B1(n_288), .B2(n_279), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_405), .A2(n_375), .B1(n_373), .B2(n_380), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_413), .B(n_277), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_404), .B(n_429), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_430), .A2(n_350), .B(n_292), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_407), .B(n_287), .Y(n_480) );
CKINVDCx11_ASAP7_75t_R g481 ( .A(n_421), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_405), .Y(n_482) );
CKINVDCx14_ASAP7_75t_R g483 ( .A(n_427), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_410), .A2(n_339), .B1(n_377), .B2(n_340), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_410), .A2(n_377), .B1(n_341), .B2(n_340), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_410), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_427), .A2(n_377), .B1(n_340), .B2(n_341), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_407), .A2(n_288), .B1(n_287), .B2(n_348), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_427), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_430), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_427), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_427), .A2(n_341), .B1(n_340), .B2(n_354), .Y(n_493) );
OAI22xp33_ASAP7_75t_SL g494 ( .A1(n_408), .A2(n_395), .B1(n_368), .B2(n_381), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_419), .A2(n_341), .B1(n_340), .B2(n_354), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_422), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_408), .A2(n_341), .B1(n_354), .B2(n_302), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_431), .B(n_392), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_423), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_432), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_431), .A2(n_376), .B(n_333), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_409), .A2(n_375), .B1(n_392), .B2(n_376), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_409), .A2(n_376), .B1(n_373), .B2(n_368), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_422), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_438), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_422), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_411), .A2(n_368), .B1(n_395), .B2(n_381), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_438), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_439), .Y(n_511) );
OAI222xp33_ASAP7_75t_L g512 ( .A1(n_411), .A2(n_395), .B1(n_381), .B2(n_368), .C1(n_302), .C2(n_319), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_476), .A2(n_389), .B1(n_396), .B2(n_388), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_441), .A2(n_389), .B1(n_396), .B2(n_388), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_449), .Y(n_515) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_448), .A2(n_350), .B(n_292), .C(n_295), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_457), .A2(n_418), .B1(n_415), .B2(n_368), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_478), .B(n_415), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_451), .A2(n_389), .B1(n_388), .B2(n_396), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_454), .A2(n_389), .B1(n_388), .B2(n_396), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_465), .A2(n_418), .B1(n_381), .B2(n_368), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_473), .B(n_292), .C(n_158), .Y(n_522) );
OAI222xp33_ASAP7_75t_L g523 ( .A1(n_486), .A2(n_381), .B1(n_395), .B2(n_439), .C1(n_436), .C2(n_426), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_462), .A2(n_295), .B1(n_269), .B2(n_266), .C(n_265), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_458), .A2(n_395), .B1(n_381), .B2(n_364), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_449), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_458), .A2(n_347), .B1(n_346), .B2(n_354), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_447), .A2(n_395), .B1(n_364), .B2(n_373), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_482), .A2(n_319), .B1(n_337), .B2(n_307), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_478), .B(n_426), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_456), .A2(n_364), .B1(n_373), .B2(n_307), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g532 ( .A1(n_494), .A2(n_295), .B(n_319), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_469), .A2(n_364), .B1(n_373), .B2(n_307), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_453), .A2(n_307), .B1(n_337), .B2(n_346), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_452), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g536 ( .A1(n_455), .A2(n_251), .B1(n_337), .B2(n_301), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_450), .A2(n_287), .B1(n_306), .B2(n_288), .C1(n_307), .C2(n_335), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_482), .A2(n_365), .B1(n_307), .B2(n_437), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_463), .A2(n_347), .B1(n_346), .B2(n_341), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_482), .A2(n_365), .B1(n_437), .B2(n_362), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_484), .A2(n_365), .B1(n_437), .B2(n_362), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_491), .B(n_440), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_468), .A2(n_347), .B1(n_346), .B2(n_365), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_483), .A2(n_362), .B1(n_257), .B2(n_329), .Y(n_544) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_479), .A2(n_440), .B(n_329), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_485), .A2(n_329), .B1(n_352), .B2(n_353), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_475), .B(n_360), .Y(n_547) );
OAI222xp33_ASAP7_75t_L g548 ( .A1(n_467), .A2(n_335), .B1(n_440), .B2(n_306), .C1(n_343), .C2(n_353), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_467), .A2(n_347), .B1(n_352), .B2(n_353), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_452), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_488), .A2(n_348), .B1(n_363), .B2(n_336), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_498), .A2(n_363), .B1(n_336), .B2(n_338), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_496), .A2(n_363), .B1(n_345), .B2(n_349), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_445), .A2(n_363), .B1(n_345), .B2(n_349), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_493), .A2(n_363), .B1(n_345), .B2(n_349), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_480), .A2(n_363), .B1(n_345), .B2(n_349), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_470), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_442), .A2(n_271), .B1(n_287), .B2(n_288), .C(n_306), .Y(n_558) );
NAND3xp33_ASAP7_75t_SL g559 ( .A(n_502), .B(n_306), .C(n_335), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_443), .A2(n_289), .B1(n_293), .B2(n_335), .C(n_304), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_511), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_509), .A2(n_338), .B1(n_358), .B2(n_342), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_504), .A2(n_342), .B1(n_345), .B2(n_349), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_489), .A2(n_345), .B1(n_349), .B2(n_358), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g565 ( .A1(n_512), .A2(n_289), .B1(n_293), .B2(n_304), .C1(n_308), .C2(n_316), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_489), .A2(n_349), .B1(n_358), .B2(n_333), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_466), .A2(n_333), .B1(n_323), .B2(n_343), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_492), .A2(n_333), .B1(n_323), .B2(n_343), .Y(n_568) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_472), .A2(n_308), .B(n_322), .Y(n_569) );
OAI222xp33_ASAP7_75t_L g570 ( .A1(n_505), .A2(n_343), .B1(n_304), .B2(n_317), .C1(n_332), .C2(n_324), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_446), .B(n_379), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_487), .A2(n_343), .B1(n_333), .B2(n_323), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_481), .A2(n_323), .B1(n_317), .B2(n_332), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_481), .A2(n_460), .B1(n_444), .B2(n_501), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_444), .B(n_379), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_501), .A2(n_289), .B1(n_293), .B2(n_316), .C(n_308), .Y(n_576) );
AOI221xp5_ASAP7_75t_SL g577 ( .A1(n_503), .A2(n_316), .B1(n_284), .B2(n_241), .C(n_260), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_460), .A2(n_327), .B1(n_324), .B2(n_360), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_470), .B(n_153), .C(n_162), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_460), .A2(n_327), .B1(n_324), .B2(n_360), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_460), .A2(n_327), .B1(n_386), .B2(n_379), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_446), .B(n_379), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_460), .A2(n_390), .B1(n_386), .B2(n_379), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_459), .B(n_379), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_501), .A2(n_390), .B1(n_386), .B2(n_379), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_461), .A2(n_390), .B1(n_386), .B2(n_379), .Y(n_586) );
OAI222xp33_ASAP7_75t_L g587 ( .A1(n_502), .A2(n_290), .B1(n_286), .B2(n_325), .C1(n_303), .C2(n_328), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_500), .A2(n_390), .B1(n_386), .B2(n_290), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_461), .A2(n_390), .B1(n_386), .B2(n_321), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_461), .A2(n_390), .B1(n_386), .B2(n_321), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_459), .B(n_386), .Y(n_591) );
NAND2xp33_ASAP7_75t_SL g592 ( .A(n_500), .B(n_386), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_497), .A2(n_390), .B1(n_321), .B2(n_299), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_497), .A2(n_390), .B1(n_299), .B2(n_321), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_497), .A2(n_390), .B1(n_321), .B2(n_299), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_506), .A2(n_321), .B1(n_299), .B2(n_328), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_506), .A2(n_321), .B1(n_325), .B2(n_303), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_506), .A2(n_321), .B1(n_334), .B2(n_298), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_474), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_464), .A2(n_298), .B1(n_305), .B2(n_318), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_508), .A2(n_321), .B1(n_286), .B2(n_356), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_508), .A2(n_334), .B1(n_305), .B2(n_298), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_508), .A2(n_334), .B1(n_305), .B2(n_298), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_474), .A2(n_298), .B1(n_305), .B2(n_309), .Y(n_604) );
OAI22xp5_ASAP7_75t_SL g605 ( .A1(n_477), .A2(n_286), .B1(n_248), .B2(n_322), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_495), .A2(n_305), .B1(n_356), .B2(n_326), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_499), .A2(n_356), .B1(n_326), .B2(n_310), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_577), .B(n_153), .C(n_158), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_536), .A2(n_510), .B1(n_507), .B2(n_499), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_561), .B(n_507), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_522), .B(n_559), .C(n_524), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_516), .B(n_153), .C(n_158), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_561), .B(n_510), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_542), .B(n_471), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g615 ( .A(n_537), .B(n_490), .C(n_231), .D(n_326), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_518), .B(n_490), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_153), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_514), .A2(n_356), .B1(n_318), .B2(n_312), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_515), .B(n_27), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_515), .B(n_27), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_565), .B(n_153), .C(n_158), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_523), .A2(n_322), .B(n_158), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_526), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_532), .B(n_153), .C(n_158), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_535), .B(n_28), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_576), .B(n_283), .C(n_285), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_563), .A2(n_356), .B1(n_318), .B2(n_312), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_562), .B(n_153), .C(n_158), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_550), .B(n_28), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_550), .B(n_29), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_557), .B(n_158), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_557), .B(n_29), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_529), .B(n_162), .C(n_154), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_599), .B(n_30), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_530), .B(n_31), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_575), .B(n_32), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_563), .B(n_32), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_558), .B(n_283), .C(n_285), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_574), .B(n_162), .C(n_154), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_571), .B(n_34), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_517), .B(n_34), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_571), .B(n_162), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_582), .B(n_162), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_582), .B(n_35), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_552), .B(n_35), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_584), .B(n_36), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_525), .A2(n_356), .B1(n_318), .B2(n_312), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_584), .B(n_36), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_549), .B(n_162), .C(n_154), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_591), .B(n_39), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_552), .B(n_309), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_543), .B(n_255), .C(n_258), .D(n_276), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_548), .A2(n_246), .B(n_318), .Y(n_653) );
NAND2x1_ASAP7_75t_L g654 ( .A(n_540), .B(n_356), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_591), .B(n_43), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_527), .A2(n_312), .B1(n_297), .B2(n_309), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_513), .B(n_154), .C(n_309), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_519), .B(n_44), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_545), .B(n_154), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_570), .A2(n_246), .B(n_309), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_594), .A2(n_297), .B(n_258), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_551), .B(n_297), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_551), .B(n_297), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_521), .B(n_297), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_560), .A2(n_154), .B1(n_285), .B2(n_294), .C(n_310), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_547), .A2(n_285), .B(n_294), .C(n_310), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_579), .B(n_310), .C(n_294), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_527), .A2(n_285), .B1(n_253), .B2(n_310), .C(n_294), .Y(n_668) );
AND2x2_ASAP7_75t_SL g669 ( .A(n_545), .B(n_285), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g670 ( .A1(n_538), .A2(n_253), .B(n_294), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_546), .A2(n_310), .B1(n_294), .B2(n_226), .C(n_49), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_588), .B(n_310), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_541), .A2(n_310), .B1(n_294), .B2(n_47), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_600), .B(n_294), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_592), .B(n_310), .C(n_50), .Y(n_675) );
NAND4xp25_ASAP7_75t_L g676 ( .A(n_534), .B(n_46), .C(n_51), .D(n_54), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_586), .B(n_55), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_592), .B(n_56), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_520), .B(n_57), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_569), .B(n_59), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_569), .B(n_61), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_604), .B(n_62), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_553), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_569), .B(n_585), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_604), .B(n_67), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_583), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g687 ( .A1(n_531), .A2(n_69), .B(n_71), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_607), .B(n_72), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_589), .B(n_73), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_605), .B(n_76), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_606), .B(n_78), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_590), .B(n_79), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_544), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_601), .B(n_80), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_581), .B(n_81), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_528), .B(n_82), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_578), .B(n_85), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_533), .B(n_89), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_554), .A2(n_90), .B1(n_92), .B2(n_93), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_564), .A2(n_96), .B1(n_98), .B2(n_99), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_580), .B(n_100), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_539), .B(n_103), .C(n_104), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_609), .B(n_572), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_614), .B(n_556), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_614), .B(n_555), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_693), .B(n_587), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_684), .B(n_595), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_669), .B(n_567), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_684), .B(n_593), .Y(n_709) );
OA21x2_ASAP7_75t_L g710 ( .A1(n_686), .A2(n_566), .B(n_573), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_611), .B(n_598), .C(n_568), .Y(n_711) );
NAND4xp75_ASAP7_75t_L g712 ( .A(n_694), .B(n_596), .C(n_597), .D(n_602), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_635), .B(n_603), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_622), .B(n_105), .C(n_621), .Y(n_714) );
BUFx3_ASAP7_75t_L g715 ( .A(n_617), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_615), .B(n_637), .C(n_645), .D(n_652), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_613), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_641), .A2(n_636), .B1(n_630), .B2(n_625), .C(n_634), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_616), .B(n_623), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_690), .B(n_639), .C(n_687), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_690), .B(n_676), .C(n_694), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_657), .B(n_633), .C(n_629), .Y(n_722) );
AO22x1_ASAP7_75t_L g723 ( .A1(n_640), .A2(n_644), .B1(n_646), .B2(n_648), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_642), .B(n_643), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_653), .B(n_670), .C(n_612), .Y(n_725) );
NAND4xp75_ASAP7_75t_L g726 ( .A(n_678), .B(n_689), .C(n_680), .D(n_681), .Y(n_726) );
OR2x2_ASAP7_75t_SL g727 ( .A(n_675), .B(n_628), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_660), .A2(n_661), .B1(n_654), .B2(n_627), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_631), .B(n_659), .Y(n_729) );
NAND4xp75_ASAP7_75t_L g730 ( .A(n_678), .B(n_689), .C(n_701), .D(n_658), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g731 ( .A(n_619), .B(n_620), .C(n_632), .Y(n_731) );
NAND4xp75_ASAP7_75t_L g732 ( .A(n_701), .B(n_696), .C(n_671), .D(n_698), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_651), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_650), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_672), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_655), .B(n_664), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_696), .B(n_698), .C(n_679), .D(n_677), .Y(n_737) );
NAND3xp33_ASAP7_75t_SL g738 ( .A(n_626), .B(n_666), .C(n_683), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_662), .B(n_663), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_677), .B(n_674), .Y(n_740) );
AO21x2_ASAP7_75t_L g741 ( .A1(n_608), .A2(n_624), .B(n_667), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_649), .B(n_683), .C(n_699), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_656), .B(n_618), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_647), .B(n_697), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_702), .A2(n_699), .B(n_668), .Y(n_745) );
AOI221x1_ASAP7_75t_L g746 ( .A1(n_697), .A2(n_692), .B1(n_688), .B2(n_685), .C(n_682), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_697), .B(n_691), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_665), .B(n_638), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_695), .B(n_673), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_695), .B(n_700), .Y(n_750) );
NOR2x1_ASAP7_75t_L g751 ( .A(n_622), .B(n_653), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_609), .B(n_611), .C(n_622), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_621), .B(n_450), .C(n_690), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_611), .A2(n_615), .B1(n_476), .B2(n_693), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_610), .B(n_613), .Y(n_755) );
NAND4xp75_ASAP7_75t_L g756 ( .A(n_694), .B(n_690), .C(n_398), .D(n_684), .Y(n_756) );
OR2x2_ASAP7_75t_SL g757 ( .A(n_693), .B(n_486), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_609), .B(n_611), .C(n_622), .Y(n_758) );
NAND4xp75_ASAP7_75t_L g759 ( .A(n_694), .B(n_690), .C(n_398), .D(n_684), .Y(n_759) );
INVx3_ASAP7_75t_L g760 ( .A(n_654), .Y(n_760) );
AND2x4_ASAP7_75t_SL g761 ( .A(n_614), .B(n_482), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_610), .B(n_613), .Y(n_762) );
AOI21x1_ASAP7_75t_L g763 ( .A1(n_690), .A2(n_694), .B(n_678), .Y(n_763) );
NAND4xp75_ASAP7_75t_L g764 ( .A(n_694), .B(n_690), .C(n_398), .D(n_684), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_614), .B(n_684), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_728), .B(n_760), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_752), .B(n_758), .C(n_728), .Y(n_767) );
NAND4xp75_ASAP7_75t_SL g768 ( .A(n_763), .B(n_706), .C(n_710), .D(n_747), .Y(n_768) );
NAND4xp75_ASAP7_75t_SL g769 ( .A(n_706), .B(n_710), .C(n_747), .D(n_759), .Y(n_769) );
INVx1_ASAP7_75t_SL g770 ( .A(n_761), .Y(n_770) );
XOR2x2_ASAP7_75t_L g771 ( .A(n_723), .B(n_712), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_760), .B(n_761), .Y(n_772) );
AND2x4_ASAP7_75t_SL g773 ( .A(n_721), .B(n_729), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_707), .B(n_709), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_765), .B(n_755), .Y(n_775) );
OR2x2_ASAP7_75t_L g776 ( .A(n_762), .B(n_717), .Y(n_776) );
NAND4xp75_ASAP7_75t_L g777 ( .A(n_751), .B(n_703), .C(n_745), .D(n_746), .Y(n_777) );
NAND4xp75_ASAP7_75t_SL g778 ( .A(n_710), .B(n_764), .C(n_756), .D(n_753), .Y(n_778) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_738), .B(n_703), .C(n_711), .Y(n_779) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_757), .B(n_754), .Y(n_780) );
NAND3xp33_ASAP7_75t_SL g781 ( .A(n_720), .B(n_754), .C(n_725), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_719), .Y(n_782) );
XNOR2xp5_ASAP7_75t_L g783 ( .A(n_737), .B(n_726), .Y(n_783) );
XNOR2xp5_ASAP7_75t_L g784 ( .A(n_716), .B(n_730), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_715), .Y(n_785) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_715), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_760), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_735), .B(n_733), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_739), .B(n_735), .Y(n_789) );
NAND4xp75_ASAP7_75t_L g790 ( .A(n_708), .B(n_718), .C(n_749), .D(n_750), .Y(n_790) );
XOR2x2_ASAP7_75t_L g791 ( .A(n_732), .B(n_742), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_724), .B(n_705), .Y(n_792) );
XNOR2x2_ASAP7_75t_L g793 ( .A(n_714), .B(n_708), .Y(n_793) );
XOR2x2_ASAP7_75t_L g794 ( .A(n_734), .B(n_731), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_729), .Y(n_795) );
XOR2x2_ASAP7_75t_L g796 ( .A(n_734), .B(n_704), .Y(n_796) );
INVx1_ASAP7_75t_SL g797 ( .A(n_770), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_788), .Y(n_798) );
BUFx2_ASAP7_75t_L g799 ( .A(n_772), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_772), .Y(n_800) );
XOR2x2_ASAP7_75t_L g801 ( .A(n_771), .B(n_713), .Y(n_801) );
XNOR2xp5_ASAP7_75t_L g802 ( .A(n_771), .B(n_736), .Y(n_802) );
XOR2x2_ASAP7_75t_L g803 ( .A(n_791), .B(n_713), .Y(n_803) );
XNOR2x1_ASAP7_75t_L g804 ( .A(n_791), .B(n_743), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_788), .Y(n_805) );
INVx1_ASAP7_75t_SL g806 ( .A(n_772), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_789), .Y(n_807) );
INVxp67_ASAP7_75t_L g808 ( .A(n_781), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_795), .Y(n_809) );
XNOR2xp5_ASAP7_75t_L g810 ( .A(n_783), .B(n_736), .Y(n_810) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_784), .B(n_748), .Y(n_811) );
INVx1_ASAP7_75t_SL g812 ( .A(n_773), .Y(n_812) );
INVx1_ASAP7_75t_SL g813 ( .A(n_773), .Y(n_813) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_766), .B(n_741), .Y(n_814) );
XNOR2x1_ASAP7_75t_L g815 ( .A(n_784), .B(n_744), .Y(n_815) );
INVx1_ASAP7_75t_SL g816 ( .A(n_794), .Y(n_816) );
XNOR2x2_ASAP7_75t_L g817 ( .A(n_777), .B(n_727), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_786), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_775), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_783), .B(n_740), .Y(n_820) );
XOR2x2_ASAP7_75t_L g821 ( .A(n_780), .B(n_722), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_775), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_792), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_818), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_817), .A2(n_793), .B1(n_767), .B2(n_768), .Y(n_825) );
INVx4_ASAP7_75t_L g826 ( .A(n_799), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_798), .Y(n_827) );
OA22x2_ASAP7_75t_L g828 ( .A1(n_816), .A2(n_780), .B1(n_777), .B2(n_778), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_801), .B(n_790), .Y(n_829) );
XOR2x2_ASAP7_75t_L g830 ( .A(n_801), .B(n_790), .Y(n_830) );
INVx1_ASAP7_75t_SL g831 ( .A(n_797), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_805), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_809), .Y(n_833) );
BUFx3_ASAP7_75t_L g834 ( .A(n_817), .Y(n_834) );
OAI22x1_ASAP7_75t_L g835 ( .A1(n_802), .A2(n_794), .B1(n_787), .B2(n_785), .Y(n_835) );
OA22x2_ASAP7_75t_L g836 ( .A1(n_808), .A2(n_769), .B1(n_779), .B2(n_774), .Y(n_836) );
OAI22x1_ASAP7_75t_L g837 ( .A1(n_808), .A2(n_785), .B1(n_796), .B2(n_776), .Y(n_837) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_812), .Y(n_838) );
AO22x2_ASAP7_75t_L g839 ( .A1(n_804), .A2(n_776), .B1(n_782), .B2(n_792), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_824), .Y(n_840) );
XOR2xp5_ASAP7_75t_L g841 ( .A(n_829), .B(n_804), .Y(n_841) );
OAI322xp33_ASAP7_75t_L g842 ( .A1(n_828), .A2(n_815), .A3(n_813), .B1(n_820), .B2(n_810), .C1(n_800), .C2(n_806), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g843 ( .A(n_831), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_838), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_838), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_826), .Y(n_846) );
BUFx2_ASAP7_75t_L g847 ( .A(n_826), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_842), .A2(n_834), .B1(n_839), .B2(n_837), .C(n_835), .Y(n_848) );
AOI31xp33_ASAP7_75t_L g849 ( .A1(n_841), .A2(n_825), .A3(n_814), .B(n_815), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_845), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_845), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_844), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_848), .A2(n_828), .B1(n_830), .B2(n_834), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_851), .A2(n_836), .B1(n_825), .B2(n_839), .Y(n_854) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_850), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_853), .A2(n_836), .B1(n_843), .B2(n_839), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_854), .A2(n_843), .B1(n_821), .B2(n_846), .Y(n_857) );
NOR2x1_ASAP7_75t_L g858 ( .A(n_856), .B(n_847), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_857), .A2(n_847), .B1(n_821), .B2(n_811), .Y(n_859) );
OAI22x1_ASAP7_75t_L g860 ( .A1(n_859), .A2(n_855), .B1(n_852), .B2(n_850), .Y(n_860) );
NOR2x1_ASAP7_75t_L g861 ( .A(n_858), .B(n_849), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_860), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_861), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_863), .A2(n_811), .B1(n_803), .B2(n_840), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_864), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_865), .A2(n_862), .B1(n_840), .B2(n_803), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_866), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_867), .A2(n_833), .B1(n_832), .B2(n_827), .Y(n_868) );
INVx1_ASAP7_75t_SL g869 ( .A(n_868), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_869), .A2(n_833), .B1(n_832), .B2(n_827), .C(n_823), .Y(n_870) );
AOI211xp5_ASAP7_75t_L g871 ( .A1(n_870), .A2(n_822), .B(n_819), .C(n_807), .Y(n_871) );
endmodule