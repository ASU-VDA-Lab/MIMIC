module real_jpeg_19033_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_37),
.B1(n_50),
.B2(n_53),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_0),
.A2(n_37),
.B1(n_66),
.B2(n_67),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_1),
.A2(n_44),
.B1(n_66),
.B2(n_67),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_44),
.B1(n_50),
.B2(n_53),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_31),
.B(n_34),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_2),
.B(n_101),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_53),
.B(n_84),
.C(n_153),
.D(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_2),
.B(n_53),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_2),
.B(n_49),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_69),
.B(n_168),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_33),
.B(n_46),
.C(n_55),
.D(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_33),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_3),
.A2(n_66),
.B1(n_67),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_50),
.B1(n_53),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_82),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_7),
.B(n_169),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_9),
.A2(n_29),
.B1(n_50),
.B2(n_53),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_9),
.A2(n_29),
.B1(n_66),
.B2(n_67),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_50),
.B1(n_53),
.B2(n_72),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_12),
.A2(n_50),
.B1(n_53),
.B2(n_68),
.Y(n_89)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_105),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_91),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_22),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_41),
.B1(n_42),
.B2(n_58),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_25),
.A2(n_30),
.B1(n_39),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_30),
.B(n_32),
.C(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_32),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_32),
.B(n_62),
.C(n_63),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_36),
.B(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_38),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_41),
.B(n_58),
.C(n_59),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_54),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_43),
.A2(n_45),
.B1(n_57),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_46),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_48),
.Y(n_208)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_85),
.B(n_86),
.C(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_50),
.B(n_52),
.Y(n_207)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_53),
.A2(n_202),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_57),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_57),
.A2(n_104),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

AOI22x1_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_62),
.B(n_90),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_62),
.B(n_70),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_64),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_67),
.B1(n_85),
.B2(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_66),
.B(n_85),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_66),
.B(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_67),
.A2(n_86),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_70),
.B1(n_78),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_69),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_69),
.B(n_170),
.Y(n_186)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_70),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_70),
.A2(n_175),
.B(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_91),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_80),
.Y(n_115)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_77),
.A2(n_186),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_90),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_83),
.A2(n_90),
.B1(n_165),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_83),
.A2(n_200),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_95),
.Y(n_94)
);

CKINVDCx9p33_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_96),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_90),
.A2(n_94),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_102),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_93),
.B1(n_102),
.B2(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_126),
.B2(n_127),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_126),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_146),
.B(n_231),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_144),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_131),
.B(n_144),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_132),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_134),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_138),
.A2(n_139),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_140),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_225),
.B(n_230),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_213),
.B(n_224),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_194),
.B(n_212),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_171),
.B(n_193),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_159),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_151),
.B(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_155),
.B1(n_156),
.B2(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_181),
.B(n_192),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_179),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_187),
.B(n_191),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_184),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_205),
.B2(n_211),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_199),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_204),
.C(n_211),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_209),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_221),
.C(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);


endmodule