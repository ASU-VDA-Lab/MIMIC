module fake_jpeg_18996_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_2),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_9),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_19),
.B1(n_7),
.B2(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_17),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_19),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_14),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.C(n_30),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_22),
.C(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_22),
.C(n_23),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

OAI21x1_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_37),
.B(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_10),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_25),
.C(n_21),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_35),
.C(n_7),
.Y(n_42)
);

AOI31xp67_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.A3(n_11),
.B(n_20),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.A3(n_11),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_0),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_3),
.B(n_1),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);


endmodule