module fake_jpeg_2621_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_29),
.B(n_1),
.C(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_8),
.Y(n_25)
);

INVx5_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_1),
.B1(n_7),
.B2(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_28),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_37),
.C(n_17),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_17),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_45),
.B1(n_35),
.B2(n_21),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_45),
.A3(n_48),
.B1(n_19),
.B2(n_47),
.C1(n_31),
.C2(n_27),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_53),
.B(n_50),
.Y(n_54)
);


endmodule