module real_jpeg_21421_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_0),
.A2(n_10),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_0),
.A2(n_19),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_10),
.B1(n_13),
.B2(n_18),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_4),
.B(n_18),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_3),
.A2(n_13),
.B1(n_36),
.B2(n_40),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_4),
.A2(n_10),
.B1(n_18),
.B2(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_4),
.A2(n_28),
.B1(n_36),
.B2(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_30),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_24),
.B(n_29),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_14),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_11),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_18),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_12),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_28),
.B(n_35),
.C(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_32),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B(n_21),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_47),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_46),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B(n_42),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);


endmodule