module real_jpeg_32519_n_13 (n_123, n_8, n_116, n_0, n_2, n_125, n_10, n_9, n_12, n_124, n_6, n_121, n_11, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_120, n_13);

input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_125;
input n_10;
input n_9;
input n_12;
input n_124;
input n_6;
input n_121;
input n_11;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_120;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_0),
.B(n_28),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_3),
.B1(n_44),
.B2(n_51),
.C(n_56),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_44),
.C(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_78),
.A3(n_80),
.B1(n_86),
.B2(n_108),
.C1(n_110),
.C2(n_125),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_5),
.B(n_88),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_7),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_8),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_8),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_12),
.B(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_24),
.B2(n_113),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_70),
.B(n_103),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_36),
.B(n_69),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_60),
.B(n_68),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_118),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR4xp25_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_85),
.C(n_94),
.D(n_99),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_104),
.B(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_99),
.C(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_121),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OA21x2_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_115),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_116),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_117),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_119),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_120),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_122),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_123),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_124),
.Y(n_101)
);


endmodule