module fake_jpeg_26889_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_70),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_63),
.B1(n_55),
.B2(n_47),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_49),
.B1(n_58),
.B2(n_53),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_47),
.B1(n_55),
.B2(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_50),
.B1(n_51),
.B2(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_83),
.B1(n_58),
.B2(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_60),
.B1(n_56),
.B2(n_57),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_93),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_46),
.C(n_59),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_96),
.C(n_99),
.Y(n_108)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_17),
.A3(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_13),
.B1(n_35),
.B2(n_33),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_15),
.B(n_42),
.Y(n_104)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_12),
.C(n_32),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_106),
.Y(n_109)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_93),
.B1(n_98),
.B2(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_81),
.B1(n_80),
.B2(n_94),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_95),
.B(n_99),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_97),
.B(n_6),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_120),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_108),
.C(n_101),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_128),
.C(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_29),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_3),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_3),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_5),
.B(n_6),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_130),
.B1(n_5),
.B2(n_7),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_27),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_28),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_26),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_135),
.C(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_23),
.C(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_25),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_130),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_133),
.C(n_141),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_146),
.B1(n_132),
.B2(n_144),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_132),
.B(n_118),
.Y(n_146)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_148),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_142),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_131),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_136),
.C(n_121),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);


endmodule