module fake_ibex_1973_n_1187 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_132, n_174, n_210, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1187);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_132;
input n_174;
input n_210;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1187;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_1148;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_510;
wire n_256;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1044;
wire n_1106;
wire n_1018;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1138;
wire n_727;
wire n_1134;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_647;
wire n_531;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_698;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1112;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_732;
wire n_673;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1068;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_787;
wire n_694;
wire n_1075;
wire n_1136;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_1168;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_933;
wire n_1081;
wire n_215;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_669;
wire n_538;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_1082;
wire n_1137;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_1180;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_1171;
wire n_438;
wire n_851;
wire n_1028;
wire n_1012;
wire n_993;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_234;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_439;
wire n_262;
wire n_704;
wire n_949;
wire n_1126;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_955;
wire n_1170;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1057;
wire n_1049;
wire n_763;
wire n_1086;
wire n_745;
wire n_1158;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_562;
wire n_444;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_1160;
wire n_615;
wire n_512;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_283;
wire n_366;
wire n_803;
wire n_894;
wire n_1118;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_288;
wire n_379;
wire n_247;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_977;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1095;
wire n_361;
wire n_1085;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1102;
wire n_1005;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_1150;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_912;
wire n_921;
wire n_890;
wire n_874;
wire n_1105;
wire n_1058;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_565;
wire n_424;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_1000;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1038;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_1186;
wire n_657;
wire n_764;
wire n_1156;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_63),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_89),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_67),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_26),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_39),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_184),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_76),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_115),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_112),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_49),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_85),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_70),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_38),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_27),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_81),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_109),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_125),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_57),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_29),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_117),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_203),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_71),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_102),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_161),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_126),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_90),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_65),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_54),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_120),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_167),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_38),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_31),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_133),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_169),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_140),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_55),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_20),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_36),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_141),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_26),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_180),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_162),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_134),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_155),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_96),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_146),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_170),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_45),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_156),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_147),
.B(n_75),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_86),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_187),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_139),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_178),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_84),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_107),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_188),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_16),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_61),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_106),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_72),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_110),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_73),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_195),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_33),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_186),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_128),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_52),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_20),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_59),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_157),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_193),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_100),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_42),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_99),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_91),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_113),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_37),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_132),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_31),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_104),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_148),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_137),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_142),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_64),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_19),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_208),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_191),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_58),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_127),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_114),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_97),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_196),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_181),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_24),
.B(n_123),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_204),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_17),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_2),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_30),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_168),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_32),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_88),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_135),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_62),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_122),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_48),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_3),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_46),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_93),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_13),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_214),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_124),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_3),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_24),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_98),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_12),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_29),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_216),
.Y(n_364)
);

OAI21x1_ASAP7_75t_L g365 ( 
.A1(n_218),
.A2(n_80),
.B(n_206),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_293),
.B(n_0),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g367 ( 
.A1(n_218),
.A2(n_77),
.B(n_205),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_216),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_274),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_227),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_216),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_222),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_222),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_255),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_239),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_255),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_239),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_255),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_278),
.B(n_4),
.Y(n_382)
);

BUFx8_ASAP7_75t_L g383 ( 
.A(n_255),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_359),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_270),
.A2(n_87),
.B(n_199),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_271),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_6),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_255),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_8),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_335),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_255),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_238),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_238),
.B(n_9),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_345),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_270),
.A2(n_103),
.B(n_198),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_219),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_275),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_346),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_275),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_216),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_299),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_300),
.B(n_13),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_287),
.A2(n_357),
.B(n_350),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_278),
.B(n_15),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_299),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_287),
.A2(n_105),
.B(n_197),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_217),
.Y(n_416)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_301),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_345),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_237),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_220),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_252),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_22),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_229),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_350),
.A2(n_118),
.B(n_194),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_231),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_232),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_315),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_235),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_301),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_315),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_241),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_243),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_269),
.B(n_23),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_277),
.B(n_286),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_322),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_244),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_234),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_329),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_248),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_329),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_245),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_290),
.B(n_25),
.Y(n_442)
);

CKINVDCx6p67_ASAP7_75t_R g443 ( 
.A(n_301),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_322),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_226),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_266),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_246),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_322),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_322),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_357),
.A2(n_119),
.B(n_192),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_302),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_250),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_254),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_226),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_257),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_258),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_259),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_249),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_261),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_314),
.B(n_319),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_332),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_383),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_370),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_395),
.A2(n_343),
.B1(n_344),
.B2(n_354),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_L g465 ( 
.A(n_386),
.B(n_362),
.C(n_289),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_409),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_409),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_375),
.B(n_304),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_383),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_395),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_376),
.A2(n_353),
.B1(n_253),
.B2(n_340),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_L g477 ( 
.A(n_401),
.B(n_215),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_408),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_383),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_364),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_383),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_373),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_416),
.B(n_264),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_373),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_406),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_373),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_455),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_387),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_372),
.Y(n_496)
);

BUFx6f_ASAP7_75t_SL g497 ( 
.A(n_375),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_416),
.A2(n_356),
.B1(n_323),
.B2(n_310),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_372),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_377),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_377),
.Y(n_504)
);

BUFx6f_ASAP7_75t_SL g505 ( 
.A(n_375),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_412),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_420),
.B(n_265),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_389),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_399),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_382),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_420),
.B(n_267),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_397),
.B(n_215),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_364),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_455),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_399),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_417),
.B(n_341),
.Y(n_520)
);

INVx11_ASAP7_75t_L g521 ( 
.A(n_417),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_411),
.B(n_369),
.C(n_375),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_423),
.A2(n_313),
.B1(n_298),
.B2(n_355),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_422),
.B(n_309),
.C(n_280),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_429),
.B(n_338),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_370),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_455),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_429),
.B(n_339),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_445),
.B(n_253),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_410),
.B(n_326),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_423),
.A2(n_312),
.B1(n_279),
.B2(n_352),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_443),
.B(n_233),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_451),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_438),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_458),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_425),
.A2(n_268),
.B1(n_283),
.B2(n_351),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_410),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_461),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_429),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_425),
.B(n_426),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_427),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_376),
.B(n_418),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_439),
.B(n_233),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_426),
.B(n_272),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_440),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_418),
.A2(n_353),
.B1(n_337),
.B2(n_340),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_428),
.B(n_282),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_446),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_384),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_430),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_431),
.B(n_348),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_431),
.B(n_432),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_422),
.B(n_285),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_432),
.B(n_436),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_374),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_364),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_436),
.B(n_295),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_364),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_452),
.Y(n_570)
);

INVx6_ASAP7_75t_L g571 ( 
.A(n_458),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_441),
.A2(n_303),
.B1(n_330),
.B2(n_331),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_374),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_364),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_441),
.B(n_242),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_440),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_378),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_385),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_378),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_456),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_380),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_447),
.B(n_347),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_447),
.B(n_360),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_380),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_SL g587 ( 
.A1(n_379),
.A2(n_263),
.B1(n_273),
.B2(n_296),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_453),
.A2(n_325),
.B1(n_320),
.B2(n_317),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_368),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_453),
.B(n_221),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_368),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_385),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_457),
.B(n_306),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_457),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_459),
.A2(n_333),
.B1(n_336),
.B2(n_358),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_393),
.B(n_223),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_381),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_365),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_381),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_393),
.B(n_225),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_434),
.B(n_292),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_388),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_388),
.B(n_228),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_460),
.B(n_458),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_392),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_392),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_400),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_400),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_368),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_379),
.A2(n_288),
.B1(n_316),
.B2(n_337),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_402),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_394),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_402),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_393),
.B(n_230),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_394),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_458),
.B(n_236),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_405),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_405),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_404),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_404),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_458),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_413),
.Y(n_623)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_558),
.B(n_458),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_559),
.B(n_494),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_510),
.B(n_390),
.Y(n_626)
);

OAI221xp5_ASAP7_75t_L g627 ( 
.A1(n_464),
.A2(n_433),
.B1(n_442),
.B2(n_396),
.C(n_391),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_466),
.A2(n_365),
.B(n_450),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_587),
.A2(n_421),
.B(n_419),
.C(n_366),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_575),
.B(n_470),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_562),
.A2(n_435),
.B(n_407),
.C(n_449),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_520),
.B(n_367),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_522),
.B(n_470),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_526),
.B(n_413),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_549),
.B(n_414),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_544),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_464),
.A2(n_513),
.B1(n_471),
.B2(n_474),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_535),
.Y(n_638)
);

AND2x6_ASAP7_75t_SL g639 ( 
.A(n_552),
.B(n_414),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_611),
.B(n_556),
.C(n_476),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_563),
.A2(n_288),
.B1(n_321),
.B2(n_316),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_462),
.B(n_407),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_549),
.B(n_240),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_519),
.B(n_445),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_472),
.B(n_435),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_535),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_544),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_549),
.B(n_247),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_479),
.B(n_251),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_543),
.B(n_454),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_560),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_256),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_561),
.B(n_260),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_561),
.B(n_262),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_529),
.B(n_276),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_483),
.B(n_281),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_584),
.B(n_291),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_585),
.B(n_294),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_534),
.B(n_297),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_492),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_563),
.A2(n_321),
.B1(n_396),
.B2(n_454),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_473),
.A2(n_449),
.B1(n_448),
.B2(n_444),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_563),
.A2(n_444),
.B1(n_448),
.B2(n_349),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_536),
.B(n_602),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_497),
.B(n_305),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_469),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_602),
.B(n_318),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_532),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_516),
.B(n_327),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_497),
.B(n_328),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_466),
.B(n_467),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_537),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_553),
.B(n_334),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_550),
.B(n_385),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_550),
.B(n_415),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_547),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_467),
.A2(n_450),
.B(n_367),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_545),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_546),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_544),
.B(n_398),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_505),
.B(n_415),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_565),
.B(n_424),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_521),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_525),
.B(n_403),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_475),
.B(n_403),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_465),
.B(n_477),
.C(n_485),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_489),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_520),
.B(n_403),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_468),
.B(n_371),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_491),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_478),
.B(n_403),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_468),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_480),
.B(n_371),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_551),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_488),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_605),
.B(n_28),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_596),
.B(n_30),
.C(n_32),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_520),
.B(n_33),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_463),
.B(n_34),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_597),
.B(n_34),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_601),
.B(n_37),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_480),
.B(n_129),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_480),
.B(n_130),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_615),
.B(n_40),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_527),
.B(n_40),
.Y(n_708)
);

NOR2x1p5_ASAP7_75t_L g709 ( 
.A(n_527),
.B(n_41),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_488),
.B(n_41),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_604),
.B(n_131),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_570),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_596),
.B(n_143),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_580),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_484),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_604),
.B(n_144),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_477),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_524),
.B(n_43),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_524),
.B(n_44),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_L g720 ( 
.A(n_484),
.B(n_46),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_484),
.Y(n_721)
);

AND2x4_ASAP7_75t_SL g722 ( 
.A(n_552),
.B(n_47),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_599),
.A2(n_150),
.B(n_50),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_608),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_582),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_594),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_484),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_533),
.B(n_47),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_595),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_533),
.B(n_51),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_498),
.A2(n_53),
.B1(n_56),
.B2(n_60),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_552),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_485),
.B(n_74),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_508),
.B(n_82),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_508),
.B(n_92),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_493),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_541),
.B(n_94),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_496),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_498),
.B(n_101),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_541),
.B(n_108),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_514),
.B(n_111),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_599),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_572),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_669),
.B(n_530),
.Y(n_744)
);

INVx8_ASAP7_75t_L g745 ( 
.A(n_691),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_669),
.B(n_514),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_672),
.A2(n_579),
.B(n_592),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_625),
.B(n_572),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_678),
.A2(n_592),
.B(n_579),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_682),
.B(n_588),
.C(n_592),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_633),
.A2(n_501),
.B(n_502),
.C(n_504),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_684),
.B(n_588),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_633),
.A2(n_507),
.B(n_509),
.C(n_621),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_672),
.A2(n_554),
.B(n_557),
.Y(n_754)
);

NAND2x1p5_ASAP7_75t_L g755 ( 
.A(n_636),
.B(n_609),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_742),
.B(n_593),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_695),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_660),
.B(n_612),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_626),
.B(n_554),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_692),
.A2(n_557),
.B(n_568),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_627),
.A2(n_637),
.B(n_629),
.C(n_718),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_692),
.A2(n_568),
.B(n_586),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_647),
.B(n_617),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_691),
.B(n_622),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_626),
.B(n_614),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_675),
.A2(n_581),
.B(n_583),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_676),
.A2(n_581),
.B(n_583),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_695),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_683),
.A2(n_606),
.B(n_586),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_689),
.A2(n_593),
.B1(n_617),
.B2(n_623),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_644),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_738),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_641),
.A2(n_620),
.B1(n_603),
.B2(n_566),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_691),
.Y(n_774)
);

BUFx12f_ASAP7_75t_L g775 ( 
.A(n_639),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_685),
.B(n_593),
.Y(n_776)
);

AO32x1_ASAP7_75t_L g777 ( 
.A1(n_731),
.A2(n_538),
.A3(n_531),
.B1(n_539),
.B2(n_523),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_724),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_660),
.B(n_153),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_689),
.A2(n_566),
.B1(n_573),
.B2(n_578),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_719),
.A2(n_619),
.B(n_618),
.C(n_616),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_630),
.A2(n_573),
.B1(n_566),
.B2(n_607),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_628),
.A2(n_613),
.B(n_598),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_742),
.B(n_603),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_685),
.B(n_540),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_634),
.B(n_573),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_650),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_634),
.A2(n_578),
.B(n_607),
.C(n_600),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_682),
.A2(n_616),
.B(n_613),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_642),
.A2(n_600),
.B(n_506),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_642),
.A2(n_506),
.B(n_523),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_665),
.B(n_571),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_661),
.Y(n_793)
);

INVx11_ASAP7_75t_L g794 ( 
.A(n_709),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_659),
.B(n_528),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_635),
.B(n_528),
.Y(n_796)
);

BUFx8_ASAP7_75t_L g797 ( 
.A(n_701),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_631),
.A2(n_500),
.B(n_577),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_499),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_727),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_670),
.B(n_499),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_645),
.A2(n_531),
.B(n_512),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_728),
.A2(n_518),
.B(n_499),
.C(n_515),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_645),
.A2(n_490),
.B(n_512),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_732),
.B(n_490),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_708),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_681),
.B(n_515),
.C(n_518),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_712),
.B(n_486),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_714),
.B(n_486),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_725),
.B(n_487),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_624),
.B(n_487),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_695),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_643),
.B(n_542),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_677),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_632),
.A2(n_555),
.B(n_481),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_632),
.A2(n_564),
.B(n_503),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_673),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_715),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_632),
.A2(n_564),
.B(n_503),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_733),
.A2(n_548),
.B(n_495),
.C(n_538),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_640),
.B(n_576),
.Y(n_822)
);

AO21x1_ASAP7_75t_L g823 ( 
.A1(n_732),
.A2(n_548),
.B(n_159),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_715),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_648),
.B(n_663),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_722),
.B(n_610),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_695),
.A2(n_739),
.B1(n_740),
.B2(n_698),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_668),
.B(n_154),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_726),
.B(n_729),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_674),
.B(n_160),
.C(n_163),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_733),
.A2(n_610),
.B(n_591),
.C(n_589),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_653),
.B(n_164),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_654),
.B(n_166),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_657),
.B(n_171),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_658),
.B(n_172),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_652),
.B(n_482),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_710),
.A2(n_173),
.B(n_174),
.C(n_175),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_666),
.B(n_179),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_662),
.A2(n_517),
.B(n_574),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_666),
.Y(n_840)
);

O2A1O1Ixp5_ASAP7_75t_SL g841 ( 
.A1(n_705),
.A2(n_706),
.B(n_686),
.C(n_713),
.Y(n_841)
);

OAI321xp33_ASAP7_75t_L g842 ( 
.A1(n_717),
.A2(n_482),
.A3(n_567),
.B1(n_569),
.B2(n_574),
.C(n_591),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_671),
.B(n_189),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_655),
.B(n_213),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_667),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_679),
.B(n_569),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_702),
.B(n_680),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_690),
.B(n_693),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_703),
.B(n_704),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_698),
.A2(n_662),
.B1(n_700),
.B2(n_737),
.Y(n_850)
);

BUFx4f_ASAP7_75t_L g851 ( 
.A(n_721),
.Y(n_851)
);

AOI33xp33_ASAP7_75t_L g852 ( 
.A1(n_688),
.A2(n_697),
.A3(n_646),
.B1(n_651),
.B2(n_638),
.B3(n_664),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_SL g853 ( 
.A(n_807),
.B(n_707),
.C(n_699),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_787),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_758),
.B(n_649),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_765),
.B(n_656),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_761),
.A2(n_711),
.B(n_716),
.C(n_735),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_749),
.A2(n_750),
.B(n_747),
.Y(n_858)
);

AO31x2_ASAP7_75t_L g859 ( 
.A1(n_823),
.A2(n_723),
.A3(n_743),
.B(n_716),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_771),
.A2(n_730),
.B(n_696),
.C(n_694),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_772),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_746),
.A2(n_741),
.B1(n_735),
.B2(n_734),
.C(n_694),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_759),
.B(n_687),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_744),
.B(n_720),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_818),
.B(n_736),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_793),
.B(n_755),
.Y(n_866)
);

AO31x2_ASAP7_75t_L g867 ( 
.A1(n_850),
.A2(n_788),
.A3(n_821),
.B(n_831),
.Y(n_867)
);

OAI21x1_ASAP7_75t_SL g868 ( 
.A1(n_829),
.A2(n_848),
.B(n_832),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_745),
.Y(n_869)
);

AO31x2_ASAP7_75t_L g870 ( 
.A1(n_816),
.A2(n_820),
.A3(n_817),
.B(n_753),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_845),
.B(n_752),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_800),
.B(n_822),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_774),
.B(n_776),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_778),
.B(n_776),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_775),
.A2(n_797),
.B1(n_828),
.B2(n_745),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_757),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_774),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_774),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_773),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_840),
.B(n_797),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_798),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_847),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_786),
.B(n_828),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_751),
.B(n_785),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_794),
.B(n_826),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_798),
.B(n_801),
.Y(n_886)
);

BUFx4_ASAP7_75t_SL g887 ( 
.A(n_808),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_766),
.A2(n_769),
.B(n_767),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_798),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_764),
.B(n_779),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_825),
.A2(n_754),
.B(n_762),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_780),
.B(n_770),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_760),
.A2(n_789),
.B(n_814),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_764),
.B(n_851),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_756),
.A2(n_844),
.B(n_790),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_836),
.A2(n_846),
.B(n_781),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_784),
.A2(n_811),
.B(n_809),
.Y(n_897)
);

AND3x4_ASAP7_75t_L g898 ( 
.A(n_830),
.B(n_812),
.C(n_815),
.Y(n_898)
);

NOR4xp25_ASAP7_75t_L g899 ( 
.A(n_804),
.B(n_842),
.C(n_852),
.D(n_837),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_802),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_841),
.A2(n_782),
.B(n_799),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_791),
.A2(n_803),
.B(n_805),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_796),
.A2(n_810),
.B(n_833),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_806),
.A2(n_834),
.B(n_835),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_L g905 ( 
.A(n_768),
.B(n_813),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_795),
.B(n_792),
.Y(n_906)
);

OAI22x1_ASAP7_75t_L g907 ( 
.A1(n_838),
.A2(n_843),
.B1(n_824),
.B2(n_819),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_824),
.B(n_763),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_812),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_777),
.A2(n_742),
.B(n_692),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_744),
.B(n_519),
.Y(n_911)
);

INVx3_ASAP7_75t_SL g912 ( 
.A(n_745),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_747),
.A2(n_742),
.B(n_692),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_758),
.B(n_625),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_744),
.B(n_519),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_772),
.Y(n_916)
);

NOR2x1_ASAP7_75t_SL g917 ( 
.A(n_774),
.B(n_691),
.Y(n_917)
);

AO21x2_ASAP7_75t_L g918 ( 
.A1(n_839),
.A2(n_749),
.B(n_783),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_749),
.A2(n_750),
.B(n_747),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_774),
.B(n_625),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_761),
.A2(n_633),
.B(n_849),
.C(n_634),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_794),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_745),
.Y(n_923)
);

AO21x2_ASAP7_75t_L g924 ( 
.A1(n_839),
.A2(n_749),
.B(n_783),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_761),
.A2(n_587),
.B(n_627),
.C(n_669),
.Y(n_925)
);

OA21x2_ASAP7_75t_L g926 ( 
.A1(n_839),
.A2(n_783),
.B(n_678),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_758),
.B(n_669),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_749),
.A2(n_750),
.B(n_747),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_749),
.A2(n_750),
.B(n_747),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_758),
.B(n_625),
.Y(n_930)
);

AO21x2_ASAP7_75t_L g931 ( 
.A1(n_839),
.A2(n_749),
.B(n_783),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_756),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_SL g933 ( 
.A1(n_748),
.A2(n_640),
.B(n_556),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_758),
.B(n_625),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_771),
.B(n_627),
.C(n_640),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_839),
.A2(n_749),
.B(n_783),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_772),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_758),
.B(n_625),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_745),
.Y(n_939)
);

AO31x2_ASAP7_75t_L g940 ( 
.A1(n_823),
.A2(n_827),
.A3(n_850),
.B(n_788),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_827),
.A2(n_640),
.B1(n_746),
.B2(n_748),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_749),
.A2(n_750),
.B(n_747),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_758),
.B(n_625),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_747),
.A2(n_742),
.B(n_692),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_758),
.B(n_625),
.Y(n_945)
);

INVx8_ASAP7_75t_L g946 ( 
.A(n_745),
.Y(n_946)
);

NOR4xp25_ASAP7_75t_L g947 ( 
.A(n_761),
.B(n_732),
.C(n_822),
.D(n_800),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_747),
.A2(n_750),
.B(n_749),
.Y(n_948)
);

OA21x2_ASAP7_75t_L g949 ( 
.A1(n_839),
.A2(n_783),
.B(n_678),
.Y(n_949)
);

OA21x2_ASAP7_75t_L g950 ( 
.A1(n_839),
.A2(n_783),
.B(n_678),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_772),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_774),
.B(n_636),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_758),
.B(n_625),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_758),
.B(n_669),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_747),
.A2(n_750),
.B(n_749),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_748),
.A2(n_827),
.B1(n_641),
.B2(n_829),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_757),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_749),
.A2(n_750),
.B(n_747),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_745),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_758),
.B(n_669),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_861),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_920),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_901),
.A2(n_910),
.B(n_858),
.Y(n_963)
);

BUFx2_ASAP7_75t_R g964 ( 
.A(n_922),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_921),
.B(n_941),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_911),
.B(n_915),
.Y(n_966)
);

NAND2x1p5_ASAP7_75t_L g967 ( 
.A(n_939),
.B(n_881),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_927),
.B(n_960),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_941),
.A2(n_872),
.B1(n_933),
.B2(n_956),
.Y(n_969)
);

OAI21x1_ASAP7_75t_SL g970 ( 
.A1(n_868),
.A2(n_917),
.B(n_883),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_935),
.B(n_933),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_871),
.B(n_925),
.C(n_864),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_912),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_914),
.B(n_930),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_934),
.B(n_938),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_943),
.B(n_945),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_946),
.Y(n_977)
);

AO31x2_ASAP7_75t_L g978 ( 
.A1(n_907),
.A2(n_891),
.A3(n_895),
.B(n_893),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_916),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_953),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_888),
.A2(n_904),
.B(n_948),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_937),
.Y(n_982)
);

AO31x2_ASAP7_75t_L g983 ( 
.A1(n_879),
.A2(n_896),
.A3(n_884),
.B(n_892),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_946),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_954),
.B(n_866),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_939),
.B(n_886),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_951),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_919),
.A2(n_958),
.B(n_929),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_947),
.B(n_904),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_946),
.Y(n_990)
);

BUFx4f_ASAP7_75t_SL g991 ( 
.A(n_959),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_882),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_955),
.A2(n_928),
.B(n_929),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_902),
.A2(n_942),
.B(n_928),
.Y(n_994)
);

NOR2x1_ASAP7_75t_SL g995 ( 
.A(n_939),
.B(n_890),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_854),
.B(n_923),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_926),
.A2(n_950),
.B(n_949),
.Y(n_997)
);

INVx6_ASAP7_75t_L g998 ( 
.A(n_909),
.Y(n_998)
);

AO21x2_ASAP7_75t_L g999 ( 
.A1(n_918),
.A2(n_936),
.B(n_924),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_880),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_865),
.Y(n_1001)
);

NOR2x1_ASAP7_75t_SL g1002 ( 
.A(n_890),
.B(n_894),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_900),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_931),
.A2(n_936),
.B(n_903),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_875),
.B(n_869),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_947),
.B(n_906),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_952),
.B(n_855),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_899),
.B(n_957),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_913),
.A2(n_944),
.A3(n_897),
.B(n_940),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_898),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_940),
.B(n_856),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_881),
.B(n_889),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_853),
.B(n_874),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_931),
.A2(n_899),
.B(n_932),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_877),
.Y(n_1015)
);

CKINVDCx11_ASAP7_75t_R g1016 ( 
.A(n_909),
.Y(n_1016)
);

AOI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_885),
.A2(n_863),
.B1(n_908),
.B2(n_862),
.C(n_860),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_873),
.B(n_878),
.Y(n_1018)
);

AO31x2_ASAP7_75t_L g1019 ( 
.A1(n_867),
.A2(n_859),
.A3(n_870),
.B(n_905),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_SL g1020 ( 
.A(n_890),
.B(n_957),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_886),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_887),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_876),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_859),
.B(n_876),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_921),
.B(n_941),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_868),
.A2(n_742),
.B(n_857),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_960),
.B(n_927),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_911),
.B(n_915),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_935),
.A2(n_454),
.B1(n_445),
.B2(n_669),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_921),
.B(n_941),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_861),
.Y(n_1031)
);

AO222x2_ASAP7_75t_L g1032 ( 
.A1(n_927),
.A2(n_744),
.B1(n_552),
.B2(n_640),
.C1(n_650),
.C2(n_644),
.Y(n_1032)
);

BUFx8_ASAP7_75t_L g1033 ( 
.A(n_923),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_970),
.B(n_969),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_965),
.B(n_1025),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_980),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_986),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_986),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_971),
.B(n_974),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1011),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_980),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_971),
.B(n_976),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_972),
.A2(n_1006),
.B(n_1010),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_994),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_997),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_983),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_1032),
.B(n_1010),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_1012),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_967),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_969),
.B(n_1026),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_975),
.A2(n_1017),
.B1(n_1030),
.B2(n_1013),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1001),
.B(n_968),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1027),
.B(n_1003),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_967),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_961),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_966),
.B(n_1028),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_981),
.A2(n_993),
.B(n_1014),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_998),
.Y(n_1058)
);

AO21x2_ASAP7_75t_L g1059 ( 
.A1(n_1004),
.A2(n_1008),
.B(n_989),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_989),
.B(n_988),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_987),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_1024),
.A2(n_1013),
.A3(n_1020),
.B(n_1023),
.Y(n_1062)
);

CKINVDCx6p67_ASAP7_75t_R g1063 ( 
.A(n_973),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_985),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_988),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1040),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1040),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1046),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_1042),
.B(n_1019),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1057),
.B(n_963),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_SL g1071 ( 
.A(n_1047),
.B(n_962),
.C(n_1017),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_1062),
.Y(n_1072)
);

INVx4_ASAP7_75t_R g1073 ( 
.A(n_1054),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1034),
.B(n_1044),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1050),
.B(n_999),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1042),
.B(n_999),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_1034),
.B(n_978),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1045),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_L g1079 ( 
.A(n_1054),
.B(n_1021),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1035),
.B(n_1009),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_1054),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1068),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1068),
.Y(n_1083)
);

NAND2x1_ASAP7_75t_L g1084 ( 
.A(n_1073),
.B(n_1034),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1066),
.B(n_1039),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1078),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1066),
.B(n_1039),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_1076),
.B(n_1060),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1081),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1076),
.B(n_1060),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1074),
.B(n_1065),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1081),
.B(n_1049),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1080),
.B(n_1059),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1081),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_1073),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1071),
.B(n_1032),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1067),
.B(n_1048),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1076),
.B(n_1059),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1080),
.B(n_1059),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1094),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1082),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1082),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1086),
.Y(n_1103)
);

NOR2xp67_ASAP7_75t_L g1104 ( 
.A(n_1095),
.B(n_1036),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1093),
.B(n_1080),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1088),
.B(n_1069),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1083),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_1094),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1091),
.B(n_1077),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1085),
.B(n_1087),
.Y(n_1110)
);

AND2x2_ASAP7_75t_SL g1111 ( 
.A(n_1091),
.B(n_1072),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1095),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1101),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1109),
.B(n_1091),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_1105),
.A2(n_1096),
.B(n_1093),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1105),
.B(n_1099),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1103),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1106),
.B(n_1098),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1110),
.B(n_1099),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_1104),
.B(n_1063),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1103),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1106),
.B(n_1098),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1109),
.B(n_1075),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1101),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1109),
.B(n_1075),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1109),
.B(n_1075),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1116),
.B(n_1100),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1120),
.A2(n_1092),
.B(n_1108),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1115),
.A2(n_1111),
.B(n_1084),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1116),
.B(n_1102),
.Y(n_1130)
);

OAI32xp33_ASAP7_75t_L g1131 ( 
.A1(n_1118),
.A2(n_1089),
.A3(n_1041),
.B1(n_1111),
.B2(n_1037),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1113),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_1117),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1113),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1114),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1124),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1118),
.B(n_1088),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1123),
.A2(n_1111),
.B1(n_1071),
.B2(n_1091),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1123),
.B(n_1070),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1131),
.A2(n_1119),
.B1(n_1043),
.B2(n_1125),
.C(n_1126),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1129),
.A2(n_1084),
.B(n_1112),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1139),
.B(n_1122),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1132),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_SL g1144 ( 
.A(n_1128),
.B(n_1112),
.C(n_1122),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_1135),
.A2(n_1064),
.B(n_1038),
.C(n_1063),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1138),
.A2(n_1022),
.B(n_1005),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1135),
.A2(n_1114),
.B1(n_1126),
.B2(n_1125),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1143),
.Y(n_1148)
);

NOR4xp25_ASAP7_75t_L g1149 ( 
.A(n_1144),
.B(n_1140),
.C(n_1146),
.D(n_1147),
.Y(n_1149)
);

AOI211xp5_ASAP7_75t_L g1150 ( 
.A1(n_1145),
.A2(n_1043),
.B(n_1137),
.C(n_1114),
.Y(n_1150)
);

AOI211x1_ASAP7_75t_L g1151 ( 
.A1(n_1141),
.A2(n_1127),
.B(n_1130),
.C(n_1139),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1142),
.A2(n_1133),
.B1(n_1134),
.B2(n_1136),
.C(n_1124),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1140),
.B(n_1133),
.C(n_1079),
.Y(n_1153)
);

AND4x1_ASAP7_75t_L g1154 ( 
.A(n_1141),
.B(n_1029),
.C(n_964),
.D(n_1051),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1142),
.B(n_1090),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_1151),
.B(n_1033),
.C(n_1000),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_1149),
.B(n_1033),
.C(n_1079),
.Y(n_1157)
);

NOR4xp25_ASAP7_75t_L g1158 ( 
.A(n_1153),
.B(n_1015),
.C(n_1056),
.D(n_1055),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1148),
.Y(n_1159)
);

AOI221xp5_ASAP7_75t_L g1160 ( 
.A1(n_1150),
.A2(n_1114),
.B1(n_1097),
.B2(n_1107),
.C(n_1102),
.Y(n_1160)
);

AOI211xp5_ASAP7_75t_L g1161 ( 
.A1(n_1152),
.A2(n_990),
.B(n_1051),
.C(n_1053),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_964),
.Y(n_1162)
);

NAND4xp75_ASAP7_75t_L g1163 ( 
.A(n_1162),
.B(n_977),
.C(n_984),
.D(n_1007),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1157),
.B(n_1156),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_SL g1165 ( 
.A(n_1158),
.B(n_1161),
.C(n_1160),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1159),
.B(n_1155),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1161),
.B(n_1117),
.Y(n_1167)
);

AND4x1_ASAP7_75t_L g1168 ( 
.A(n_1157),
.B(n_991),
.C(n_1018),
.D(n_1016),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1157),
.B(n_1016),
.C(n_992),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1164),
.B(n_991),
.Y(n_1170)
);

NAND3x1_ASAP7_75t_SL g1171 ( 
.A(n_1168),
.B(n_1163),
.C(n_1165),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1169),
.B(n_1121),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_1166),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_R g1174 ( 
.A(n_1167),
.B(n_996),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1165),
.A2(n_1058),
.B(n_979),
.C(n_982),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1170),
.B(n_1053),
.Y(n_1176)
);

OAI211xp5_ASAP7_75t_L g1177 ( 
.A1(n_1175),
.A2(n_1058),
.B(n_1018),
.C(n_1038),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1176),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1177),
.A2(n_1173),
.B1(n_1171),
.B2(n_1174),
.Y(n_1179)
);

INVxp67_ASAP7_75t_SL g1180 ( 
.A(n_1179),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1178),
.A2(n_1172),
.B(n_1058),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1180),
.B(n_1052),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1182),
.A2(n_1181),
.B(n_995),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1182),
.A2(n_1002),
.B(n_1031),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1183),
.B(n_1055),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1185),
.A2(n_1184),
.B(n_1061),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1186),
.A2(n_1052),
.B(n_998),
.Y(n_1187)
);


endmodule