module real_jpeg_15508_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_560),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_0),
.B(n_561),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_1),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_1),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_1),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_1),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_1),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_1),
.A2(n_3),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_1),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_2),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_3),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_3),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_3),
.B(n_370),
.Y(n_369)
);

AOI31xp33_ASAP7_75t_SL g402 ( 
.A1(n_3),
.A2(n_301),
.A3(n_403),
.B(n_405),
.Y(n_402)
);

NAND2x1_ASAP7_75t_SL g444 ( 
.A(n_3),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_3),
.B(n_108),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_3),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_3),
.B(n_517),
.Y(n_516)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_4),
.Y(n_423)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_5),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_5),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_6),
.Y(n_181)
);

NAND2x1_ASAP7_75t_SL g183 ( 
.A(n_6),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_6),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g320 ( 
.A(n_6),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_6),
.B(n_108),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_6),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_6),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_7),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_7),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_7),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_7),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_7),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g367 ( 
.A(n_7),
.B(n_258),
.Y(n_367)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_8),
.Y(n_226)
);

BUFx4f_ASAP7_75t_L g412 ( 
.A(n_8),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_8),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_9),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_9),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_9),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_9),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_9),
.B(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_9),
.B(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_9),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_10),
.B(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_11),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_12),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_12),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_13),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_13),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_13),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_13),
.B(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_14),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_14),
.Y(n_146)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_14),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_15),
.B(n_67),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_15),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_15),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_15),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_15),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_15),
.B(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_15),
.B(n_325),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_16),
.B(n_93),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_16),
.B(n_84),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_16),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_16),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_16),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_16),
.B(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g184 ( 
.A(n_18),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_117),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_116),
.Y(n_21)
);

NAND2x1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_72),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_72),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_54),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.C(n_35),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_32),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_30),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_31),
.Y(n_163)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_31),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_64),
.C(n_69),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_32),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_45),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_107),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_46),
.B(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_63),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_55),
.A2(n_56),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_62),
.Y(n_222)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_62),
.Y(n_323)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

XOR2x1_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_69),
.A2(n_70),
.B1(n_106),
.B2(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_103),
.C(n_106),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_111),
.C(n_112),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_102),
.C(n_109),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_74),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_91),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_92),
.C(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_82),
.C(n_87),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_173)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_79),
.Y(n_336)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_80),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_81),
.Y(n_306)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_87),
.B(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_102),
.B(n_109),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_103),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_106),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_158),
.C(n_166),
.Y(n_190)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_291),
.B(n_555),
.Y(n_118)
);

NOR3x1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_195),
.C(n_285),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_120),
.A2(n_556),
.B(n_559),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_121),
.B(n_123),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_187),
.C(n_192),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_124),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_172),
.C(n_174),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_126),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_140),
.C(n_157),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_127),
.B(n_140),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_130),
.C(n_135),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_139),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.C(n_152),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_141),
.B(n_152),
.Y(n_218)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_145),
.Y(n_446)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_147),
.B(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_151),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_156),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_162),
.Y(n_269)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_166),
.A2(n_167),
.B1(n_177),
.B2(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_177),
.C(n_180),
.Y(n_176)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_172),
.B(n_174),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_183),
.C(n_185),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_176),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_220),
.C(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_177),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_177),
.A2(n_223),
.B1(n_231),
.B2(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_179),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_180),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_180),
.A2(n_228),
.B1(n_313),
.B2(n_362),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_185),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_183),
.B(n_257),
.C(n_261),
.Y(n_256)
);

XNOR2x2_ASAP7_75t_SL g298 ( 
.A(n_183),
.B(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_185),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_185),
.A2(n_214),
.B1(n_215),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_187),
.A2(n_192),
.B1(n_193),
.B2(n_289),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_187),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_190),
.B(n_191),
.Y(n_280)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_274),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_196),
.B(n_274),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_232),
.C(n_235),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_197),
.B(n_232),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_216),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_202),
.B(n_276),
.C(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_214),
.C(n_215),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_203),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_213),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_213),
.Y(n_254)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_208),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_227),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_217),
.B(n_219),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_226),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_308),
.C(n_313),
.Y(n_307)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_235),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_255),
.C(n_270),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_236),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.C(n_253),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_237),
.B(n_240),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.C(n_248),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_241),
.A2(n_248),
.B1(n_249),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_241),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_245),
.B(n_381),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_248),
.B(n_440),
.C(n_444),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_248),
.A2(n_249),
.B1(n_440),
.B2(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g354 ( 
.A(n_253),
.B(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_255),
.B(n_271),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_264),
.C(n_267),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_256),
.B(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_261),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_260),
.Y(n_416)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_264),
.B(n_268),
.Y(n_339)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_265),
.Y(n_523)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_267),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_267),
.A2(n_268),
.B1(n_418),
.B2(n_419),
.Y(n_539)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_279),
.C(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_286),
.A2(n_557),
.B(n_558),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_287),
.B(n_290),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_389),
.B(n_552),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_383),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_348),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_294),
.B(n_348),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_340),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_295),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_317),
.C(n_337),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_307),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_298),
.B(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_300),
.A2(n_301),
.B1(n_307),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_303),
.B(n_406),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_307),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_312),
.Y(n_464)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_318),
.A2(n_337),
.B1(n_338),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_328),
.C(n_335),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.C(n_324),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_320),
.B(n_324),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_320),
.B(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_320),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_322),
.B(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_329),
.B1(n_335),
.B2(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_343),
.B1(n_346),
.B2(n_347),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_341),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_346),
.B(n_387),
.C(n_388),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.C(n_356),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_350),
.A2(n_351),
.B1(n_354),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_377),
.C(n_380),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_358),
.B(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.C(n_368),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_SL g449 ( 
.A(n_360),
.B(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_363),
.B(n_368),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_364),
.B(n_367),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_366),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_373),
.C(n_374),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_369),
.A2(n_373),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_373),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_373),
.B(n_504),
.C(n_506),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_373),
.A2(n_437),
.B1(n_506),
.B2(n_507),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_374),
.B(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_376),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_380),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_383),
.A2(n_553),
.B(n_554),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_384),
.B(n_386),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_451),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.C(n_427),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.C(n_424),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_424),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.C(n_407),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_402),
.Y(n_432)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_432),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_417),
.C(n_418),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_408),
.B(n_539),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_413),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_409),
.B(n_413),
.Y(n_490)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_409),
.A2(n_515),
.B1(n_516),
.B2(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_430),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.C(n_449),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_431),
.B(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_433),
.B(n_449),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_438),
.C(n_447),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_434),
.B(n_544),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_439),
.B(n_448),
.Y(n_544)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

INVx8_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XOR2x2_ASAP7_75t_L g495 ( 
.A(n_444),
.B(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND3xp33_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_453),
.C(n_454),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_455),
.A2(n_547),
.B(n_551),
.Y(n_454)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_533),
.B(n_546),
.Y(n_455)
);

OAI21x1_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_498),
.B(n_532),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_486),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_458),
.B(n_486),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_466),
.C(n_475),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_459),
.B(n_501),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_465),
.C(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_467),
.B1(n_475),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_472),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_468),
.B(n_472),
.Y(n_505)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

AO22x1_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_481),
.B1(n_484),
.B2(n_485),
.Y(n_475)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_476),
.Y(n_484)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_481),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_484),
.Y(n_488)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_482),
.Y(n_518)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_527),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_492),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_487),
.B(n_493),
.C(n_495),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

MAJx2_ASAP7_75t_L g541 ( 
.A(n_488),
.B(n_490),
.C(n_491),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_495),
.Y(n_492)
);

AOI21x1_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_509),
.B(n_531),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_503),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g531 ( 
.A(n_500),
.B(n_503),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_504),
.A2(n_505),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_510),
.A2(n_519),
.B(n_530),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_514),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_514),
.Y(n_530)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_516),
.Y(n_525)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_526),
.B(n_529),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_524),
.Y(n_529)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_534),
.B(n_545),
.Y(n_533)
);

NOR2x1p5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_545),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_535),
.A2(n_536),
.B1(n_542),
.B2(n_543),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_538),
.B1(n_540),
.B2(n_541),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_541),
.C(n_542),
.Y(n_548)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_SL g547 ( 
.A(n_548),
.B(n_549),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_549),
.Y(n_551)
);


endmodule