module real_jpeg_28075_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_106)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_20),
.B1(n_45),
.B2(n_46),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_20),
.B1(n_38),
.B2(n_39),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_5),
.A2(n_26),
.B(n_30),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_6),
.B(n_39),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_5),
.B(n_59),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_5),
.A2(n_8),
.B(n_29),
.C(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_87)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_92),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_91),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_80),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.C(n_67),
.Y(n_15)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_16),
.B(n_62),
.CI(n_67),
.CON(n_112),
.SN(n_112)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_31),
.B2(n_32),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_17),
.A2(n_18),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_17),
.A2(n_18),
.B1(n_70),
.B2(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_17),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_17),
.B(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_17),
.A2(n_18),
.B1(n_65),
.B2(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_17),
.A2(n_18),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_18),
.A2(n_68),
.B(n_79),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_18),
.B(n_33),
.C(n_50),
.Y(n_90)
);

AOI211xp5_ASAP7_75t_L g120 ( 
.A1(n_18),
.A2(n_109),
.B(n_111),
.C(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_20),
.A2(n_21),
.B(n_27),
.C(n_135),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_20),
.A2(n_41),
.B(n_46),
.C(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_20),
.B(n_37),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_20),
.B(n_171),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_20),
.A2(n_45),
.B(n_57),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_26),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_28),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_29),
.A2(n_30),
.B1(n_55),
.B2(n_57),
.Y(n_58)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_33),
.A2(n_34),
.B1(n_85),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_47),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_36),
.B(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_42),
.B1(n_47),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_37),
.A2(n_42),
.B1(n_64),
.B2(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_38),
.B(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_73),
.Y(n_74)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_46),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_54),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_63),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_65),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_103),
.B1(n_109),
.B2(n_122),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_136),
.C(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_65),
.A2(n_103),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_69),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_70),
.A2(n_76),
.B1(n_79),
.B2(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_73),
.A2(n_74),
.B1(n_106),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_75),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_76),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_113),
.B(n_235),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_112),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_94),
.B(n_112),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.C(n_99),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_95),
.B(n_98),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_99),
.A2(n_100),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B(n_110),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_101),
.A2(n_110),
.B(n_211),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_102),
.A2(n_111),
.B(n_138),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_122),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_103),
.A2(n_122),
.B(n_183),
.C(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_104),
.A2(n_130),
.B1(n_131),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_104),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_105),
.A2(n_109),
.B1(n_122),
.B2(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_105),
.Y(n_214)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_122),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_109),
.A2(n_122),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_122),
.B1(n_157),
.B2(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_136),
.C(n_161),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_109),
.A2(n_122),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_189),
.C(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_109),
.B(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_112),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_229),
.B(n_234),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_219),
.B(n_228),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_150),
.B(n_206),
.C(n_218),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_139),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_139),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_129),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_119),
.B(n_124),
.C(n_129),
.Y(n_207)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_138),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_130),
.A2(n_131),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_137),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_137),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_136),
.A2(n_137),
.B1(n_147),
.B2(n_148),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_146),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_141),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_143),
.B1(n_179),
.B2(n_183),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_205),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_198),
.B(n_204),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_185),
.B(n_197),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_176),
.B(n_184),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_164),
.B(n_175),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_172),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_208),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_217),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_215),
.C(n_217),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_225),
.C(n_227),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);


endmodule