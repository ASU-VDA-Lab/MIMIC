module fake_jpeg_2293_n_553 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_553);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_3),
.B(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_64),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_9),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_73),
.B(n_99),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_75),
.Y(n_192)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_52),
.Y(n_123)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_88),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_26),
.B(n_10),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_39),
.B(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_117),
.Y(n_136)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_43),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_103),
.B(n_35),
.Y(n_182)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_46),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_48),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_116),
.Y(n_164)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g173 ( 
.A(n_118),
.Y(n_173)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_121),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_122),
.B(n_17),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_17),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_123),
.B(n_129),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_37),
.B1(n_32),
.B2(n_58),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_124),
.A2(n_134),
.B1(n_147),
.B2(n_155),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_31),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_133),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_37),
.B1(n_32),
.B2(n_58),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_57),
.C(n_56),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_140),
.B(n_196),
.C(n_178),
.Y(n_266)
);

NAND2x1_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_56),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_142),
.B(n_17),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_37),
.B1(n_54),
.B2(n_53),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_54),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_148),
.B(n_176),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_59),
.A2(n_23),
.B1(n_52),
.B2(n_47),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_153),
.A2(n_7),
.B1(n_15),
.B2(n_4),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_95),
.A2(n_57),
.B1(n_53),
.B2(n_31),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_156),
.A2(n_196),
.B(n_186),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_95),
.A2(n_19),
.B1(n_27),
.B2(n_20),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_158),
.A2(n_183),
.B1(n_197),
.B2(n_198),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_47),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_82),
.B(n_45),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_86),
.B(n_45),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_177),
.B(n_182),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_23),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_91),
.A2(n_48),
.B1(n_19),
.B2(n_20),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_110),
.B(n_35),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_199),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_93),
.A2(n_27),
.B1(n_17),
.B2(n_0),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_60),
.A2(n_17),
.B1(n_38),
.B2(n_36),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_96),
.B(n_12),
.Y(n_199)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_206),
.Y(n_298)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_208),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_136),
.A2(n_69),
.B1(n_63),
.B2(n_65),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_209),
.B(n_212),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_210),
.B(n_216),
.Y(n_282)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_213),
.Y(n_273)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_214),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_133),
.Y(n_216)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx11_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_75),
.B1(n_66),
.B2(n_74),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_221),
.A2(n_249),
.B1(n_250),
.B2(n_257),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_124),
.Y(n_222)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_164),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_226),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_237),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_162),
.B(n_0),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_228),
.B(n_236),
.Y(n_302)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_230),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_131),
.B(n_98),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_231),
.B(n_234),
.Y(n_300)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_142),
.B(n_125),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_143),
.Y(n_235)
);

BUFx4f_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_127),
.B(n_87),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_240),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_61),
.B1(n_97),
.B2(n_118),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_255),
.B1(n_261),
.B2(n_268),
.Y(n_275)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_242),
.B(n_243),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_125),
.A2(n_44),
.B1(n_38),
.B2(n_118),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_244),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_269)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_245),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_191),
.Y(n_246)
);

BUFx8_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_162),
.B(n_44),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_248),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_138),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_146),
.A2(n_11),
.B1(n_15),
.B2(n_6),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_149),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_251),
.Y(n_316)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_141),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_134),
.A2(n_6),
.B(n_7),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_264),
.B(n_169),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_183),
.A2(n_0),
.B1(n_2),
.B2(n_7),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_138),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_147),
.A2(n_11),
.B1(n_13),
.B2(n_2),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_263),
.B1(n_267),
.B2(n_160),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_151),
.B(n_187),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_262),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_155),
.A2(n_2),
.B1(n_11),
.B2(n_158),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_190),
.B(n_179),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_167),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_192),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_247),
.Y(n_310)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_137),
.A2(n_161),
.B1(n_195),
.B2(n_152),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_271),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_222),
.A2(n_160),
.B1(n_126),
.B2(n_150),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_279),
.A2(n_306),
.B1(n_309),
.B2(n_318),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_169),
.C(n_184),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_310),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_283),
.A2(n_308),
.B(n_273),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_287),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_239),
.A2(n_216),
.B1(n_212),
.B2(n_225),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_307),
.B1(n_209),
.B2(n_254),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_161),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_137),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_210),
.B(n_150),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_317),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_223),
.A2(n_152),
.B1(n_172),
.B2(n_174),
.Y(n_297)
);

AO21x2_ASAP7_75t_L g355 ( 
.A1(n_297),
.A2(n_314),
.B(n_301),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_226),
.A2(n_126),
.B1(n_172),
.B2(n_174),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_249),
.A2(n_184),
.B1(n_192),
.B2(n_217),
.Y(n_307)
);

AOI22x1_ASAP7_75t_SL g308 ( 
.A1(n_217),
.A2(n_261),
.B1(n_209),
.B2(n_262),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_201),
.A2(n_268),
.B1(n_204),
.B2(n_208),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_205),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_265),
.A2(n_242),
.B1(n_235),
.B2(n_237),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_215),
.B(n_219),
.C(n_207),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_230),
.C(n_233),
.Y(n_327)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_322),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_348),
.Y(n_382)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_292),
.A2(n_236),
.B1(n_255),
.B2(n_229),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_326),
.A2(n_328),
.B1(n_331),
.B2(n_343),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_236),
.B1(n_232),
.B2(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_317),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_330),
.B(n_359),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_292),
.A2(n_206),
.B1(n_211),
.B2(n_251),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_275),
.A2(n_220),
.B1(n_252),
.B2(n_203),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_333),
.A2(n_341),
.B1(n_342),
.B2(n_347),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_213),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_202),
.B(n_246),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_338),
.A2(n_351),
.B(n_357),
.Y(n_389)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_275),
.A2(n_253),
.B1(n_267),
.B2(n_227),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_243),
.B1(n_214),
.B2(n_258),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_218),
.B1(n_281),
.B2(n_293),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_344),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_281),
.A2(n_296),
.B1(n_291),
.B2(n_295),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_345),
.A2(n_349),
.B1(n_355),
.B2(n_361),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_294),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_350),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_285),
.A2(n_310),
.B1(n_302),
.B2(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_295),
.A2(n_302),
.B1(n_270),
.B2(n_269),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_280),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_353),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_273),
.B(n_300),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_312),
.A2(n_311),
.B(n_290),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_321),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_299),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_304),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_360),
.B(n_315),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_305),
.A2(n_304),
.B1(n_314),
.B2(n_316),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_276),
.C(n_316),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_368),
.C(n_274),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_347),
.A2(n_305),
.B1(n_313),
.B2(n_299),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_371),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_276),
.C(n_278),
.Y(n_368)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

O2A1O1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_343),
.A2(n_288),
.B(n_294),
.C(n_286),
.Y(n_375)
);

OAI31xp33_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_387),
.A3(n_334),
.B(n_288),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_358),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_376),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_278),
.Y(n_377)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_345),
.B(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_379),
.B(n_388),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_335),
.B(n_298),
.Y(n_384)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_315),
.Y(n_385)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_351),
.A2(n_288),
.B(n_286),
.C(n_274),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_361),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_353),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_390),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_346),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_392),
.A2(n_322),
.B(n_337),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_340),
.B(n_320),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_393),
.B(n_339),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_370),
.B(n_357),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_370),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_382),
.A2(n_323),
.B1(n_352),
.B2(n_333),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_401),
.B1(n_413),
.B2(n_411),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_382),
.A2(n_355),
.B1(n_341),
.B2(n_338),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_381),
.Y(n_402)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_402),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_403),
.A2(n_373),
.B(n_387),
.Y(n_438)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_407),
.A2(n_410),
.B1(n_380),
.B2(n_394),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_389),
.A2(n_334),
.B(n_332),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_408),
.A2(n_418),
.B(n_424),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_327),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_364),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_380),
.A2(n_349),
.B1(n_326),
.B2(n_328),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_342),
.B(n_331),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_416),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_412),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_382),
.A2(n_355),
.B1(n_339),
.B2(n_356),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_414),
.Y(n_436)
);

OAI32xp33_ASAP7_75t_L g416 ( 
.A1(n_369),
.A2(n_324),
.A3(n_329),
.B1(n_348),
.B2(n_360),
.Y(n_416)
);

A2O1A1O1Ixp25_ASAP7_75t_L g418 ( 
.A1(n_390),
.A2(n_350),
.B(n_355),
.C(n_344),
.D(n_336),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_420),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_425),
.C(n_368),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_389),
.A2(n_320),
.B(n_355),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_368),
.B(n_284),
.C(n_365),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_426),
.A2(n_428),
.B1(n_429),
.B2(n_441),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_400),
.A2(n_413),
.B1(n_424),
.B2(n_401),
.Y(n_428)
);

AOI22x1_ASAP7_75t_L g429 ( 
.A1(n_415),
.A2(n_367),
.B1(n_363),
.B2(n_387),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_430),
.B(n_372),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_381),
.C(n_386),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_392),
.Y(n_432)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_432),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_419),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_438),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_365),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_452),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_377),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_408),
.A2(n_376),
.B(n_395),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_407),
.Y(n_455)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_399),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_451),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_394),
.B1(n_388),
.B2(n_363),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_446),
.A2(n_447),
.B1(n_396),
.B2(n_417),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_421),
.A2(n_394),
.B1(n_366),
.B2(n_395),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_397),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_409),
.B(n_384),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_432),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_460),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_449),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_457),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_425),
.Y(n_459)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_462),
.C(n_467),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_414),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_465),
.C(n_466),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_417),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_474),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_404),
.C(n_397),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_404),
.C(n_385),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_443),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_410),
.C(n_422),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_471),
.C(n_391),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_470),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_422),
.C(n_393),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_379),
.Y(n_473)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_366),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_461),
.Y(n_476)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_494),
.Y(n_495)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_478),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_444),
.B(n_427),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_479),
.A2(n_483),
.B(n_466),
.Y(n_506)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_482),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_472),
.A2(n_444),
.B(n_438),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_464),
.B(n_427),
.Y(n_484)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_489),
.C(n_490),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_469),
.A2(n_429),
.B1(n_366),
.B2(n_411),
.Y(n_485)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_485),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_486),
.B(n_465),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_458),
.B(n_418),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_391),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_463),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_468),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_496),
.B(n_506),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_501),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_454),
.Y(n_500)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_500),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_483),
.A2(n_474),
.B1(n_471),
.B2(n_467),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_480),
.C(n_492),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_505),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_493),
.C(n_487),
.Y(n_505)
);

MAJx2_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_458),
.C(n_462),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_482),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_479),
.A2(n_375),
.B(n_439),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_486),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_488),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_511),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_487),
.C(n_491),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_434),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_514),
.B(n_515),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_489),
.C(n_484),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_495),
.A2(n_478),
.B(n_434),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_516),
.A2(n_519),
.B(n_512),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_518),
.B(n_506),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_507),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_439),
.C(n_450),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_509),
.C(n_502),
.Y(n_524)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_526),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_520),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_496),
.C(n_508),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_527),
.B(n_528),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_500),
.B1(n_499),
.B2(n_501),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_530),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_412),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_531),
.B(n_525),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_535),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_522),
.A2(n_517),
.B(n_515),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_533),
.A2(n_539),
.B(n_504),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_527),
.B(n_517),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_530),
.A2(n_504),
.B(n_362),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_537),
.B(n_523),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_541),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_534),
.B(n_526),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_543),
.B(n_536),
.C(n_420),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_538),
.B(n_450),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_544),
.A2(n_536),
.B(n_374),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_546),
.A2(n_374),
.B(n_383),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_540),
.B1(n_545),
.B2(n_542),
.Y(n_548)
);

AO21x1_ASAP7_75t_L g550 ( 
.A1(n_548),
.A2(n_549),
.B(n_383),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_372),
.C(n_405),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_371),
.C(n_375),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_284),
.Y(n_553)
);


endmodule