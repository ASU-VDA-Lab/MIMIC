module fake_jpeg_9568_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_38),
.B1(n_21),
.B2(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_0),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_21),
.B1(n_17),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_50),
.B1(n_56),
.B2(n_59),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_17),
.B1(n_35),
.B2(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_17),
.B1(n_20),
.B2(n_19),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_28),
.B1(n_24),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_67),
.B1(n_44),
.B2(n_38),
.Y(n_88)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_94),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_47),
.B(n_49),
.C(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_35),
.B(n_31),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_82),
.A3(n_93),
.B1(n_33),
.B2(n_60),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_83),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_33),
.B(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_95),
.B1(n_58),
.B2(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_59),
.B1(n_38),
.B2(n_44),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_37),
.C(n_46),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.C(n_75),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_33),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_32),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_110),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_51),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_115),
.C(n_71),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_48),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_103),
.B(n_112),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_107),
.B1(n_80),
.B2(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_0),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_44),
.B1(n_58),
.B2(n_52),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_114),
.B1(n_90),
.B2(n_70),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_60),
.B1(n_54),
.B2(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_122),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_54),
.B1(n_60),
.B2(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_80),
.B1(n_84),
.B2(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_54),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_97),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_135),
.B(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_121),
.C(n_30),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_137),
.B1(n_140),
.B2(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_124),
.B(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_89),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_144),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_115),
.B1(n_102),
.B2(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_151),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_141),
.B1(n_117),
.B2(n_33),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_72),
.B1(n_76),
.B2(n_79),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_43),
.B1(n_77),
.B2(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_32),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_43),
.B1(n_36),
.B2(n_29),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_150),
.B1(n_155),
.B2(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_32),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_27),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_96),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_87),
.B1(n_36),
.B2(n_53),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_108),
.B(n_29),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_33),
.B(n_30),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_123),
.B(n_116),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_167),
.B1(n_187),
.B2(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_162),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_121),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_171),
.C(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_173),
.B(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_186),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_118),
.B1(n_27),
.B2(n_29),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_11),
.B(n_16),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_22),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_154),
.B1(n_155),
.B2(n_150),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_121),
.B(n_22),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_121),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_30),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_146),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_155),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_142),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_138),
.A2(n_117),
.B1(n_30),
.B2(n_23),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_157),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_137),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_209),
.C(n_4),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_126),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_134),
.B1(n_145),
.B2(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_205),
.B1(n_187),
.B2(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_150),
.B1(n_154),
.B2(n_152),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_150),
.B1(n_147),
.B2(n_133),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_156),
.A2(n_160),
.B1(n_178),
.B2(n_169),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_207),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_150),
.B(n_135),
.C(n_130),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_212),
.B1(n_216),
.B2(n_172),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_128),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_135),
.B(n_144),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_135),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_30),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_162),
.B1(n_163),
.B2(n_176),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_23),
.B1(n_22),
.B2(n_9),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_161),
.B(n_23),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_22),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_180),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_228),
.C(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_208),
.B1(n_204),
.B2(n_202),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_235),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_171),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_174),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_236),
.C(n_237),
.Y(n_252)
);

AOI22x1_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_22),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_243),
.B1(n_206),
.B2(n_207),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_234),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_10),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_4),
.C(n_5),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_242),
.C(n_200),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_11),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_11),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_211),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_5),
.C(n_6),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_243)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_206),
.B(n_194),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_258),
.B(n_231),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_260),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_227),
.B1(n_205),
.B2(n_236),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_214),
.C(n_195),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_263),
.C(n_237),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_195),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_218),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_223),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_205),
.C(n_212),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_13),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_224),
.C(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_279),
.C(n_281),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_248),
.Y(n_286)
);

XOR2x1_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_256),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_258),
.B(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_250),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_235),
.C(n_5),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_7),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_292),
.C(n_295),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_289),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_272),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_255),
.B(n_252),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_253),
.C(n_252),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_262),
.CI(n_12),
.CON(n_293),
.SN(n_293)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_8),
.CI(n_12),
.CON(n_294),
.SN(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_13),
.C(n_15),
.Y(n_295)
);

O2A1O1Ixp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_278),
.B(n_276),
.C(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_268),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_270),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_282),
.A2(n_265),
.B1(n_279),
.B2(n_268),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_13),
.C(n_15),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_291),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_297),
.B(n_290),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_291),
.B(n_287),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_301),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_294),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_300),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_320),
.A2(n_323),
.B(n_311),
.C(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_303),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_322),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_324),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_326),
.B(n_295),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_320),
.B(n_15),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_16),
.B(n_317),
.Y(n_331)
);


endmodule