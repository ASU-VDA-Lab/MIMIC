module fake_jpeg_2868_n_644 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_60),
.Y(n_206)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_63),
.Y(n_162)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_67),
.B(n_81),
.Y(n_138)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g201 ( 
.A(n_75),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_78),
.Y(n_178)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_110),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_37),
.B(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_10),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_12),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_39),
.B(n_12),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_12),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_121),
.Y(n_157)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_57),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_45),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_20),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_18),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_16),
.Y(n_167)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_21),
.Y(n_128)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_81),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_153),
.B(n_183),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_63),
.A2(n_43),
.B1(n_27),
.B2(n_36),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_155),
.A2(n_160),
.B1(n_168),
.B2(n_182),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_36),
.B1(n_47),
.B2(n_29),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_187),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_70),
.A2(n_27),
.B1(n_47),
.B2(n_43),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_170),
.B(n_0),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_116),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_59),
.B(n_32),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_94),
.B(n_40),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_62),
.A2(n_57),
.B1(n_52),
.B2(n_54),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_189),
.A2(n_198),
.B1(n_210),
.B2(n_211),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_54),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_55),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_55),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_199),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_109),
.A2(n_43),
.B1(n_27),
.B2(n_49),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_68),
.B(n_49),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_98),
.Y(n_203)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_124),
.A2(n_45),
.B1(n_41),
.B2(n_40),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_219),
.B1(n_118),
.B2(n_110),
.Y(n_254)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_72),
.A2(n_41),
.B1(n_34),
.B2(n_32),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_123),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_66),
.A2(n_73),
.B1(n_85),
.B2(n_30),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_97),
.B1(n_108),
.B2(n_95),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_126),
.A2(n_31),
.B1(n_28),
.B2(n_34),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_118),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_66),
.B(n_26),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_215),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_73),
.B(n_26),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_85),
.B(n_28),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_220),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_76),
.A2(n_77),
.B1(n_104),
.B2(n_103),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_78),
.B(n_28),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_221),
.B(n_240),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_142),
.B(n_83),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_222),
.B(n_255),
.Y(n_301)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_228),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_229),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_135),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_230),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_231),
.Y(n_326)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_232),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_160),
.A2(n_88),
.B1(n_90),
.B2(n_101),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_233),
.A2(n_250),
.B1(n_292),
.B2(n_297),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_140),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_234),
.B(n_279),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_236),
.A2(n_291),
.B1(n_295),
.B2(n_296),
.Y(n_303)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_238),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_239),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_201),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_241),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_243),
.Y(n_308)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_170),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_245),
.B(n_253),
.Y(n_305)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_247),
.B(n_293),
.Y(n_355)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_149),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_248),
.Y(n_339)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_158),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_254),
.A2(n_180),
.B1(n_179),
.B2(n_144),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_130),
.B(n_6),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_133),
.B(n_6),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_260),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_138),
.A2(n_6),
.B(n_17),
.C(n_15),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_258),
.B(n_276),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_213),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_259),
.A2(n_298),
.B1(n_163),
.B2(n_175),
.Y(n_349)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_139),
.A2(n_18),
.B(n_17),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_261),
.B(n_262),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_156),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_263),
.B(n_268),
.Y(n_336)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_135),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_266),
.Y(n_311)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_151),
.B(n_17),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_269),
.B(n_270),
.Y(n_352)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_271),
.B(n_273),
.Y(n_357)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_206),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_129),
.B(n_13),
.C(n_1),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_137),
.C(n_159),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_132),
.B(n_13),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_200),
.Y(n_277)
);

INVx6_ASAP7_75t_SL g344 ( 
.A(n_277),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_145),
.B(n_0),
.Y(n_279)
);

AO22x1_ASAP7_75t_SL g280 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_156),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_284),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_207),
.B(n_13),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_283),
.B(n_285),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_136),
.B(n_0),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g286 ( 
.A(n_177),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_147),
.B(n_2),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_294),
.Y(n_333)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_186),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_290),
.Y(n_332)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_178),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_200),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_178),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_165),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g297 ( 
.A1(n_211),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_143),
.B(n_3),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_272),
.A2(n_146),
.B1(n_172),
.B2(n_184),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_SL g375 ( 
.A1(n_313),
.A2(n_315),
.B(n_316),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_288),
.A2(n_146),
.B1(n_172),
.B2(n_161),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_284),
.A2(n_150),
.B1(n_152),
.B2(n_173),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_250),
.A2(n_233),
.B1(n_226),
.B2(n_292),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_329),
.B1(n_347),
.B2(n_291),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_350),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_247),
.A2(n_227),
.B1(n_239),
.B2(n_248),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_321),
.A2(n_335),
.B1(n_337),
.B2(n_231),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_278),
.A2(n_164),
.B1(n_162),
.B2(n_202),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_330),
.B1(n_334),
.B2(n_346),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_247),
.A2(n_297),
.B1(n_279),
.B2(n_287),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_280),
.A2(n_164),
.B1(n_162),
.B2(n_202),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_239),
.A2(n_131),
.B1(n_134),
.B2(n_144),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_238),
.A2(n_131),
.B1(n_134),
.B2(n_180),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_280),
.A2(n_179),
.B1(n_192),
.B2(n_196),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_341),
.A2(n_348),
.B1(n_349),
.B2(n_295),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_223),
.A2(n_234),
.B1(n_264),
.B2(n_242),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_258),
.A2(n_192),
.B1(n_196),
.B2(n_165),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_265),
.A2(n_137),
.B1(n_163),
.B2(n_175),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_256),
.B(n_177),
.C(n_4),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_275),
.A2(n_5),
.B1(n_266),
.B2(n_241),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_356),
.A2(n_274),
.B1(n_224),
.B2(n_230),
.Y(n_373)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_344),
.Y(n_359)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_318),
.A2(n_249),
.B1(n_246),
.B2(n_244),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_361),
.A2(n_363),
.B1(n_371),
.B2(n_373),
.Y(n_407)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_300),
.A2(n_252),
.B1(n_225),
.B2(n_296),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_253),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_370),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_311),
.B1(n_327),
.B2(n_343),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_232),
.B(n_251),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_379),
.B(n_395),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_346),
.B(n_235),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_369),
.B(n_372),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_336),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_270),
.Y(n_372)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_301),
.B(n_263),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_305),
.B(n_336),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_377),
.B(n_380),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_228),
.B1(n_261),
.B2(n_229),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_378),
.A2(n_311),
.B1(n_342),
.B2(n_303),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_231),
.B(n_286),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_267),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_307),
.A2(n_237),
.B(n_290),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_383),
.A2(n_400),
.B(n_402),
.Y(n_427)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_352),
.Y(n_384)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_305),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_385),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_333),
.B(n_281),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_386),
.B(n_394),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_344),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_389),
.Y(n_425)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_300),
.A2(n_5),
.B1(n_286),
.B2(n_329),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_391),
.B1(n_398),
.B2(n_399),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_307),
.A2(n_347),
.B1(n_349),
.B2(n_302),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_304),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_396),
.Y(n_435)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_5),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_331),
.A2(n_328),
.B(n_302),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_355),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_397),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_320),
.A2(n_338),
.B1(n_356),
.B2(n_355),
.Y(n_398)
);

OAI22x1_ASAP7_75t_SL g399 ( 
.A1(n_355),
.A2(n_330),
.B1(n_338),
.B2(n_314),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_339),
.A2(n_353),
.B(n_304),
.C(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_340),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_401),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_332),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_332),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_343),
.B(n_342),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_391),
.A2(n_390),
.B1(n_371),
.B2(n_398),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_409),
.A2(n_310),
.B(n_304),
.C(n_374),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_414),
.A2(n_359),
.B1(n_392),
.B2(n_388),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_426),
.B1(n_431),
.B2(n_383),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_400),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_422),
.B(n_433),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_364),
.A2(n_314),
.B1(n_324),
.B2(n_332),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_358),
.B(n_340),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_436),
.C(n_438),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_363),
.B1(n_361),
.B2(n_364),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_429),
.A2(n_432),
.B1(n_378),
.B2(n_373),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_396),
.A2(n_309),
.B1(n_299),
.B2(n_317),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_380),
.A2(n_299),
.B1(n_317),
.B2(n_354),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_400),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_308),
.C(n_354),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_365),
.B(n_343),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_439),
.B(n_383),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_386),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_438),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_425),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_442),
.B(n_450),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_436),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_446),
.Y(n_480)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_372),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_377),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_449),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_448),
.B(n_459),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_395),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_416),
.B(n_369),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_451),
.B(n_455),
.Y(n_499)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_393),
.C(n_384),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_461),
.C(n_471),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_454),
.A2(n_457),
.B1(n_462),
.B2(n_463),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_437),
.B(n_370),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_405),
.Y(n_456)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_456),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_427),
.A2(n_387),
.B(n_379),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_458),
.A2(n_427),
.B(n_422),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_406),
.B(n_308),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_460),
.B(n_464),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_394),
.C(n_402),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_409),
.A2(n_403),
.B1(n_362),
.B2(n_360),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_409),
.A2(n_368),
.B1(n_383),
.B2(n_375),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_425),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_429),
.A2(n_359),
.B1(n_401),
.B2(n_382),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_465),
.A2(n_407),
.B1(n_414),
.B2(n_418),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_466),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_431),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_467),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_468),
.A2(n_474),
.B(n_433),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_381),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_469),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_430),
.B(n_374),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_470),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_439),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_419),
.B(n_397),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_475),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_405),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_419),
.B(n_397),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_345),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_432),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_443),
.B(n_412),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_479),
.B(n_487),
.Y(n_525)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_486),
.A2(n_505),
.B(n_458),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_412),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_445),
.B(n_423),
.C(n_440),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_489),
.C(n_494),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_445),
.B(n_434),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_491),
.A2(n_468),
.B1(n_474),
.B2(n_472),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_492),
.A2(n_498),
.B1(n_502),
.B2(n_503),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_446),
.B(n_434),
.C(n_415),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_449),
.B(n_415),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_495),
.B(n_496),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_408),
.C(n_426),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_454),
.A2(n_407),
.B1(n_411),
.B2(n_418),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_465),
.A2(n_408),
.B1(n_424),
.B2(n_421),
.Y(n_502)
);

AOI211xp5_ASAP7_75t_L g503 ( 
.A1(n_473),
.A2(n_410),
.B(n_417),
.C(n_420),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_420),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_504),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_448),
.A2(n_424),
.B(n_410),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_462),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_464),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_442),
.B(n_417),
.C(n_413),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_456),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_503),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_512),
.B(n_513),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_501),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_514),
.B(n_521),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_486),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_515),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_499),
.B(n_469),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_516),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_517),
.A2(n_529),
.B(n_531),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_508),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_518),
.B(n_528),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_473),
.Y(n_519)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_519),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_505),
.Y(n_522)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_495),
.B(n_470),
.Y(n_523)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_483),
.A2(n_459),
.B1(n_468),
.B2(n_463),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_498),
.B1(n_478),
.B2(n_502),
.Y(n_555)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_476),
.Y(n_527)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_527),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_491),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_497),
.A2(n_466),
.B(n_468),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_530),
.B(n_532),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_497),
.A2(n_457),
.B(n_468),
.Y(n_531)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_494),
.B(n_474),
.C(n_475),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_534),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_477),
.A2(n_413),
.B(n_452),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_441),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_535),
.B(n_538),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_510),
.B(n_441),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_345),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_539),
.B(n_484),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_480),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_543),
.B(n_544),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_480),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_549),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_514),
.B(n_481),
.Y(n_547)
);

XNOR2x1_ASAP7_75t_L g572 ( 
.A(n_547),
.B(n_558),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_511),
.B(n_489),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_540),
.B(n_481),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_563),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_555),
.A2(n_564),
.B1(n_531),
.B2(n_548),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_540),
.B(n_479),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_530),
.B(n_487),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_512),
.A2(n_483),
.B1(n_478),
.B2(n_492),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_564),
.A2(n_536),
.B1(n_519),
.B2(n_529),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_561),
.A2(n_536),
.B1(n_531),
.B2(n_518),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_565),
.A2(n_567),
.B1(n_570),
.B2(n_580),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_561),
.A2(n_531),
.B1(n_524),
.B2(n_515),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_556),
.Y(n_571)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_571),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_511),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_574),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_488),
.C(n_537),
.Y(n_574)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_557),
.A2(n_517),
.B(n_506),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_576),
.Y(n_601)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_562),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_521),
.C(n_496),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_582),
.C(n_584),
.Y(n_599)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_542),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_578),
.B(n_583),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_560),
.A2(n_513),
.B(n_534),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_581),
.B(n_559),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_541),
.A2(n_522),
.B(n_528),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_544),
.B(n_504),
.C(n_485),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_563),
.B(n_485),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_520),
.C(n_539),
.Y(n_584)
);

BUFx24_ASAP7_75t_SL g585 ( 
.A(n_573),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_566),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_568),
.B(n_545),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_588),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_577),
.B(n_545),
.C(n_558),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_596),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_559),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_589),
.A2(n_594),
.B(n_598),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_569),
.B(n_552),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_600),
.Y(n_604)
);

OAI321xp33_ASAP7_75t_L g594 ( 
.A1(n_565),
.A2(n_553),
.A3(n_516),
.B1(n_490),
.B2(n_551),
.C(n_535),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_SL g595 ( 
.A(n_572),
.B(n_520),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_595),
.B(n_528),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_575),
.Y(n_596)
);

OAI321xp33_ASAP7_75t_L g598 ( 
.A1(n_570),
.A2(n_527),
.A3(n_554),
.B1(n_523),
.B2(n_555),
.C(n_538),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_546),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_593),
.A2(n_581),
.B1(n_528),
.B2(n_554),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_602),
.B(n_611),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_599),
.B(n_582),
.C(n_566),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_609),
.C(n_610),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_606),
.B(n_614),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_590),
.B(n_526),
.Y(n_608)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_608),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_586),
.C(n_574),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_587),
.B(n_583),
.C(n_584),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_601),
.A2(n_528),
.B1(n_572),
.B2(n_325),
.Y(n_611)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_612),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_325),
.Y(n_613)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_613),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_592),
.A2(n_325),
.B1(n_326),
.B2(n_339),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_607),
.A2(n_588),
.B(n_595),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_619),
.A2(n_611),
.B(n_602),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_605),
.B(n_600),
.Y(n_621)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_621),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_607),
.A2(n_326),
.B1(n_345),
.B2(n_323),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_615),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_609),
.B(n_310),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_625),
.B(n_615),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_627),
.Y(n_633)
);

BUFx4f_ASAP7_75t_SL g627 ( 
.A(n_617),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_603),
.C(n_610),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_629),
.B(n_631),
.Y(n_634)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_630),
.A2(n_624),
.B(n_616),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_620),
.B(n_604),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_632),
.A2(n_618),
.B(n_619),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_635),
.B(n_636),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_634),
.B(n_628),
.C(n_626),
.Y(n_638)
);

OAI21x1_ASAP7_75t_SL g639 ( 
.A1(n_638),
.A2(n_633),
.B(n_624),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_639),
.A2(n_627),
.B1(n_637),
.B2(n_623),
.Y(n_640)
);

NAND4xp25_ASAP7_75t_L g641 ( 
.A(n_640),
.B(n_627),
.C(n_622),
.D(n_625),
.Y(n_641)
);

AOI321xp33_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_604),
.A3(n_351),
.B1(n_310),
.B2(n_319),
.C(n_323),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_642),
.A2(n_351),
.B(n_319),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_351),
.B(n_392),
.Y(n_644)
);


endmodule