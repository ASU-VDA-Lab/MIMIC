module fake_jpeg_26720_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.C(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_17),
.B(n_27),
.C(n_23),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_22),
.B(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_17),
.B(n_27),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_54),
.B(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

OAI22x1_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_19),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_58),
.B1(n_29),
.B2(n_28),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_16),
.B1(n_26),
.B2(n_29),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_26),
.B1(n_16),
.B2(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_40),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_36),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_72),
.B(n_83),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_33),
.B1(n_30),
.B2(n_19),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_55),
.B(n_60),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_33),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_84),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_32),
.B1(n_24),
.B2(n_28),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_44),
.B(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_92),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_71),
.B1(n_49),
.B2(n_81),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_74),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_73),
.B(n_72),
.C(n_84),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_122),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_132),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_85),
.B1(n_76),
.B2(n_78),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_128),
.B1(n_107),
.B2(n_109),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_67),
.B1(n_70),
.B2(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_131),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_86),
.B(n_66),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_100),
.B(n_19),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_79),
.B1(n_71),
.B2(n_69),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_83),
.B1(n_75),
.B2(n_64),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_136),
.B1(n_94),
.B2(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_93),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_83),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_75),
.B1(n_49),
.B2(n_22),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_93),
.C(n_104),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_128),
.C(n_129),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

OAI211xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_96),
.B(n_95),
.C(n_104),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_156),
.B(n_157),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_90),
.B1(n_107),
.B2(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_103),
.B1(n_112),
.B2(n_18),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_96),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_106),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_130),
.B1(n_129),
.B2(n_114),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_124),
.C(n_123),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_119),
.B(n_134),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_147),
.B(n_144),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_164),
.C(n_138),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_165),
.B1(n_169),
.B2(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_131),
.C(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_135),
.B1(n_121),
.B2(n_103),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_121),
.A3(n_31),
.B1(n_18),
.B2(n_13),
.C1(n_15),
.C2(n_63),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_140),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_112),
.B1(n_31),
.B2(n_63),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_18),
.A3(n_47),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_165),
.B1(n_163),
.B2(n_150),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_175),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_183),
.B1(n_160),
.B2(n_161),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_178),
.C(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_144),
.C(n_154),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_185),
.B(n_146),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_173),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_137),
.B1(n_169),
.B2(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_145),
.B(n_147),
.C(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_191),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_168),
.C(n_158),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_195),
.C(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_158),
.C(n_167),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_184),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_189),
.B(n_8),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_180),
.B(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_9),
.C(n_10),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_142),
.B1(n_3),
.B2(n_4),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_189),
.B1(n_6),
.B2(n_7),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_2),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_210),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_2),
.C(n_9),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_210),
.CI(n_213),
.CON(n_217),
.SN(n_217)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_199),
.B(n_203),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_199),
.CI(n_208),
.CON(n_218),
.SN(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_208),
.Y(n_219)
);

OAI322xp33_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_220),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_217),
.C2(n_216),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_217),
.B(n_218),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_11),
.Y(n_222)
);


endmodule