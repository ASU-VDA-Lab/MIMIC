module real_aes_7155_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g231 ( .A1(n_0), .A2(n_232), .B(n_233), .C(n_237), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_1), .B(n_173), .Y(n_238) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_3), .B(n_145), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_4), .A2(n_131), .B(n_136), .C(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_5), .A2(n_126), .B(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_6), .A2(n_126), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_7), .B(n_173), .Y(n_544) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_8), .A2(n_161), .B(n_177), .Y(n_176) );
AND2x6_ASAP7_75t_L g131 ( .A(n_9), .B(n_132), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_10), .A2(n_131), .B(n_136), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g482 ( .A(n_11), .Y(n_482) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_12), .B(n_41), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_13), .B(n_236), .Y(n_502) );
INVx1_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_15), .B(n_145), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_16), .A2(n_146), .B(n_490), .C(n_492), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_17), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_18), .B(n_173), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_19), .B(n_210), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_20), .A2(n_136), .B(n_187), .C(n_206), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_21), .A2(n_185), .B(n_235), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_22), .B(n_236), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_23), .B(n_236), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_24), .Y(n_529) );
INVx1_ASAP7_75t_L g521 ( .A(n_25), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_26), .A2(n_136), .B(n_180), .C(n_187), .Y(n_179) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_27), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_28), .Y(n_498) );
INVx1_ASAP7_75t_L g578 ( .A(n_29), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_30), .A2(n_126), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g129 ( .A(n_31), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_32), .A2(n_134), .B(n_149), .C(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_33), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_34), .A2(n_235), .B(n_541), .C(n_543), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_35), .A2(n_100), .B1(n_111), .B2(n_749), .Y(n_99) );
INVxp67_ASAP7_75t_L g579 ( .A(n_36), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_37), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_38), .A2(n_136), .B(n_187), .C(n_520), .Y(n_519) );
CKINVDCx14_ASAP7_75t_R g539 ( .A(n_39), .Y(n_539) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_40), .A2(n_98), .B1(n_463), .B2(n_741), .C1(n_742), .C2(n_745), .Y(n_462) );
INVx1_ASAP7_75t_L g741 ( .A(n_40), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_41), .B(n_105), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_42), .A2(n_237), .B(n_480), .C(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_43), .B(n_204), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_44), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_45), .A2(n_118), .B1(n_119), .B2(n_449), .Y(n_117) );
INVx1_ASAP7_75t_L g449 ( .A(n_45), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_46), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_47), .B(n_126), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_48), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_49), .Y(n_575) );
A2O1A1Ixp33_ASAP7_75t_L g133 ( .A1(n_50), .A2(n_134), .B(n_139), .C(n_149), .Y(n_133) );
INVx1_ASAP7_75t_L g234 ( .A(n_51), .Y(n_234) );
INVx1_ASAP7_75t_L g140 ( .A(n_52), .Y(n_140) );
INVx1_ASAP7_75t_L g510 ( .A(n_53), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_54), .B(n_126), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_55), .Y(n_213) );
CKINVDCx14_ASAP7_75t_R g478 ( .A(n_56), .Y(n_478) );
INVx1_ASAP7_75t_L g132 ( .A(n_57), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_58), .B(n_126), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_59), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_60), .A2(n_167), .B(n_169), .C(n_171), .Y(n_166) );
INVx1_ASAP7_75t_L g154 ( .A(n_61), .Y(n_154) );
INVx1_ASAP7_75t_SL g542 ( .A(n_62), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_64), .B(n_145), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_65), .B(n_173), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_66), .B(n_146), .Y(n_248) );
INVx1_ASAP7_75t_L g532 ( .A(n_67), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_68), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_69), .B(n_142), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_70), .A2(n_136), .B(n_149), .C(n_219), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_71), .Y(n_165) );
INVx1_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_73), .A2(n_126), .B(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_74), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_75), .A2(n_126), .B(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_76), .A2(n_204), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g488 ( .A(n_77), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_78), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_79), .B(n_141), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_80), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_81), .A2(n_126), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g491 ( .A(n_82), .Y(n_491) );
INVx2_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
INVx1_ASAP7_75t_L g501 ( .A(n_84), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_85), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_86), .B(n_236), .Y(n_249) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_87), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g453 ( .A(n_87), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g469 ( .A(n_87), .Y(n_469) );
OR2x2_ASAP7_75t_L g740 ( .A(n_87), .B(n_455), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_88), .A2(n_136), .B(n_149), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_89), .B(n_126), .Y(n_193) );
INVx1_ASAP7_75t_L g196 ( .A(n_90), .Y(n_196) );
INVxp67_ASAP7_75t_L g170 ( .A(n_91), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_92), .B(n_161), .Y(n_483) );
INVx2_ASAP7_75t_L g513 ( .A(n_93), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_94), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g220 ( .A(n_95), .Y(n_220) );
INVx1_ASAP7_75t_L g244 ( .A(n_96), .Y(n_244) );
AND2x2_ASAP7_75t_L g156 ( .A(n_97), .B(n_151), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx5_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_103), .Y(n_750) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g455 ( .A(n_107), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_461), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g748 ( .A(n_115), .Y(n_748) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_450), .B(n_457), .Y(n_116) );
AOI22x1_ASAP7_75t_SL g746 ( .A1(n_118), .A2(n_465), .B1(n_737), .B2(n_747), .Y(n_746) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_119), .A2(n_465), .B1(n_470), .B2(n_737), .Y(n_464) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR5x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_322), .C(n_400), .D(n_424), .E(n_441), .Y(n_120) );
OAI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_188), .B(n_239), .C(n_299), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_157), .Y(n_122) );
AND2x2_ASAP7_75t_L g253 ( .A(n_123), .B(n_159), .Y(n_253) );
INVx5_ASAP7_75t_SL g281 ( .A(n_123), .Y(n_281) );
AND2x2_ASAP7_75t_L g317 ( .A(n_123), .B(n_302), .Y(n_317) );
OR2x2_ASAP7_75t_L g356 ( .A(n_123), .B(n_158), .Y(n_356) );
OR2x2_ASAP7_75t_L g387 ( .A(n_123), .B(n_278), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_123), .B(n_291), .Y(n_423) );
AND2x2_ASAP7_75t_L g435 ( .A(n_123), .B(n_278), .Y(n_435) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_156), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_133), .B(n_151), .Y(n_124) );
BUFx2_ASAP7_75t_L g204 ( .A(n_126), .Y(n_204) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_131), .Y(n_126) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_127), .B(n_131), .Y(n_245) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
INVx1_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
INVx1_ASAP7_75t_L g186 ( .A(n_129), .Y(n_186) );
INVx1_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_130), .Y(n_143) );
INVx3_ASAP7_75t_L g146 ( .A(n_130), .Y(n_146) );
INVx1_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_130), .Y(n_236) );
INVx4_ASAP7_75t_SL g150 ( .A(n_131), .Y(n_150) );
BUFx3_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_135), .A2(n_150), .B(n_165), .C(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g229 ( .A1(n_135), .A2(n_150), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_135), .A2(n_150), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g487 ( .A1(n_135), .A2(n_150), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_135), .A2(n_150), .B(n_510), .C(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_135), .A2(n_150), .B(n_539), .C(n_540), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_SL g574 ( .A1(n_135), .A2(n_150), .B(n_575), .C(n_576), .Y(n_574) );
INVx5_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx3_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_137), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_144), .C(n_147), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_141), .A2(n_147), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp5_ASAP7_75t_L g500 ( .A1(n_141), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_141), .A2(n_503), .B(n_532), .C(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_145), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g232 ( .A(n_145), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_145), .A2(n_209), .B(n_521), .C(n_522), .Y(n_520) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_145), .A2(n_168), .B1(n_578), .B2(n_579), .Y(n_577) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_146), .B(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g237 ( .A(n_148), .Y(n_237) );
INVx1_ASAP7_75t_L g492 ( .A(n_148), .Y(n_492) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_151), .A2(n_193), .B(n_194), .Y(n_192) );
INVx2_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
INVx1_ASAP7_75t_L g214 ( .A(n_151), .Y(n_214) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_151), .A2(n_476), .B(n_483), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_151), .A2(n_245), .B(n_518), .C(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_L g162 ( .A(n_152), .B(n_153), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g434 ( .A(n_157), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g297 ( .A(n_158), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_175), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_159), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_159), .Y(n_290) );
INVx3_ASAP7_75t_L g305 ( .A(n_159), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_159), .B(n_175), .Y(n_329) );
OR2x2_ASAP7_75t_L g338 ( .A(n_159), .B(n_281), .Y(n_338) );
AND2x2_ASAP7_75t_L g342 ( .A(n_159), .B(n_302), .Y(n_342) );
AND2x2_ASAP7_75t_L g348 ( .A(n_159), .B(n_349), .Y(n_348) );
INVxp67_ASAP7_75t_L g385 ( .A(n_159), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_159), .B(n_242), .Y(n_399) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_163), .B(n_172), .Y(n_159) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_160), .A2(n_486), .B(n_493), .Y(n_485) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_160), .A2(n_508), .B(n_514), .Y(n_507) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_160), .A2(n_537), .B(n_544), .Y(n_536) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_161), .A2(n_178), .B(n_179), .Y(n_177) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g252 ( .A(n_162), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_167), .A2(n_220), .B(n_221), .C(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_168), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_168), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_171), .B(n_577), .Y(n_576) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_173), .A2(n_228), .B(n_238), .Y(n_227) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_174), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_174), .A2(n_217), .B(n_225), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_174), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_174), .A2(n_243), .B(n_250), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_174), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_174), .B(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_174), .A2(n_528), .B(n_534), .Y(n_527) );
OR2x2_ASAP7_75t_L g291 ( .A(n_175), .B(n_242), .Y(n_291) );
AND2x2_ASAP7_75t_L g302 ( .A(n_175), .B(n_278), .Y(n_302) );
AND2x2_ASAP7_75t_L g314 ( .A(n_175), .B(n_305), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_175), .B(n_242), .Y(n_337) );
INVx1_ASAP7_75t_SL g349 ( .A(n_175), .Y(n_349) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g241 ( .A(n_176), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_176), .B(n_281), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .B(n_184), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_184), .A2(n_248), .B(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_200), .Y(n_189) );
AND2x2_ASAP7_75t_L g262 ( .A(n_190), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_190), .B(n_215), .Y(n_266) );
AND2x2_ASAP7_75t_L g269 ( .A(n_190), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_190), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g294 ( .A(n_190), .B(n_285), .Y(n_294) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_190), .Y(n_313) );
AND2x2_ASAP7_75t_L g334 ( .A(n_190), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g344 ( .A(n_190), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g390 ( .A(n_190), .B(n_273), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_190), .B(n_296), .Y(n_417) );
INVx5_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g287 ( .A(n_191), .Y(n_287) );
AND2x2_ASAP7_75t_L g353 ( .A(n_191), .B(n_285), .Y(n_353) );
AND2x2_ASAP7_75t_L g437 ( .A(n_191), .B(n_305), .Y(n_437) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_198), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_200), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_200), .Y(n_426) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_215), .Y(n_200) );
AND2x2_ASAP7_75t_L g256 ( .A(n_201), .B(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g265 ( .A(n_201), .B(n_263), .Y(n_265) );
INVx5_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
AND2x2_ASAP7_75t_L g296 ( .A(n_201), .B(n_227), .Y(n_296) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_201), .Y(n_333) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
AOI21xp5_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_205), .B(n_210), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .Y(n_206) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_211), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_214), .A2(n_497), .B(n_504), .Y(n_496) );
INVx1_ASAP7_75t_L g374 ( .A(n_215), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_215), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g407 ( .A(n_215), .B(n_273), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_215), .A2(n_330), .B(n_437), .C(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_227), .Y(n_215) );
BUFx2_ASAP7_75t_L g257 ( .A(n_216), .Y(n_257) );
INVx2_ASAP7_75t_L g261 ( .A(n_216), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g543 ( .A(n_223), .Y(n_543) );
INVx2_ASAP7_75t_L g263 ( .A(n_227), .Y(n_263) );
AND2x2_ASAP7_75t_L g270 ( .A(n_227), .B(n_261), .Y(n_270) );
AND2x2_ASAP7_75t_L g361 ( .A(n_227), .B(n_273), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_235), .B(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g480 ( .A(n_236), .Y(n_480) );
INVx2_ASAP7_75t_L g503 ( .A(n_237), .Y(n_503) );
AOI211x1_ASAP7_75t_SL g239 ( .A1(n_240), .A2(n_254), .B(n_267), .C(n_292), .Y(n_239) );
INVx1_ASAP7_75t_L g358 ( .A(n_240), .Y(n_358) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_253), .Y(n_240) );
INVx5_ASAP7_75t_SL g278 ( .A(n_242), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_242), .B(n_348), .Y(n_347) );
AOI311xp33_ASAP7_75t_L g366 ( .A1(n_242), .A2(n_367), .A3(n_369), .B(n_370), .C(n_376), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_242), .A2(n_314), .B(n_402), .C(n_405), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_246), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_245), .A2(n_498), .B(n_499), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_245), .A2(n_529), .B(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g571 ( .A(n_252), .Y(n_571) );
INVxp67_ASAP7_75t_L g321 ( .A(n_253), .Y(n_321) );
NAND4xp25_ASAP7_75t_SL g254 ( .A(n_255), .B(n_258), .C(n_264), .D(n_266), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_255), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g312 ( .A(n_256), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_259), .B(n_265), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_259), .B(n_272), .Y(n_392) );
BUFx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_260), .B(n_273), .Y(n_410) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g285 ( .A(n_261), .Y(n_285) );
INVxp67_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
AND2x4_ASAP7_75t_L g272 ( .A(n_263), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g346 ( .A(n_263), .B(n_285), .Y(n_346) );
INVx1_ASAP7_75t_L g373 ( .A(n_263), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_263), .B(n_360), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_264), .B(n_334), .Y(n_354) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_265), .B(n_287), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_265), .B(n_334), .Y(n_433) );
INVx1_ASAP7_75t_L g444 ( .A(n_266), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_274), .C(n_282), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g286 ( .A(n_270), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g324 ( .A(n_270), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g306 ( .A(n_271), .Y(n_306) );
AND2x2_ASAP7_75t_L g283 ( .A(n_272), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_272), .B(n_334), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_272), .B(n_353), .Y(n_377) );
OR2x2_ASAP7_75t_L g293 ( .A(n_273), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g325 ( .A(n_273), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_273), .B(n_285), .Y(n_340) );
AND2x2_ASAP7_75t_L g397 ( .A(n_273), .B(n_353), .Y(n_397) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_273), .Y(n_404) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_275), .A2(n_287), .B1(n_409), .B2(n_411), .C(n_414), .Y(n_408) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g298 ( .A(n_278), .B(n_281), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_278), .B(n_348), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_278), .B(n_305), .Y(n_413) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g398 ( .A(n_280), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g412 ( .A(n_280), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_281), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g309 ( .A(n_281), .B(n_302), .Y(n_309) );
AND2x2_ASAP7_75t_L g379 ( .A(n_281), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_281), .B(n_328), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_281), .B(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_286), .B(n_288), .Y(n_282) );
INVx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g335 ( .A(n_285), .Y(n_335) );
OR2x2_ASAP7_75t_L g339 ( .A(n_287), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g442 ( .A(n_287), .B(n_410), .Y(n_442) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI21xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_L g446 ( .A(n_293), .Y(n_446) );
INVx2_ASAP7_75t_SL g360 ( .A(n_294), .Y(n_360) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_297), .A2(n_378), .B(n_442), .C(n_443), .Y(n_441) );
OAI322xp33_ASAP7_75t_SL g310 ( .A1(n_298), .A2(n_311), .A3(n_314), .B1(n_315), .B2(n_316), .C1(n_318), .C2(n_321), .Y(n_310) );
INVx2_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_307), .B2(n_309), .C(n_310), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI22xp33_ASAP7_75t_SL g376 ( .A1(n_301), .A2(n_377), .B1(n_378), .B2(n_381), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_302), .B(n_305), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_302), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g375 ( .A(n_304), .B(n_337), .Y(n_375) );
INVx1_ASAP7_75t_L g365 ( .A(n_305), .Y(n_365) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_309), .A2(n_419), .B(n_421), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_311), .A2(n_344), .B(n_347), .Y(n_343) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp67_ASAP7_75t_SL g372 ( .A(n_313), .B(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_313), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g429 ( .A(n_314), .Y(n_429) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND4xp25_ASAP7_75t_L g322 ( .A(n_323), .B(n_350), .C(n_366), .D(n_382), .Y(n_322) );
AOI211xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B(n_331), .C(n_343), .Y(n_323) );
INVx1_ASAP7_75t_L g415 ( .A(n_324), .Y(n_415) );
AND2x2_ASAP7_75t_L g363 ( .A(n_325), .B(n_346), .Y(n_363) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_330), .B(n_365), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_336), .B1(n_339), .B2(n_341), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_333), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_334), .A2(n_373), .B(n_396), .C(n_398), .Y(n_395) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
INVx1_ASAP7_75t_L g440 ( .A(n_338), .Y(n_440) );
NAND2xp33_ASAP7_75t_SL g430 ( .A(n_339), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B(n_355), .C(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_362), .B2(n_364), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_360), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_365), .B(n_386), .Y(n_448) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI21xp33_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_374), .B(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_388), .B1(n_391), .B2(n_393), .C(n_395), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_398), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_414) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_408), .C(n_418), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B(n_427), .C(n_436), .Y(n_424) );
INVx1_ASAP7_75t_L g445 ( .A(n_425), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_432), .B2(n_434), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g460 ( .A(n_453), .Y(n_460) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_454), .B(n_469), .Y(n_744) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g468 ( .A(n_455), .B(n_469), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_457), .B(n_462), .C(n_748), .Y(n_461) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g747 ( .A(n_470), .Y(n_747) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_667), .Y(n_470) );
NAND5xp2_ASAP7_75t_L g471 ( .A(n_472), .B(n_582), .C(n_614), .D(n_631), .E(n_654), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_515), .B1(n_545), .B2(n_549), .C(n_553), .Y(n_472) );
INVx1_ASAP7_75t_L g694 ( .A(n_473), .Y(n_694) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_494), .Y(n_473) );
AND3x2_ASAP7_75t_L g669 ( .A(n_474), .B(n_496), .C(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_475), .B(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g560 ( .A(n_475), .Y(n_560) );
AND2x2_ASAP7_75t_L g564 ( .A(n_475), .B(n_506), .Y(n_564) );
INVx2_ASAP7_75t_L g591 ( .A(n_475), .Y(n_591) );
OR2x2_ASAP7_75t_L g602 ( .A(n_475), .B(n_507), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_475), .B(n_495), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_475), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g681 ( .A(n_475), .B(n_507), .Y(n_681) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_484), .Y(n_563) );
AND2x2_ASAP7_75t_L g622 ( .A(n_484), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_484), .B(n_495), .Y(n_641) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g552 ( .A(n_485), .B(n_495), .Y(n_552) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
AND2x2_ASAP7_75t_L g608 ( .A(n_485), .B(n_507), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_485), .B(n_494), .C(n_591), .Y(n_633) );
AND2x2_ASAP7_75t_L g698 ( .A(n_485), .B(n_496), .Y(n_698) );
AND2x2_ASAP7_75t_L g732 ( .A(n_485), .B(n_495), .Y(n_732) );
INVxp67_ASAP7_75t_L g561 ( .A(n_494), .Y(n_561) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_495), .B(n_591), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_495), .B(n_622), .Y(n_630) );
AND2x2_ASAP7_75t_L g680 ( .A(n_495), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g708 ( .A(n_495), .Y(n_708) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g615 ( .A(n_496), .B(n_608), .Y(n_615) );
BUFx3_ASAP7_75t_L g647 ( .A(n_496), .Y(n_647) );
INVx2_ASAP7_75t_L g623 ( .A(n_506), .Y(n_623) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_507), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_515), .A2(n_683), .B1(n_685), .B2(n_686), .Y(n_682) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
AND2x2_ASAP7_75t_L g545 ( .A(n_516), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_SL g556 ( .A(n_516), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_516), .B(n_586), .Y(n_618) );
OR2x2_ASAP7_75t_L g637 ( .A(n_516), .B(n_526), .Y(n_637) );
AND2x2_ASAP7_75t_L g642 ( .A(n_516), .B(n_594), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_516), .B(n_587), .Y(n_645) );
AND2x2_ASAP7_75t_L g657 ( .A(n_516), .B(n_536), .Y(n_657) );
AND2x2_ASAP7_75t_L g673 ( .A(n_516), .B(n_527), .Y(n_673) );
AND2x4_ASAP7_75t_L g676 ( .A(n_516), .B(n_547), .Y(n_676) );
OR2x2_ASAP7_75t_L g693 ( .A(n_516), .B(n_629), .Y(n_693) );
OR2x2_ASAP7_75t_L g724 ( .A(n_516), .B(n_569), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_516), .B(n_652), .Y(n_726) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
AND2x2_ASAP7_75t_L g600 ( .A(n_525), .B(n_567), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_525), .B(n_587), .Y(n_719) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_536), .Y(n_525) );
AND2x2_ASAP7_75t_L g555 ( .A(n_526), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g586 ( .A(n_526), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g594 ( .A(n_526), .B(n_569), .Y(n_594) );
AND2x2_ASAP7_75t_L g612 ( .A(n_526), .B(n_547), .Y(n_612) );
OR2x2_ASAP7_75t_L g629 ( .A(n_526), .B(n_587), .Y(n_629) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g548 ( .A(n_527), .Y(n_548) );
AND2x2_ASAP7_75t_L g652 ( .A(n_527), .B(n_536), .Y(n_652) );
INVx2_ASAP7_75t_L g547 ( .A(n_536), .Y(n_547) );
INVx1_ASAP7_75t_L g664 ( .A(n_536), .Y(n_664) );
AND2x2_ASAP7_75t_L g714 ( .A(n_536), .B(n_556), .Y(n_714) );
AND2x2_ASAP7_75t_L g566 ( .A(n_546), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g598 ( .A(n_546), .B(n_556), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_546), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g585 ( .A(n_547), .B(n_556), .Y(n_585) );
OR2x2_ASAP7_75t_L g701 ( .A(n_548), .B(n_675), .Y(n_701) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_551), .B(n_681), .Y(n_687) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_552), .A2(n_644), .A3(n_646), .B1(n_648), .B2(n_649), .Y(n_643) );
OR2x2_ASAP7_75t_L g660 ( .A(n_552), .B(n_602), .Y(n_660) );
OAI21xp33_ASAP7_75t_SL g685 ( .A1(n_552), .A2(n_562), .B(n_590), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_557), .B1(n_562), .B2(n_565), .Y(n_553) );
INVxp33_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_555), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_556), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_556), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g711 ( .A(n_556), .B(n_652), .Y(n_711) );
OR2x2_ASAP7_75t_L g735 ( .A(n_556), .B(n_629), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g718 ( .A1(n_557), .A2(n_617), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g595 ( .A(n_559), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_559), .B(n_564), .Y(n_613) );
AND2x2_ASAP7_75t_L g635 ( .A(n_560), .B(n_608), .Y(n_635) );
INVx1_ASAP7_75t_L g648 ( .A(n_560), .Y(n_648) );
OR2x2_ASAP7_75t_L g653 ( .A(n_560), .B(n_587), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_563), .B(n_602), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_564), .A2(n_584), .B1(n_589), .B2(n_593), .Y(n_583) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_567), .A2(n_626), .B1(n_633), .B2(n_634), .Y(n_632) );
AND2x2_ASAP7_75t_L g710 ( .A(n_567), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_569), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g729 ( .A(n_569), .B(n_612), .Y(n_729) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B(n_580), .Y(n_569) );
INVx1_ASAP7_75t_L g588 ( .A(n_570), .Y(n_588) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_573), .A2(n_581), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_595), .B1(n_596), .B2(n_601), .C(n_603), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_585), .B(n_587), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_585), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g604 ( .A(n_586), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_586), .A2(n_692), .B(n_693), .C(n_694), .Y(n_691) );
AND2x2_ASAP7_75t_L g696 ( .A(n_586), .B(n_676), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_SL g734 ( .A1(n_586), .A2(n_675), .B(n_735), .C(n_736), .Y(n_734) );
BUFx3_ASAP7_75t_L g626 ( .A(n_587), .Y(n_626) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_590), .B(n_647), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_590), .A2(n_710), .B(n_712), .C(n_718), .Y(n_709) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVxp67_ASAP7_75t_L g670 ( .A(n_592), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_594), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g614 ( .A1(n_598), .A2(n_615), .B(n_616), .C(n_624), .Y(n_614) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g699 ( .A(n_602), .Y(n_699) );
OR2x2_ASAP7_75t_L g716 ( .A(n_602), .B(n_646), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_610), .B2(n_613), .Y(n_603) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_605), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
OR2x2_ASAP7_75t_L g703 ( .A(n_607), .B(n_647), .Y(n_703) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g658 ( .A(n_608), .B(n_648), .Y(n_658) );
INVx1_ASAP7_75t_L g666 ( .A(n_609), .Y(n_666) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_612), .B(n_626), .Y(n_674) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_622), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g731 ( .A(n_623), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_630), .Y(n_624) );
INVx1_ASAP7_75t_L g661 ( .A(n_625), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_626), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_626), .B(n_657), .Y(n_656) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_626), .B(n_652), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_626), .B(n_673), .Y(n_684) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_626), .A2(n_636), .B(n_676), .C(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_636), .B1(n_638), .B2(n_642), .C(n_643), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_640), .B(n_648), .Y(n_722) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g733 ( .A1(n_642), .A2(n_657), .B(n_659), .C(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_645), .B(n_652), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_646), .B(n_699), .Y(n_736) );
CKINVDCx16_ASAP7_75t_R g646 ( .A(n_647), .Y(n_646) );
INVxp33_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
AOI21xp33_ASAP7_75t_SL g662 ( .A1(n_651), .A2(n_663), .B(n_665), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_651), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_652), .B(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_659), .B2(n_661), .C(n_662), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_658), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g692 ( .A(n_664), .Y(n_692) );
NAND5xp2_ASAP7_75t_L g667 ( .A(n_668), .B(n_695), .C(n_709), .D(n_720), .E(n_733), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_678), .C(n_691), .Y(n_668) );
INVx2_ASAP7_75t_SL g715 ( .A(n_669), .Y(n_715) );
NAND4xp25_ASAP7_75t_SL g671 ( .A(n_672), .B(n_674), .C(n_675), .D(n_677), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g678 ( .A1(n_677), .A2(n_679), .B(n_682), .C(n_688), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_680), .A2(n_721), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_720) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_697), .B1(n_700), .B2(n_702), .C(n_704), .Y(n_695) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_703), .A2(n_726), .B1(n_728), .B2(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
endmodule