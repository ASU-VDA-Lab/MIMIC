module fake_jpeg_2774_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_10),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_14),
.B(n_2),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_46),
.Y(n_130)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_53),
.B(n_64),
.Y(n_105)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_56),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx3_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_63),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_33),
.B(n_12),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_11),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_80),
.Y(n_96)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_84),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_79),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_25),
.B(n_11),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_10),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_85),
.B(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_34),
.B(n_0),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_93),
.Y(n_98)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_28),
.B1(n_41),
.B2(n_30),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_0),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_28),
.B1(n_41),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_108),
.A2(n_112),
.B1(n_117),
.B2(n_119),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_46),
.A2(n_40),
.B1(n_35),
.B2(n_26),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_129),
.B1(n_135),
.B2(n_147),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_40),
.B1(n_35),
.B2(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_74),
.A2(n_42),
.B1(n_39),
.B2(n_20),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_122),
.A2(n_128),
.B1(n_8),
.B2(n_124),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_52),
.A2(n_39),
.B1(n_62),
.B2(n_36),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_126),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_54),
.A2(n_36),
.B1(n_20),
.B2(n_35),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_57),
.A2(n_40),
.B1(n_26),
.B2(n_23),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_49),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_23),
.B1(n_2),
.B2(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_58),
.B1(n_61),
.B2(n_82),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_49),
.A2(n_0),
.B1(n_4),
.B2(n_7),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_9),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_8),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_0),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_50),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_50),
.A2(n_8),
.B1(n_58),
.B2(n_81),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_149),
.B(n_151),
.Y(n_194)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_91),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_154),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_70),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_159),
.B(n_188),
.Y(n_223)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_130),
.B1(n_58),
.B2(n_115),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_165),
.A2(n_176),
.B1(n_175),
.B2(n_153),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_78),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_167),
.B(n_172),
.Y(n_229)
);

BUFx2_ASAP7_75t_SL g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2x1_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_83),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_176),
.B(n_187),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_98),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_84),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_65),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_123),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_96),
.B(n_8),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_186),
.Y(n_224)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_97),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_99),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_133),
.B1(n_125),
.B2(n_120),
.Y(n_227)
);

CKINVDCx12_ASAP7_75t_R g182 ( 
.A(n_104),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_190),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_95),
.B(n_116),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_138),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_119),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_132),
.B1(n_121),
.B2(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_141),
.Y(n_188)
);

NAND2x1_ASAP7_75t_SL g189 ( 
.A(n_106),
.B(n_148),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_113),
.B(n_140),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_113),
.Y(n_201)
);

NOR4xp25_ASAP7_75t_SL g192 ( 
.A(n_99),
.B(n_97),
.C(n_138),
.D(n_140),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_202),
.B(n_215),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_134),
.B1(n_103),
.B2(n_143),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_227),
.B1(n_187),
.B2(n_162),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_138),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_100),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_210),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_100),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_133),
.C(n_143),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_214),
.C(n_226),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_114),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_120),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_184),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_114),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_189),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_174),
.B(n_114),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_239),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_231),
.B(n_232),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

AO21x2_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_192),
.B(n_165),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_188),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_247),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_244),
.B1(n_217),
.B2(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_166),
.B1(n_175),
.B2(n_181),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_245),
.A2(n_246),
.B(n_251),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_193),
.A2(n_189),
.B(n_171),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_150),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_256),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_193),
.A2(n_180),
.B(n_154),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_152),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_254),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_163),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_160),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_258),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_201),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_259),
.A2(n_213),
.B1(n_196),
.B2(n_226),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_279),
.B1(n_257),
.B2(n_242),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_196),
.B(n_199),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_264),
.B(n_270),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_199),
.B(n_220),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_227),
.B1(n_226),
.B2(n_229),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_229),
.B(n_194),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_194),
.B1(n_145),
.B2(n_125),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_145),
.B1(n_195),
.B2(n_208),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_285),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_237),
.A2(n_195),
.B1(n_219),
.B2(n_221),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_230),
.B(n_239),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_237),
.A2(n_228),
.B1(n_208),
.B2(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_237),
.A2(n_238),
.B1(n_243),
.B2(n_248),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_240),
.B1(n_236),
.B2(n_241),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_237),
.A2(n_228),
.A3(n_203),
.B1(n_206),
.B2(n_178),
.C1(n_225),
.C2(n_200),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_283),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_294),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_252),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_289),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_249),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_304),
.B1(n_311),
.B2(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_258),
.B1(n_250),
.B2(n_234),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_260),
.B1(n_278),
.B2(n_280),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_254),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_249),
.C(n_231),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_275),
.A2(n_233),
.B(n_235),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_301),
.A2(n_296),
.B1(n_276),
.B2(n_271),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_256),
.C(n_255),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_200),
.C(n_225),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_278),
.A2(n_221),
.B1(n_228),
.B2(n_197),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_197),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_305),
.B(n_308),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_225),
.C(n_206),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_280),
.C(n_286),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_222),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_307),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_267),
.B(n_270),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_275),
.A2(n_203),
.B(n_179),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_264),
.C(n_267),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_332),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_263),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_314),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_288),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_297),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_315),
.B(n_293),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_316),
.A2(n_320),
.B1(n_311),
.B2(n_294),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_272),
.B1(n_273),
.B2(n_269),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_261),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_SL g343 ( 
.A(n_322),
.B(n_328),
.C(n_309),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_329),
.Y(n_336)
);

XOR2x2_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_262),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_263),
.C(n_271),
.Y(n_329)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_276),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_330),
.A2(n_296),
.B1(n_301),
.B2(n_300),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_306),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_337),
.B(n_349),
.Y(n_355)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_348),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_307),
.Y(n_341)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_333),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_342),
.B(n_344),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_312),
.B(n_326),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_265),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_313),
.B(n_329),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_310),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_321),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_332),
.Y(n_352)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_347),
.A2(n_317),
.B1(n_328),
.B2(n_322),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_353),
.A2(n_334),
.B1(n_346),
.B2(n_191),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_362),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_335),
.A2(n_283),
.B(n_291),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_345),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_360),
.B(n_365),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_286),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_277),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_277),
.C(n_222),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_366),
.B(n_334),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_336),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_369),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_347),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_374),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_351),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_373),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_345),
.B1(n_343),
.B2(n_340),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_376),
.A2(n_377),
.B1(n_363),
.B2(n_354),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_356),
.C(n_366),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_382),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_357),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_370),
.B(n_362),
.Y(n_383)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_383),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_384),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_370),
.B(n_361),
.Y(n_385)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_385),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_353),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_386),
.A2(n_387),
.B(n_164),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_359),
.B(n_179),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_381),
.B(n_373),
.CI(n_157),
.CON(n_389),
.SN(n_389)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_389),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_391),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_157),
.C(n_379),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_394),
.A2(n_395),
.B(n_391),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_157),
.C(n_386),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_392),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_397),
.B(n_398),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_392),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_400),
.A2(n_393),
.B1(n_388),
.B2(n_389),
.Y(n_403)
);

AOI322xp5_ASAP7_75t_L g402 ( 
.A1(n_396),
.A2(n_388),
.A3(n_389),
.B1(n_393),
.B2(n_394),
.C1(n_395),
.C2(n_399),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_402),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_403),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_401),
.B(n_388),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_405),
.Y(n_407)
);


endmodule