module fake_jpeg_9195_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_24),
.B1(n_14),
.B2(n_15),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_16),
.B2(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_33),
.B(n_2),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_47),
.B(n_25),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_26),
.B(n_21),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_57),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_19),
.B1(n_44),
.B2(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_60),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_13),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_65),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_21),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_13),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_83),
.B(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_58),
.B1(n_57),
.B2(n_35),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_86),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_28),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_28),
.C(n_13),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_55),
.C(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_12),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_12),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_93),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_68),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_59),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_101),
.C(n_26),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_66),
.B1(n_62),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_85),
.B1(n_22),
.B2(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_100),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_106),
.B(n_22),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_66),
.A3(n_54),
.B1(n_21),
.B2(n_22),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_80),
.B1(n_69),
.B2(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_35),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_11),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_72),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_113),
.B(n_118),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_69),
.B1(n_103),
.B2(n_76),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_119),
.C(n_101),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_73),
.B1(n_56),
.B2(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_121),
.B1(n_106),
.B2(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_11),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_124),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_98),
.B(n_93),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_137),
.B1(n_112),
.B2(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_131),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_134),
.C(n_115),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_94),
.C(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_96),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_136),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_102),
.C(n_91),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_116),
.B(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_72),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_145),
.B(n_146),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_133),
.B(n_122),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_147),
.C(n_134),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_116),
.C(n_121),
.Y(n_147)
);

OAI31xp33_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_130),
.A3(n_137),
.B(n_138),
.Y(n_151)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_130),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_154),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_6),
.B(n_7),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_146),
.B(n_145),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_5),
.C(n_6),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_7),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_156),
.C(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_154),
.B(n_8),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_157),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_167),
.B1(n_160),
.B2(n_8),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_150),
.C(n_9),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_10),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_10),
.B(n_160),
.C(n_168),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_10),
.B(n_171),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_173),
.Y(n_176)
);


endmodule