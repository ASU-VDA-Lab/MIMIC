module fake_ariane_2768_n_1868 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_457, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_1868);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_1868;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_533;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1716;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_489;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1208;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_673;
wire n_1038;
wire n_571;
wire n_1521;
wire n_1694;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_946;
wire n_757;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_1299;
wire n_782;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g459 ( 
.A(n_250),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_288),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_305),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_204),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_430),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_424),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_302),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_378),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_335),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_143),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_307),
.Y(n_470)
);

BUFx5_ASAP7_75t_L g471 ( 
.A(n_72),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_169),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_53),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_98),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_249),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_245),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_161),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_121),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_281),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_139),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_20),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_237),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_269),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_78),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_258),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_94),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_238),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_85),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_264),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_75),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_452),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_216),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_209),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_73),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_54),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_370),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_271),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_70),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_12),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_314),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_215),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_225),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_179),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_27),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_317),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_223),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_219),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_323),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_59),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_360),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_297),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_189),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_299),
.Y(n_515)
);

BUFx5_ASAP7_75t_L g516 ( 
.A(n_273),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_201),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_268),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_112),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_243),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_457),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_295),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_311),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_139),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_35),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_220),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_165),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_137),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_287),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_60),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_188),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_35),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_87),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_254),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_255),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_5),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_168),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_455),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_200),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_29),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_419),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_224),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_75),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_189),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_244),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_313),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_285),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_218),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_193),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_262),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_66),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_284),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_202),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_355),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_414),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_372),
.Y(n_558)
);

BUFx10_ASAP7_75t_L g559 ( 
.A(n_300),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_228),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_195),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_214),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_130),
.Y(n_563)
);

XNOR2x1_ASAP7_75t_L g564 ( 
.A(n_261),
.B(n_308),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_61),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_55),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_150),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_84),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_278),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_16),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_458),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_283),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_319),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_445),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_451),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_332),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_83),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_10),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_272),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_453),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_337),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_324),
.Y(n_582)
);

BUFx5_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_156),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_333),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_399),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_136),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_303),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_279),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_294),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_183),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_446),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_301),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_420),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_208),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_428),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_309),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_363),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_184),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_263),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_129),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_253),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_61),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_89),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_374),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_213),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_233),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_231),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_346),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_9),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_197),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_210),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_405),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_298),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_235),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_227),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_182),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_293),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_13),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_267),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_246),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_111),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_142),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_296),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_384),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_4),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_450),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_198),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_40),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_280),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_230),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_622),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_604),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_469),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

INVxp33_ASAP7_75t_SL g637 ( 
.A(n_604),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_469),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_569),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_473),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_620),
.Y(n_642)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_487),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_620),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_471),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_471),
.Y(n_646)
);

INVxp67_ASAP7_75t_SL g647 ( 
.A(n_542),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_472),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_578),
.B(n_0),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_477),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_481),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_492),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_513),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_500),
.Y(n_654)
);

INVxp33_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_543),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_519),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_529),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_524),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_530),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_551),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_532),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_534),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_535),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_524),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_546),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_577),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_542),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_574),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_624),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_601),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_603),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_506),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_542),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_542),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_511),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_525),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_571),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_501),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_580),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_531),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_531),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_578),
.Y(n_686)
);

CKINVDCx16_ASAP7_75t_R g687 ( 
.A(n_557),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_556),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_557),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_559),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_564),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_585),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_559),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_514),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_600),
.Y(n_695)
);

INVxp33_ASAP7_75t_SL g696 ( 
.A(n_474),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_600),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_502),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_459),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_556),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_462),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_478),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_598),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_598),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_465),
.Y(n_705)
);

CKINVDCx16_ASAP7_75t_R g706 ( 
.A(n_625),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_475),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_479),
.Y(n_708)
);

INVxp33_ASAP7_75t_SL g709 ( 
.A(n_480),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_484),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_491),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_631),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_498),
.Y(n_713)
);

INVxp33_ASAP7_75t_L g714 ( 
.A(n_482),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_504),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_517),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_637),
.A2(n_563),
.B1(n_545),
.B2(n_496),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_645),
.A2(n_527),
.B(n_526),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_703),
.B(n_528),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_643),
.B(n_655),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_640),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_640),
.Y(n_722)
);

INVx6_ASAP7_75t_L g723 ( 
.A(n_640),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_643),
.B(n_605),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_638),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_698),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_647),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_SL g728 ( 
.A(n_687),
.B(n_486),
.Y(n_728)
);

BUFx8_ASAP7_75t_L g729 ( 
.A(n_649),
.Y(n_729)
);

BUFx12f_ASAP7_75t_L g730 ( 
.A(n_653),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_670),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_698),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_698),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_714),
.B(n_549),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_677),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_714),
.B(n_550),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_646),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_678),
.Y(n_738)
);

OAI22x1_ASAP7_75t_L g739 ( 
.A1(n_633),
.A2(n_497),
.B1(n_505),
.B2(n_485),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_688),
.B(n_558),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_634),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_691),
.A2(n_673),
.B1(n_635),
.B2(n_641),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_655),
.B(n_538),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_634),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_688),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_700),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_700),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_704),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_650),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_704),
.B(n_502),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_699),
.B(n_483),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_701),
.Y(n_752)
);

BUFx12f_ASAP7_75t_L g753 ( 
.A(n_656),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_705),
.B(n_490),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_686),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_651),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_707),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_708),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_654),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_710),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_657),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_711),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_702),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_713),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_715),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_755),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_R g767 ( 
.A(n_725),
.B(n_661),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_749),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_730),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_730),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_R g771 ( 
.A(n_720),
.B(n_672),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_741),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_753),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_756),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_720),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_R g776 ( 
.A(n_743),
.B(n_683),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_741),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_724),
.B(n_684),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_753),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_759),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_725),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_717),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_724),
.B(n_685),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_763),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_761),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_762),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_742),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_746),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_728),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_729),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_729),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_729),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_744),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_743),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_751),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_757),
.B(n_692),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_765),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_765),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_737),
.B(n_689),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_734),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_765),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_746),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_736),
.A2(n_639),
.B1(n_642),
.B2(n_636),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_746),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_747),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_747),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_748),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_751),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_747),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_744),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_745),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_752),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_R g814 ( 
.A(n_718),
.B(n_712),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_744),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_748),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_752),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_R g818 ( 
.A(n_757),
.B(n_706),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_752),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_739),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_758),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_739),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_727),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_744),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_745),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_731),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_735),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_719),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_745),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_738),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_738),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_772),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_828),
.B(n_751),
.Y(n_833)
);

XOR2xp5_ASAP7_75t_L g834 ( 
.A(n_766),
.B(n_652),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_783),
.B(n_754),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_819),
.B(n_794),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_777),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_768),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_797),
.B(n_696),
.Y(n_839)
);

OAI22xp33_ASAP7_75t_L g840 ( 
.A1(n_782),
.A2(n_644),
.B1(n_666),
.B2(n_659),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_784),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_775),
.B(n_709),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_767),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_774),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_780),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_801),
.B(n_690),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_785),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_821),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_767),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_808),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_816),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_783),
.B(n_760),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_812),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_823),
.B(n_826),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_829),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_825),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_803),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_830),
.Y(n_858)
);

BUFx4f_ASAP7_75t_L g859 ( 
.A(n_786),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_796),
.B(n_764),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_805),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_831),
.Y(n_862)
);

AND2x6_ASAP7_75t_L g863 ( 
.A(n_815),
.B(n_764),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_793),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_813),
.B(n_658),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_781),
.B(n_693),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_769),
.Y(n_867)
);

AO22x2_ASAP7_75t_L g868 ( 
.A1(n_789),
.A2(n_681),
.B1(n_697),
.B2(n_695),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_778),
.B(n_666),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_791),
.B(n_660),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_809),
.B(n_716),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_827),
.B(n_740),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_815),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_809),
.B(n_818),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_811),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_804),
.B(n_539),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_770),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_800),
.B(n_682),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_795),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_824),
.B(n_503),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_773),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_787),
.B(n_682),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_818),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_779),
.Y(n_884)
);

AO22x2_ASAP7_75t_L g885 ( 
.A1(n_820),
.A2(n_694),
.B1(n_674),
.B2(n_648),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_798),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_792),
.B(n_632),
.Y(n_887)
);

INVx6_ASAP7_75t_L g888 ( 
.A(n_811),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_771),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_799),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_802),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_790),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_788),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_806),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_771),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_807),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_776),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_810),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_822),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_662),
.Y(n_900)
);

AND2x2_ASAP7_75t_SL g901 ( 
.A(n_814),
.B(n_694),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_814),
.B(n_553),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_R g903 ( 
.A(n_767),
.B(n_663),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_811),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_784),
.B(n_664),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_784),
.B(n_665),
.Y(n_906)
);

INVx5_ASAP7_75t_L g907 ( 
.A(n_809),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_768),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_793),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_782),
.A2(n_584),
.B1(n_565),
.B2(n_566),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_784),
.B(n_667),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_768),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_768),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_772),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_772),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_768),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_766),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_811),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_793),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_772),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_784),
.B(n_668),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_784),
.B(n_669),
.Y(n_922)
);

OAI22xp33_ASAP7_75t_SL g923 ( 
.A1(n_782),
.A2(n_570),
.B1(n_599),
.B2(n_587),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_817),
.B(n_568),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_828),
.B(n_610),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_832),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_838),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_841),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_843),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_867),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_844),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_854),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_856),
.A2(n_619),
.B1(n_623),
.B2(n_617),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_867),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_845),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_917),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_837),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_907),
.B(n_671),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_847),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_907),
.B(n_675),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_902),
.B(n_626),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_L g942 ( 
.A(n_849),
.B(n_629),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_907),
.B(n_874),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_842),
.A2(n_562),
.B(n_572),
.C(n_560),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_908),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_SL g946 ( 
.A1(n_834),
.A2(n_679),
.B1(n_680),
.B2(n_676),
.Y(n_946)
);

OR2x6_ASAP7_75t_L g947 ( 
.A(n_883),
.B(n_509),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_921),
.B(n_0),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_912),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_900),
.B(n_630),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_835),
.B(n_573),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_877),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_SL g953 ( 
.A1(n_882),
.A2(n_846),
.B1(n_878),
.B2(n_897),
.Y(n_953)
);

AO22x2_ASAP7_75t_L g954 ( 
.A1(n_900),
.A2(n_588),
.B1(n_592),
.B2(n_576),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_905),
.B(n_1),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_857),
.B(n_721),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_913),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_881),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_916),
.Y(n_959)
);

AO22x2_ASAP7_75t_L g960 ( 
.A1(n_901),
.A2(n_594),
.B1(n_595),
.B2(n_593),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_914),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_859),
.A2(n_607),
.B1(n_609),
.B2(n_602),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_905),
.B(n_2),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_859),
.A2(n_616),
.B1(n_621),
.B2(n_611),
.Y(n_964)
);

AO22x2_ASAP7_75t_L g965 ( 
.A1(n_865),
.A2(n_627),
.B1(n_523),
.B2(n_596),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_835),
.B(n_750),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_915),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_895),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_922),
.B(n_2),
.Y(n_969)
);

OAI22xp33_ASAP7_75t_SL g970 ( 
.A1(n_833),
.A2(n_520),
.B1(n_518),
.B2(n_510),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_848),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_857),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_920),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_850),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_886),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_862),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_851),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_903),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_922),
.B(n_3),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_894),
.B(n_618),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_SL g981 ( 
.A1(n_910),
.A2(n_461),
.B1(n_463),
.B2(n_460),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_836),
.A2(n_466),
.B1(n_467),
.B2(n_464),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_877),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_925),
.A2(n_470),
.B1(n_476),
.B2(n_468),
.Y(n_984)
);

BUFx8_ASAP7_75t_L g985 ( 
.A(n_870),
.Y(n_985)
);

AO22x2_ASAP7_75t_L g986 ( 
.A1(n_865),
.A2(n_628),
.B1(n_5),
.B2(n_3),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_860),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_852),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_889),
.B(n_896),
.Y(n_989)
);

OAI221xp5_ASAP7_75t_L g990 ( 
.A1(n_869),
.A2(n_494),
.B1(n_495),
.B2(n_493),
.C(n_488),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_870),
.B(n_499),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_853),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_860),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_861),
.B(n_750),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_839),
.B(n_508),
.C(n_507),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_855),
.Y(n_996)
);

INVx3_ASAP7_75t_R g997 ( 
.A(n_906),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_884),
.Y(n_998)
);

BUFx8_ASAP7_75t_L g999 ( 
.A(n_887),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_884),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_858),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_911),
.A2(n_512),
.B1(n_522),
.B2(n_521),
.C(n_515),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_879),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_890),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_891),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_873),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_893),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_864),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_898),
.B(n_722),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_909),
.Y(n_1010)
);

AO22x2_ASAP7_75t_L g1011 ( 
.A1(n_876),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_909),
.Y(n_1012)
);

CKINVDCx14_ASAP7_75t_R g1013 ( 
.A(n_899),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_840),
.B(n_536),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_919),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_898),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_863),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_875),
.Y(n_1018)
);

AO22x2_ASAP7_75t_L g1019 ( 
.A1(n_885),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_899),
.B(n_8),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_868),
.A2(n_540),
.B1(n_541),
.B2(n_537),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_892),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_868),
.A2(n_547),
.B1(n_548),
.B2(n_544),
.Y(n_1023)
);

AOI211xp5_ASAP7_75t_L g1024 ( 
.A1(n_923),
.A2(n_554),
.B(n_555),
.C(n_552),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_863),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_863),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_885),
.B(n_9),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_866),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_863),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_888),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_888),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_875),
.Y(n_1032)
);

AO22x2_ASAP7_75t_L g1033 ( 
.A1(n_871),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_924),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_SL g1035 ( 
.A(n_875),
.B(n_561),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_904),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_904),
.Y(n_1037)
);

BUFx8_ASAP7_75t_L g1038 ( 
.A(n_918),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_918),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_918),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_880),
.Y(n_1041)
);

NAND3x1_ASAP7_75t_L g1042 ( 
.A(n_880),
.B(n_11),
.C(n_14),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_880),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_880),
.A2(n_579),
.B1(n_581),
.B2(n_575),
.Y(n_1044)
);

OAI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_854),
.A2(n_582),
.B1(n_590),
.B2(n_589),
.C(n_586),
.Y(n_1045)
);

NAND3x1_ASAP7_75t_L g1046 ( 
.A(n_854),
.B(n_14),
.C(n_15),
.Y(n_1046)
);

OAI221xp5_ASAP7_75t_L g1047 ( 
.A1(n_854),
.A2(n_597),
.B1(n_612),
.B2(n_608),
.C(n_606),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_841),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_838),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_907),
.B(n_726),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_849),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_838),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_854),
.A2(n_614),
.B1(n_615),
.B2(n_613),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_838),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_854),
.B(n_15),
.Y(n_1055)
);

NAND2x1p5_ASAP7_75t_L g1056 ( 
.A(n_907),
.B(n_733),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_907),
.B(n_16),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_841),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_849),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_905),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_841),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_838),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_841),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_838),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_832),
.Y(n_1065)
);

INVx8_ASAP7_75t_L g1066 ( 
.A(n_905),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_907),
.B(n_726),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_854),
.B(n_516),
.Y(n_1068)
);

AO22x2_ASAP7_75t_L g1069 ( 
.A1(n_834),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_854),
.B(n_516),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_849),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_872),
.B(n_18),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_841),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_907),
.B(n_726),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_872),
.B(n_19),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_907),
.B(n_20),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_907),
.B(n_726),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_917),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_832),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_854),
.B(n_516),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_872),
.B(n_21),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_832),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_975),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_932),
.B(n_21),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1060),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_943),
.B(n_22),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_953),
.B(n_23),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_927),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_1068),
.A2(n_723),
.B(n_26),
.C(n_24),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_991),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_978),
.B(n_25),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_989),
.B(n_25),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_941),
.B(n_26),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1072),
.A2(n_1081),
.B(n_1075),
.C(n_1014),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_948),
.B(n_27),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_988),
.B(n_28),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1060),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_SL g1098 ( 
.A(n_1055),
.B(n_28),
.C(n_29),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1070),
.A2(n_733),
.B(n_732),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_931),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_981),
.B(n_30),
.C(n_31),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_944),
.A2(n_733),
.B(n_583),
.C(n_32),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_935),
.A2(n_723),
.B1(n_32),
.B2(n_30),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_990),
.A2(n_31),
.B(n_33),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_928),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1080),
.A2(n_194),
.B(n_192),
.Y(n_1106)
);

BUFx4f_ASAP7_75t_L g1107 ( 
.A(n_1066),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_958),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_958),
.B(n_196),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1032),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_939),
.A2(n_949),
.B1(n_957),
.B2(n_945),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1022),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_959),
.B(n_33),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1049),
.B(n_34),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1052),
.B(n_34),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1048),
.B(n_36),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1018),
.Y(n_1117)
);

NAND2x1p5_ASAP7_75t_L g1118 ( 
.A(n_1078),
.B(n_199),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1054),
.B(n_37),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1062),
.B(n_37),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1064),
.B(n_38),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1010),
.A2(n_205),
.B(n_203),
.Y(n_1122)
);

AO22x1_ASAP7_75t_L g1123 ( 
.A1(n_985),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_971),
.B(n_39),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1012),
.A2(n_207),
.B(n_206),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_943),
.B(n_41),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_L g1127 ( 
.A(n_1071),
.B(n_583),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1015),
.A2(n_212),
.B(n_211),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1003),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1004),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_926),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_968),
.A2(n_583),
.B1(n_44),
.B2(n_42),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_974),
.B(n_43),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_972),
.B(n_1058),
.Y(n_1134)
);

AO21x1_ASAP7_75t_L g1135 ( 
.A1(n_962),
.A2(n_583),
.B(n_217),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_960),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_977),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_985),
.Y(n_1138)
);

OAI321xp33_ASAP7_75t_L g1139 ( 
.A1(n_1027),
.A2(n_49),
.A3(n_51),
.B1(n_47),
.B2(n_48),
.C(n_50),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1005),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1035),
.A2(n_222),
.B(n_221),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1066),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_937),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1017),
.A2(n_229),
.B(n_226),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_992),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1051),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_987),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_996),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_950),
.B(n_49),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1061),
.B(n_50),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_1045),
.B(n_52),
.C(n_53),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1063),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_942),
.B(n_52),
.C(n_54),
.Y(n_1153)
);

INVxp33_ASAP7_75t_SL g1154 ( 
.A(n_1059),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_964),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_954),
.B(n_56),
.Y(n_1156)
);

NOR2x1p5_ASAP7_75t_SL g1157 ( 
.A(n_1026),
.B(n_232),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1038),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1037),
.A2(n_236),
.B(n_234),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1034),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1073),
.A2(n_62),
.B1(n_58),
.B2(n_60),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1001),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_SL g1163 ( 
.A(n_983),
.B(n_62),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_997),
.B(n_63),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1036),
.A2(n_240),
.B(n_239),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_972),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1039),
.A2(n_242),
.B(n_241),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1000),
.B(n_63),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1040),
.A2(n_248),
.B(n_247),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1007),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_936),
.B(n_64),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_929),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_938),
.B(n_999),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1008),
.A2(n_65),
.B(n_67),
.Y(n_1175)
);

AOI33xp33_ASAP7_75t_L g1176 ( 
.A1(n_1021),
.A2(n_68),
.A3(n_69),
.B1(n_71),
.B2(n_72),
.B3(n_73),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1028),
.A2(n_938),
.B1(n_986),
.B2(n_998),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1029),
.A2(n_252),
.B(n_251),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_L g1179 ( 
.A(n_995),
.B(n_68),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_954),
.B(n_69),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1047),
.A2(n_76),
.B(n_71),
.C(n_74),
.Y(n_1181)
);

NOR2x1p5_ASAP7_75t_L g1182 ( 
.A(n_930),
.B(n_74),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_951),
.B(n_77),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1025),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1002),
.B(n_77),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1041),
.A2(n_257),
.B(n_256),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_993),
.B(n_78),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1030),
.A2(n_260),
.B(n_259),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1024),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_SL g1190 ( 
.A1(n_1016),
.A2(n_82),
.B(n_79),
.C(n_81),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_994),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1031),
.A2(n_967),
.B(n_961),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_951),
.B(n_82),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_973),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1065),
.A2(n_1082),
.B(n_1079),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_986),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1038),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_929),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1006),
.A2(n_266),
.B(n_265),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_960),
.B(n_86),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_947),
.B(n_86),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_976),
.A2(n_274),
.B(n_270),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_979),
.B(n_87),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1009),
.A2(n_276),
.B(n_275),
.Y(n_1204)
);

NOR2x1_ASAP7_75t_L g1205 ( 
.A(n_934),
.B(n_277),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1053),
.B(n_88),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1057),
.B(n_88),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_933),
.A2(n_89),
.B(n_90),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_947),
.B(n_90),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1057),
.B(n_91),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_966),
.B(n_91),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1076),
.B(n_92),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1076),
.B(n_92),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1013),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_966),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_955),
.B(n_93),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_1023),
.B(n_93),
.C(n_95),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_946),
.B(n_95),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_SL g1219 ( 
.A(n_982),
.B(n_96),
.C(n_97),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_956),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_994),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_940),
.B(n_96),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_952),
.B(n_99),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_980),
.B(n_100),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_963),
.B(n_100),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1020),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_969),
.B(n_101),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_980),
.B(n_102),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_965),
.B(n_103),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_980),
.B(n_104),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_970),
.A2(n_286),
.B(n_282),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1044),
.B(n_104),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1046),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1011),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_L g1235 ( 
.A(n_1042),
.B(n_1050),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_965),
.B(n_106),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1011),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1056),
.B(n_107),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1067),
.Y(n_1239)
);

AND2x2_ASAP7_75t_SL g1240 ( 
.A(n_1043),
.B(n_1019),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1019),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1069),
.A2(n_1033),
.B1(n_1077),
.B2(n_1074),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1033),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1069),
.A2(n_290),
.B(n_289),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1166),
.B(n_108),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_292),
.B(n_291),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1218),
.B(n_109),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1105),
.B(n_110),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1088),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1152),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1166),
.B(n_111),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1100),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1107),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1094),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1085),
.B(n_113),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1093),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1209),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1166),
.B(n_118),
.Y(n_1258)
);

NOR3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1146),
.B(n_1098),
.C(n_1084),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1211),
.B(n_118),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1140),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1206),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1262)
);

CKINVDCx14_ASAP7_75t_R g1263 ( 
.A(n_1107),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1154),
.B(n_119),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1145),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1215),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1184),
.B(n_120),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1138),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1148),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1185),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1097),
.B(n_122),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1095),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1090),
.B(n_125),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1184),
.B(n_126),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1162),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1129),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1234),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1277)
);

OR2x6_ASAP7_75t_L g1278 ( 
.A(n_1197),
.B(n_128),
.Y(n_1278)
);

INVx3_ASAP7_75t_SL g1279 ( 
.A(n_1158),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1090),
.B(n_1086),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1112),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1130),
.B(n_129),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1108),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1147),
.B(n_131),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1211),
.B(n_131),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1083),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1111),
.B(n_132),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1214),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1131),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1086),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1126),
.B(n_132),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1126),
.B(n_133),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1171),
.B(n_133),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1092),
.A2(n_134),
.B(n_135),
.C(n_136),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1215),
.B(n_134),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1216),
.B(n_135),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1191),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1225),
.B(n_137),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1208),
.A2(n_138),
.B(n_140),
.C(n_141),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1110),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1240),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1173),
.Y(n_1302)
);

NOR3xp33_ASAP7_75t_SL g1303 ( 
.A(n_1223),
.B(n_142),
.C(n_144),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1243),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1177),
.B(n_145),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_SL g1306 ( 
.A1(n_1181),
.A2(n_146),
.B(n_147),
.C(n_148),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1241),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_1307)
);

AOI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1149),
.A2(n_149),
.B(n_150),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1087),
.B(n_151),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_L g1310 ( 
.A(n_1101),
.B(n_151),
.C(n_152),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1242),
.B(n_152),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1174),
.B(n_153),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1179),
.A2(n_1189),
.B(n_1170),
.C(n_1151),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_R g1314 ( 
.A(n_1158),
.B(n_1142),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1155),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1196),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1116),
.B(n_157),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1150),
.B(n_157),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1178),
.A2(n_306),
.B(n_304),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1132),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1143),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1217),
.B(n_158),
.C(n_159),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1104),
.A2(n_160),
.B(n_161),
.C(n_162),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1183),
.B(n_162),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1203),
.B(n_163),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1194),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1113),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1122),
.A2(n_312),
.B(n_310),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1114),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1115),
.Y(n_1330)
);

CKINVDCx8_ASAP7_75t_R g1331 ( 
.A(n_1198),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1136),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1229),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1187),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1119),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1193),
.B(n_166),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1120),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1237),
.B(n_167),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1168),
.B(n_168),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1121),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1191),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1244),
.A2(n_1180),
.B1(n_1156),
.B2(n_1200),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1226),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1233),
.A2(n_1176),
.B(n_1175),
.C(n_1102),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1221),
.B(n_1118),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1221),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1124),
.B(n_170),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1168),
.B(n_171),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1231),
.A2(n_172),
.B(n_173),
.C(n_174),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1207),
.B(n_175),
.Y(n_1350)
);

O2A1O1Ixp5_ASAP7_75t_L g1351 ( 
.A1(n_1135),
.A2(n_175),
.B(n_176),
.C(n_177),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1133),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1210),
.B(n_176),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1110),
.B(n_177),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1201),
.B(n_178),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1125),
.A2(n_316),
.B(n_315),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_R g1357 ( 
.A(n_1110),
.B(n_318),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1220),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1219),
.A2(n_178),
.B(n_179),
.C(n_180),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1128),
.A2(n_382),
.B(n_454),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1212),
.B(n_180),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1096),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1091),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1213),
.Y(n_1364)
);

CKINVDCx8_ASAP7_75t_R g1365 ( 
.A(n_1117),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1134),
.B(n_181),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1232),
.A2(n_182),
.B(n_183),
.C(n_184),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1227),
.B(n_185),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1172),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1222),
.B(n_185),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1236),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1117),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1195),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1172),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1117),
.B(n_320),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1238),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1239),
.B(n_456),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1089),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1153),
.A2(n_186),
.B1(n_187),
.B2(n_190),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1204),
.A2(n_385),
.B(n_447),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1164),
.A2(n_190),
.B1(n_191),
.B2(n_321),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1106),
.A2(n_387),
.B(n_322),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1109),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1186),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1163),
.A2(n_1139),
.B1(n_1230),
.B2(n_1228),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1224),
.B(n_449),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1160),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1182),
.B(n_444),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1144),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1205),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1123),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1192),
.B(n_328),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1137),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1127),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1161),
.A2(n_1103),
.B1(n_1141),
.B2(n_1188),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1190),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1235),
.A2(n_334),
.B(n_336),
.C(n_338),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1157),
.B(n_443),
.Y(n_1398)
);

INVx3_ASAP7_75t_SL g1399 ( 
.A(n_1302),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1268),
.Y(n_1400)
);

BUFx4_ASAP7_75t_SL g1401 ( 
.A(n_1278),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1281),
.B(n_1165),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1372),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1300),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1345),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1365),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1283),
.Y(n_1407)
);

INVx8_ASAP7_75t_L g1408 ( 
.A(n_1300),
.Y(n_1408)
);

BUFx10_ASAP7_75t_L g1409 ( 
.A(n_1264),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1300),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1331),
.Y(n_1411)
);

INVx5_ASAP7_75t_L g1412 ( 
.A(n_1345),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1369),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1279),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1249),
.B(n_1202),
.Y(n_1415)
);

INVx6_ASAP7_75t_SL g1416 ( 
.A(n_1345),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1266),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1250),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1266),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1373),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1253),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1376),
.B(n_1167),
.Y(n_1422)
);

CKINVDCx6p67_ASAP7_75t_R g1423 ( 
.A(n_1278),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1374),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1288),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1290),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1383),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1247),
.B(n_339),
.Y(n_1428)
);

INVx3_ASAP7_75t_SL g1429 ( 
.A(n_1280),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1362),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1358),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1314),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1357),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1354),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1297),
.B(n_1169),
.Y(n_1435)
);

INVx3_ASAP7_75t_SL g1436 ( 
.A(n_1284),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1383),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1341),
.B(n_1159),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1252),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1383),
.Y(n_1440)
);

INVx3_ASAP7_75t_SL g1441 ( 
.A(n_1355),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1384),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1375),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1348),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1260),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1291),
.B(n_340),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_SL g1447 ( 
.A(n_1285),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1396),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1255),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1341),
.Y(n_1450)
);

BUFx12f_ASAP7_75t_L g1451 ( 
.A(n_1391),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1346),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1261),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1265),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1269),
.Y(n_1455)
);

INVx4_ASAP7_75t_L g1456 ( 
.A(n_1346),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1275),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1271),
.Y(n_1458)
);

INVx5_ASAP7_75t_L g1459 ( 
.A(n_1377),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1276),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1295),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1248),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1263),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1329),
.Y(n_1464)
);

BUFx4_ASAP7_75t_SL g1465 ( 
.A(n_1364),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1389),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1325),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1286),
.Y(n_1468)
);

BUFx8_ASAP7_75t_L g1469 ( 
.A(n_1335),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1394),
.Y(n_1470)
);

INVx6_ASAP7_75t_SL g1471 ( 
.A(n_1339),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1289),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1309),
.B(n_341),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1321),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1326),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1330),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1390),
.B(n_1199),
.Y(n_1478)
);

INVx5_ASAP7_75t_L g1479 ( 
.A(n_1389),
.Y(n_1479)
);

BUFx2_ASAP7_75t_R g1480 ( 
.A(n_1311),
.Y(n_1480)
);

BUFx8_ASAP7_75t_L g1481 ( 
.A(n_1337),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1340),
.Y(n_1482)
);

BUFx12f_ASAP7_75t_L g1483 ( 
.A(n_1389),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1282),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1352),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1273),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1338),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1293),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1378),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1398),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1347),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1259),
.B(n_342),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1334),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1366),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1292),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1392),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1303),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1363),
.Y(n_1498)
);

BUFx4_ASAP7_75t_SL g1499 ( 
.A(n_1322),
.Y(n_1499)
);

INVx8_ASAP7_75t_L g1500 ( 
.A(n_1257),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1246),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1287),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1388),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1336),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1312),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1267),
.B(n_343),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1317),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1296),
.B(n_442),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1318),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1351),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1272),
.Y(n_1511)
);

NAND2x2_ASAP7_75t_L g1512 ( 
.A(n_1298),
.B(n_1310),
.Y(n_1512)
);

BUFx12f_ASAP7_75t_L g1513 ( 
.A(n_1368),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1319),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1305),
.B(n_344),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1254),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1344),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1353),
.Y(n_1518)
);

INVx8_ASAP7_75t_L g1519 ( 
.A(n_1245),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1251),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1258),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1274),
.Y(n_1522)
);

BUFx4f_ASAP7_75t_L g1523 ( 
.A(n_1385),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1350),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1361),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1324),
.Y(n_1526)
);

BUFx2_ASAP7_75t_SL g1527 ( 
.A(n_1370),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1333),
.Y(n_1528)
);

NAND2x1p5_ASAP7_75t_L g1529 ( 
.A(n_1386),
.B(n_345),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1262),
.Y(n_1530)
);

INVx5_ASAP7_75t_L g1531 ( 
.A(n_1397),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1270),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1367),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1256),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1379),
.Y(n_1535)
);

INVx3_ASAP7_75t_SL g1536 ( 
.A(n_1342),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1313),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1332),
.Y(n_1538)
);

CKINVDCx11_ASAP7_75t_R g1539 ( 
.A(n_1307),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1294),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1528),
.A2(n_1316),
.B1(n_1320),
.B2(n_1308),
.C(n_1343),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1526),
.B(n_1277),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1420),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1420),
.Y(n_1544)
);

INVx5_ASAP7_75t_L g1545 ( 
.A(n_1459),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1425),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1439),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1483),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1454),
.B(n_1301),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1530),
.A2(n_1299),
.B1(n_1371),
.B2(n_1381),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1403),
.B(n_1359),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1523),
.A2(n_1323),
.B(n_1349),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1430),
.B(n_1304),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1493),
.B(n_1306),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1439),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1414),
.Y(n_1556)
);

AOI221x1_ASAP7_75t_L g1557 ( 
.A1(n_1532),
.A2(n_1537),
.B1(n_1516),
.B2(n_1533),
.C(n_1515),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1536),
.A2(n_1395),
.B1(n_1393),
.B2(n_1387),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1444),
.B(n_1315),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1407),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1418),
.A2(n_1360),
.B(n_1356),
.C(n_1328),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1534),
.A2(n_1380),
.B1(n_1382),
.B2(n_349),
.C(n_350),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1514),
.A2(n_347),
.B(n_348),
.Y(n_1563)
);

OAI211xp5_ASAP7_75t_L g1564 ( 
.A1(n_1539),
.A2(n_1511),
.B(n_1517),
.C(n_1500),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1445),
.B(n_351),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1514),
.A2(n_352),
.B(n_353),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1507),
.B(n_356),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1478),
.A2(n_357),
.B(n_358),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_L g1569 ( 
.A(n_1517),
.B(n_359),
.C(n_361),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1426),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1457),
.B(n_362),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_SL g1572 ( 
.A1(n_1402),
.A2(n_364),
.B(n_365),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1405),
.B(n_366),
.Y(n_1573)
);

INVx3_ASAP7_75t_SL g1574 ( 
.A(n_1399),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1509),
.B(n_367),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1490),
.A2(n_441),
.B(n_369),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1531),
.A2(n_368),
.B(n_371),
.Y(n_1577)
);

NAND2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1459),
.B(n_373),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1435),
.A2(n_375),
.B(n_376),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1502),
.B(n_377),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_SL g1581 ( 
.A1(n_1502),
.A2(n_379),
.B(n_380),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1501),
.A2(n_440),
.B(n_383),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1453),
.B(n_1455),
.Y(n_1583)
);

AO31x2_ASAP7_75t_L g1584 ( 
.A1(n_1496),
.A2(n_381),
.A3(n_388),
.B(n_389),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1438),
.A2(n_390),
.B(n_391),
.Y(n_1585)
);

AOI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1496),
.A2(n_392),
.B(n_393),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1463),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1455),
.B(n_394),
.Y(n_1588)
);

NAND2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1459),
.B(n_1406),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1405),
.B(n_396),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1442),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1489),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1463),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1498),
.B(n_397),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1500),
.A2(n_398),
.B1(n_400),
.B2(n_401),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1473),
.A2(n_402),
.B(n_403),
.C(n_404),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1531),
.A2(n_1516),
.B(n_1508),
.C(n_1494),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1498),
.B(n_406),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1540),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1512),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.C(n_413),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1441),
.B(n_415),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1450),
.Y(n_1602)
);

AOI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1535),
.A2(n_416),
.B(n_417),
.Y(n_1603)
);

OAI21xp33_ASAP7_75t_L g1604 ( 
.A1(n_1538),
.A2(n_421),
.B(n_422),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1412),
.B(n_423),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1442),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1412),
.B(n_1443),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1415),
.A2(n_425),
.B(n_426),
.Y(n_1608)
);

A2O1A1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1531),
.A2(n_427),
.B(n_429),
.C(n_431),
.Y(n_1609)
);

NOR2xp67_ASAP7_75t_L g1610 ( 
.A(n_1479),
.B(n_432),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1466),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1400),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1487),
.B(n_433),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1469),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1460),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1456),
.Y(n_1616)
);

NAND2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1412),
.B(n_434),
.Y(n_1617)
);

AO21x2_ASAP7_75t_L g1618 ( 
.A1(n_1422),
.A2(n_439),
.B(n_436),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1433),
.B(n_1411),
.Y(n_1619)
);

BUFx4f_ASAP7_75t_L g1620 ( 
.A(n_1451),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1417),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1547),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1611),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1545),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1547),
.B(n_1466),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1545),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1555),
.Y(n_1627)
);

INVx11_ASAP7_75t_L g1628 ( 
.A(n_1546),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1543),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1543),
.Y(n_1630)
);

AO21x2_ASAP7_75t_L g1631 ( 
.A1(n_1597),
.A2(n_1487),
.B(n_1474),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1544),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1552),
.A2(n_1513),
.B1(n_1525),
.B2(n_1524),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1550),
.A2(n_1486),
.B1(n_1436),
.B2(n_1458),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1614),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1541),
.A2(n_1449),
.B1(n_1475),
.B2(n_1476),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1570),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1591),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1542),
.A2(n_1475),
.B1(n_1476),
.B2(n_1431),
.Y(n_1639)
);

BUFx8_ASAP7_75t_L g1640 ( 
.A(n_1564),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1557),
.A2(n_1510),
.B(n_1448),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1583),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1558),
.A2(n_1484),
.B1(n_1468),
.B2(n_1472),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1591),
.Y(n_1644)
);

INVx6_ASAP7_75t_L g1645 ( 
.A(n_1587),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1600),
.A2(n_1447),
.B1(n_1480),
.B2(n_1505),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1606),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1615),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1582),
.B(n_1482),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1582),
.B(n_1479),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1592),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1553),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1584),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1592),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1559),
.B(n_1477),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1574),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1598),
.Y(n_1657)
);

NAND2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_1479),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1549),
.B(n_1485),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1580),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1578),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1571),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1637),
.B(n_1477),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1625),
.B(n_1560),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1628),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1628),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1656),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1638),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1629),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1493),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1647),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1651),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1630),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_SL g1674 ( 
.A(n_1646),
.B(n_1551),
.C(n_1462),
.Y(n_1674)
);

BUFx2_ASAP7_75t_SL g1675 ( 
.A(n_1654),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1634),
.A2(n_1554),
.B1(n_1595),
.B2(n_1505),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1632),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1632),
.Y(n_1678)
);

OAI222xp33_ASAP7_75t_L g1679 ( 
.A1(n_1652),
.A2(n_1464),
.B1(n_1467),
.B2(n_1488),
.C1(n_1588),
.C2(n_1491),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1635),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1641),
.A2(n_1596),
.B(n_1609),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1623),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_R g1683 ( 
.A(n_1635),
.B(n_1448),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1645),
.B(n_1556),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1640),
.Y(n_1685)
);

CKINVDCx16_ASAP7_75t_R g1686 ( 
.A(n_1659),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1645),
.Y(n_1687)
);

NOR2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1655),
.B(n_1423),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1623),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1650),
.B(n_1589),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1687),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1669),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1686),
.B(n_1642),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1690),
.B(n_1650),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1664),
.B(n_1625),
.Y(n_1696)
);

NOR2x1p5_ASAP7_75t_L g1697 ( 
.A(n_1685),
.B(n_1612),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1668),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1689),
.B(n_1659),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1674),
.A2(n_1527),
.B1(n_1649),
.B2(n_1471),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1689),
.B(n_1644),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1673),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1671),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1681),
.A2(n_1649),
.B1(n_1471),
.B2(n_1631),
.Y(n_1704)
);

OR2x6_ASAP7_75t_SL g1705 ( 
.A(n_1685),
.B(n_1660),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1673),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1699),
.B(n_1663),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1698),
.B(n_1677),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1703),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1693),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1705),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1692),
.A2(n_1641),
.B(n_1678),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1701),
.Y(n_1713)
);

AO21x1_ASAP7_75t_SL g1714 ( 
.A1(n_1700),
.A2(n_1627),
.B(n_1622),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1711),
.B(n_1705),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1709),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1708),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1708),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1707),
.B(n_1672),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1710),
.B(n_1691),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1713),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1720),
.B(n_1667),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1719),
.B(n_1694),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1716),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1718),
.B(n_1587),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1716),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1718),
.B(n_1717),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1715),
.B(n_1667),
.Y(n_1728)
);

NAND2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1715),
.B(n_1620),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1696),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1726),
.B(n_1702),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1728),
.B(n_1680),
.Y(n_1732)
);

INVxp33_ASAP7_75t_L g1733 ( 
.A(n_1722),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1726),
.B(n_1702),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1724),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1729),
.B(n_1697),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1721),
.B(n_1680),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1727),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1723),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1730),
.B(n_1665),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1725),
.B(n_1712),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1737),
.B(n_1665),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1732),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_R g1744 ( 
.A(n_1737),
.B(n_1666),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1739),
.B(n_1725),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1733),
.B(n_1666),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1736),
.B(n_1670),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1738),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1735),
.Y(n_1749)
);

OAI21xp33_ASAP7_75t_L g1750 ( 
.A1(n_1743),
.A2(n_1734),
.B(n_1731),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1748),
.B(n_1740),
.Y(n_1751)
);

NAND2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1746),
.B(n_1620),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1749),
.Y(n_1753)
);

O2A1O1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1745),
.B(n_1741),
.C(n_1747),
.Y(n_1754)
);

AOI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1751),
.A2(n_1745),
.B(n_1744),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1750),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1752),
.A2(n_1712),
.B1(n_1742),
.B2(n_1676),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1756),
.B(n_1664),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1755),
.B(n_1409),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1754),
.B(n_1757),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1756),
.B(n_1633),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1756),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1762),
.B(n_1432),
.C(n_1601),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1759),
.B(n_1758),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1761),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1760),
.B(n_1413),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1758),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1758),
.Y(n_1768)
);

XOR2xp5_ASAP7_75t_L g1769 ( 
.A(n_1761),
.B(n_1587),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1758),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1758),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1688),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1765),
.A2(n_1704),
.B1(n_1503),
.B2(n_1481),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1497),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1768),
.B(n_1770),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1771),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1769),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1766),
.A2(n_1492),
.B(n_1594),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1764),
.B(n_1481),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1772),
.B(n_1675),
.Y(n_1780)
);

AOI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1763),
.A2(n_1401),
.B(n_1492),
.C(n_1593),
.Y(n_1781)
);

NAND5xp2_ASAP7_75t_L g1782 ( 
.A(n_1766),
.B(n_1619),
.C(n_1700),
.D(n_1704),
.E(n_1446),
.Y(n_1782)
);

AO21x1_ASAP7_75t_L g1783 ( 
.A1(n_1766),
.A2(n_1683),
.B(n_1506),
.Y(n_1783)
);

OAI21xp33_ASAP7_75t_L g1784 ( 
.A1(n_1766),
.A2(n_1684),
.B(n_1548),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1779),
.A2(n_1775),
.B(n_1776),
.Y(n_1785)
);

AOI221x1_ASAP7_75t_L g1786 ( 
.A1(n_1777),
.A2(n_1593),
.B1(n_1613),
.B2(n_1506),
.C(n_1421),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1774),
.A2(n_1593),
.B(n_1519),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1781),
.B(n_1640),
.C(n_1428),
.Y(n_1788)
);

AOI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1783),
.A2(n_1567),
.B(n_1575),
.C(n_1565),
.Y(n_1789)
);

AOI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1780),
.A2(n_1424),
.B(n_1504),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1784),
.B(n_1640),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1778),
.Y(n_1792)
);

AO221x1_ASAP7_75t_L g1793 ( 
.A1(n_1782),
.A2(n_1548),
.B1(n_1421),
.B2(n_1465),
.C(n_1522),
.Y(n_1793)
);

OAI31xp33_ASAP7_75t_L g1794 ( 
.A1(n_1773),
.A2(n_1604),
.A3(n_1617),
.B(n_1529),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1775),
.A2(n_1695),
.B1(n_1636),
.B2(n_1562),
.C(n_1518),
.Y(n_1795)
);

NOR3xp33_ASAP7_75t_L g1796 ( 
.A(n_1777),
.B(n_1569),
.C(n_1586),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_L g1797 ( 
.A(n_1785),
.B(n_1469),
.C(n_1599),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1788),
.A2(n_1503),
.B1(n_1495),
.B2(n_1519),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1792),
.Y(n_1799)
);

OAI221xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1791),
.A2(n_1695),
.B1(n_1577),
.B2(n_1434),
.C(n_1521),
.Y(n_1800)
);

AOI22x1_ASAP7_75t_L g1801 ( 
.A1(n_1787),
.A2(n_1706),
.B1(n_1602),
.B2(n_1616),
.Y(n_1801)
);

AO21x1_ASAP7_75t_L g1802 ( 
.A1(n_1790),
.A2(n_1590),
.B(n_1573),
.Y(n_1802)
);

NAND4xp25_ASAP7_75t_L g1803 ( 
.A(n_1786),
.B(n_1605),
.C(n_1573),
.D(n_1590),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1796),
.A2(n_1429),
.B1(n_1650),
.B2(n_1645),
.C(n_1610),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1795),
.A2(n_1579),
.B(n_1585),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1793),
.B(n_1706),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1789),
.A2(n_1581),
.B1(n_1572),
.B2(n_1485),
.C(n_1648),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1799),
.B(n_1802),
.Y(n_1808)
);

NOR2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1797),
.B(n_1794),
.Y(n_1809)
);

AOI222xp33_ASAP7_75t_L g1810 ( 
.A1(n_1804),
.A2(n_1461),
.B1(n_1653),
.B2(n_1679),
.C1(n_1520),
.C2(n_1470),
.Y(n_1810)
);

XOR2xp5_ASAP7_75t_L g1811 ( 
.A(n_1798),
.B(n_1605),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1803),
.B(n_1654),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1520),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1805),
.A2(n_1461),
.B1(n_1561),
.B2(n_1603),
.C(n_1618),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1806),
.B(n_1801),
.Y(n_1815)
);

NAND2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1800),
.B(n_1602),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1799),
.B(n_1673),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1799),
.B(n_1687),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1808),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1815),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1818),
.B(n_1662),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1817),
.B(n_1812),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1813),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1816),
.A2(n_1610),
.B1(n_1645),
.B2(n_1563),
.C(n_1695),
.Y(n_1824)
);

INVxp67_ASAP7_75t_SL g1825 ( 
.A(n_1809),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1811),
.Y(n_1826)
);

NAND4xp75_ASAP7_75t_L g1827 ( 
.A(n_1814),
.B(n_1563),
.C(n_1437),
.D(n_1499),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1825),
.Y(n_1828)
);

CKINVDCx16_ASAP7_75t_R g1829 ( 
.A(n_1820),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1819),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1822),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1823),
.B(n_1810),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1826),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1821),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1827),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1828),
.A2(n_1824),
.B(n_1566),
.Y(n_1836)
);

XNOR2x1_ASAP7_75t_L g1837 ( 
.A(n_1831),
.B(n_1427),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1829),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1833),
.Y(n_1839)
);

OA22x2_ASAP7_75t_L g1840 ( 
.A1(n_1830),
.A2(n_1616),
.B1(n_1621),
.B2(n_1568),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1832),
.A2(n_1427),
.B1(n_1440),
.B2(n_1661),
.C(n_1690),
.Y(n_1841)
);

OAI22x1_ASAP7_75t_L g1842 ( 
.A1(n_1835),
.A2(n_1621),
.B1(n_1410),
.B2(n_1658),
.Y(n_1842)
);

CKINVDCx20_ASAP7_75t_R g1843 ( 
.A(n_1838),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1839),
.A2(n_1834),
.B1(n_1440),
.B2(n_1416),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1836),
.B(n_1661),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1837),
.A2(n_1576),
.B1(n_1661),
.B2(n_1452),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1842),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1840),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1847),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1843),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1848),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1844),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1845),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1846),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1850),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1849),
.Y(n_1856)
);

CKINVDCx20_ASAP7_75t_R g1857 ( 
.A(n_1851),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1853),
.B(n_1841),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_SL g1859 ( 
.A1(n_1856),
.A2(n_1852),
.B(n_1854),
.C(n_437),
.Y(n_1859)
);

AOI22x1_ASAP7_75t_L g1860 ( 
.A1(n_1855),
.A2(n_1857),
.B1(n_1858),
.B2(n_1452),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1855),
.A2(n_1416),
.B1(n_1661),
.B2(n_1404),
.Y(n_1861)
);

NAND4xp25_ASAP7_75t_SL g1862 ( 
.A(n_1860),
.B(n_1639),
.C(n_1643),
.D(n_1714),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1859),
.A2(n_1404),
.B1(n_1661),
.B2(n_1419),
.C(n_1417),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_1863),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1864),
.A2(n_1861),
.B1(n_1862),
.B2(n_1408),
.Y(n_1865)
);

OR2x6_ASAP7_75t_L g1866 ( 
.A(n_1865),
.B(n_1408),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1866),
.A2(n_438),
.B(n_1608),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1419),
.B(n_1624),
.C(n_1626),
.Y(n_1868)
);


endmodule