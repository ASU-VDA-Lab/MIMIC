module fake_aes_12630_n_479 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_479);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_479;
wire n_117;
wire n_361;
wire n_185;
wire n_57;
wire n_407;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_56;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_58;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g56 ( .A(n_11), .Y(n_56) );
INVx1_ASAP7_75t_L g57 ( .A(n_47), .Y(n_57) );
INVx1_ASAP7_75t_L g58 ( .A(n_48), .Y(n_58) );
INVx1_ASAP7_75t_L g59 ( .A(n_27), .Y(n_59) );
INVx1_ASAP7_75t_L g60 ( .A(n_9), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_24), .Y(n_61) );
HB1xp67_ASAP7_75t_L g62 ( .A(n_11), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_23), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_15), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_19), .Y(n_65) );
BUFx6f_ASAP7_75t_L g66 ( .A(n_19), .Y(n_66) );
CKINVDCx5p33_ASAP7_75t_R g67 ( .A(n_1), .Y(n_67) );
INVx1_ASAP7_75t_SL g68 ( .A(n_35), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_53), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_51), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_5), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_33), .Y(n_72) );
INVxp67_ASAP7_75t_L g73 ( .A(n_28), .Y(n_73) );
INVxp33_ASAP7_75t_L g74 ( .A(n_14), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_21), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_36), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_17), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_4), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_32), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_54), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_29), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_45), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_40), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_49), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_50), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_44), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_39), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_22), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_52), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVx4_ASAP7_75t_R g92 ( .A(n_25), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_0), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_8), .Y(n_94) );
INVx1_ASAP7_75t_SL g95 ( .A(n_15), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_57), .Y(n_96) );
NOR2xp33_ASAP7_75t_L g97 ( .A(n_74), .B(n_0), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_89), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_57), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_71), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_56), .B(n_1), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_59), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_59), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_62), .B(n_2), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_86), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_56), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_84), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_87), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_63), .B(n_2), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_77), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_63), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_94), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_73), .B(n_3), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_68), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_69), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_60), .B(n_3), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_95), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_69), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_70), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_70), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_76), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_96), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_104), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_96), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_104), .B(n_88), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_96), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_105), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_105), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
INVx2_ASAP7_75t_SL g137 ( .A(n_100), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_123), .Y(n_138) );
AOI22xp33_ASAP7_75t_SL g139 ( .A1(n_121), .A2(n_60), .B1(n_64), .B2(n_65), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_100), .B(n_80), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g144 ( .A(n_102), .B(n_83), .C(n_79), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_124), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_104), .B(n_72), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_126), .B(n_83), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
NAND3x1_ASAP7_75t_L g151 ( .A(n_121), .B(n_80), .C(n_91), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_103), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_109), .B(n_64), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_103), .B(n_91), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_106), .B(n_90), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_127), .Y(n_158) );
NAND2x1p5_ASAP7_75t_L g159 ( .A(n_121), .B(n_79), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_127), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_106), .B(n_90), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_111), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_111), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_109), .B(n_65), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
OR2x2_ASAP7_75t_L g167 ( .A(n_142), .B(n_117), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_131), .A2(n_108), .B1(n_99), .B2(n_101), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_165), .B(n_153), .Y(n_170) );
OR2x6_ASAP7_75t_L g171 ( .A(n_159), .B(n_107), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
O2A1O1Ixp5_ASAP7_75t_L g173 ( .A1(n_132), .A2(n_114), .B(n_118), .C(n_112), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_165), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_149), .B(n_113), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_159), .B(n_107), .Y(n_176) );
XNOR2xp5_ASAP7_75t_L g177 ( .A(n_151), .B(n_115), .Y(n_177) );
NAND2xp33_ASAP7_75t_R g178 ( .A(n_165), .B(n_98), .Y(n_178) );
HB1xp67_ASAP7_75t_SL g179 ( .A(n_131), .Y(n_179) );
AND3x1_ASAP7_75t_SL g180 ( .A(n_139), .B(n_75), .C(n_78), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_153), .A2(n_125), .B(n_120), .C(n_116), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_163), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_131), .A2(n_125), .B1(n_116), .B2(n_120), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_149), .B(n_110), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_149), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_152), .B(n_119), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_131), .B(n_118), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_165), .B(n_97), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_146), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g197 ( .A(n_144), .B(n_97), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_165), .B(n_114), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_150), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_129), .A2(n_85), .B1(n_66), .B2(n_93), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_148), .B(n_122), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_159), .B(n_81), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_137), .B(n_66), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_148), .B(n_82), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_153), .B(n_85), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_129), .A2(n_66), .B1(n_88), .B2(n_92), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_196), .B(n_137), .Y(n_210) );
AND3x1_ASAP7_75t_SL g211 ( .A(n_177), .B(n_151), .C(n_139), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_186), .A2(n_199), .B(n_194), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_176), .B(n_151), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_176), .B(n_137), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_166), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_181), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_181), .Y(n_219) );
INVx5_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
OAI221xp5_ASAP7_75t_L g221 ( .A1(n_195), .A2(n_146), .B1(n_156), .B2(n_141), .C(n_162), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_196), .B(n_132), .Y(n_223) );
CKINVDCx11_ASAP7_75t_R g224 ( .A(n_187), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_170), .B(n_168), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_191), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_170), .B(n_129), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_181), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_179), .A2(n_146), .B1(n_147), .B2(n_162), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_174), .B(n_147), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_172), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_184), .A2(n_146), .B1(n_147), .B2(n_163), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_202), .B(n_141), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_167), .B(n_156), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_208), .B(n_164), .Y(n_239) );
NAND2x1p5_ASAP7_75t_L g240 ( .A(n_188), .B(n_164), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_208), .B(n_155), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_186), .A2(n_155), .B(n_161), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_167), .A2(n_164), .B1(n_163), .B2(n_144), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_183), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_178), .A2(n_161), .B1(n_143), .B2(n_158), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_240), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_227), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_224), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_237), .A2(n_208), .B1(n_197), .B2(n_203), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_238), .A2(n_169), .B1(n_203), .B2(n_189), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_216), .B(n_169), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_224), .Y(n_254) );
OAI222xp33_ASAP7_75t_L g255 ( .A1(n_212), .A2(n_177), .B1(n_180), .B2(n_189), .C1(n_182), .C2(n_204), .Y(n_255) );
NAND2x1_ASAP7_75t_L g256 ( .A(n_230), .B(n_191), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_220), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g258 ( .A1(n_220), .A2(n_175), .B1(n_136), .B2(n_135), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_234), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_227), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_221), .A2(n_173), .B(n_190), .Y(n_261) );
NOR3xp33_ASAP7_75t_L g262 ( .A(n_226), .B(n_193), .C(n_207), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_230), .B(n_188), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_213), .A2(n_200), .B(n_190), .Y(n_264) );
BUFx2_ASAP7_75t_R g265 ( .A(n_225), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_225), .B(n_201), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_244), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_227), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_220), .A2(n_154), .B1(n_133), .B2(n_134), .Y(n_269) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_264), .A2(n_242), .B(n_244), .Y(n_270) );
AOI33xp33_ASAP7_75t_L g271 ( .A1(n_250), .A2(n_243), .A3(n_241), .B1(n_209), .B2(n_211), .B3(n_158), .Y(n_271) );
BUFx2_ASAP7_75t_SL g272 ( .A(n_246), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_264), .A2(n_232), .B(n_200), .Y(n_273) );
OAI211xp5_ASAP7_75t_L g274 ( .A1(n_250), .A2(n_185), .B(n_214), .C(n_245), .Y(n_274) );
AO31x2_ASAP7_75t_L g275 ( .A1(n_261), .A2(n_235), .A3(n_140), .B(n_145), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_262), .A2(n_218), .B1(n_212), .B2(n_222), .Y(n_276) );
AOI222xp33_ASAP7_75t_L g277 ( .A1(n_255), .A2(n_231), .B1(n_218), .B2(n_241), .C1(n_212), .C2(n_222), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g278 ( .A1(n_258), .A2(n_222), .B(n_239), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_255), .A2(n_231), .B1(n_241), .B2(n_228), .C(n_215), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_253), .B(n_220), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_253), .B(n_228), .Y(n_281) );
HB1xp67_ASAP7_75t_SL g282 ( .A(n_254), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_262), .A2(n_251), .B1(n_252), .B2(n_259), .C(n_253), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_267), .B(n_228), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_265), .B(n_236), .Y(n_285) );
AOI22xp33_ASAP7_75t_SL g286 ( .A1(n_254), .A2(n_240), .B1(n_236), .B2(n_217), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_251), .A2(n_233), .B1(n_236), .B2(n_217), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_267), .B(n_240), .Y(n_288) );
NAND2x1_ASAP7_75t_L g289 ( .A(n_246), .B(n_227), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_252), .A2(n_136), .B1(n_133), .B2(n_134), .C(n_135), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_247), .B(n_229), .Y(n_291) );
AOI33xp33_ASAP7_75t_L g292 ( .A1(n_283), .A2(n_138), .A3(n_143), .B1(n_154), .B2(n_263), .B3(n_258), .Y(n_292) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_283), .A2(n_265), .B(n_249), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_279), .A2(n_269), .B1(n_266), .B2(n_246), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_287), .A2(n_269), .B1(n_266), .B2(n_246), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_282), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_272), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_288), .B(n_246), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_272), .B(n_247), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_288), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
AOI21x1_ASAP7_75t_L g303 ( .A1(n_273), .A2(n_256), .B(n_264), .Y(n_303) );
NAND2xp33_ASAP7_75t_R g304 ( .A(n_285), .B(n_247), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_281), .A2(n_266), .B1(n_257), .B2(n_263), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_281), .A2(n_263), .B1(n_261), .B2(n_66), .C(n_257), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
OAI321xp33_ASAP7_75t_L g308 ( .A1(n_274), .A2(n_66), .A3(n_257), .B1(n_138), .B2(n_229), .C(n_206), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_277), .B(n_256), .C(n_150), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_280), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_284), .B(n_248), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_291), .B(n_268), .Y(n_315) );
OAI211xp5_ASAP7_75t_SL g316 ( .A1(n_271), .A2(n_140), .B(n_145), .C(n_157), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_275), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_302), .B(n_275), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_311), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_301), .B(n_275), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
OAI31xp33_ASAP7_75t_L g323 ( .A1(n_293), .A2(n_278), .A3(n_276), .B(n_291), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_294), .A2(n_277), .B1(n_278), .B2(n_286), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_318), .B(n_275), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_275), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_311), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_313), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_313), .Y(n_329) );
OAI321xp33_ASAP7_75t_L g330 ( .A1(n_305), .A2(n_295), .A3(n_310), .B1(n_309), .B2(n_299), .C(n_300), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_318), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_314), .B(n_275), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_273), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_306), .A2(n_256), .B1(n_290), .B2(n_233), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_300), .B(n_268), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_299), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_312), .A2(n_260), .B1(n_268), .B2(n_248), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_289), .B(n_260), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_298), .B(n_268), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_317), .B(n_248), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_316), .A2(n_150), .B1(n_160), .B2(n_145), .C(n_157), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_298), .B(n_248), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_312), .B(n_140), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_299), .B(n_157), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_299), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_315), .B(n_160), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_315), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_292), .A2(n_233), .B(n_160), .Y(n_351) );
OAI33xp33_ASAP7_75t_L g352 ( .A1(n_296), .A2(n_4), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_297), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_296), .B(n_6), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_304), .B(n_260), .Y(n_356) );
AND2x4_ASAP7_75t_SL g357 ( .A(n_347), .B(n_260), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_353), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_353), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_7), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_338), .Y(n_361) );
OAI33xp33_ASAP7_75t_L g362 ( .A1(n_354), .A2(n_9), .A3(n_10), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_332), .B(n_10), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_338), .B(n_260), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_328), .B(n_13), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_328), .Y(n_366) );
OAI31xp33_ASAP7_75t_L g367 ( .A1(n_355), .A2(n_217), .A3(n_219), .B(n_210), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_16), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_320), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_354), .B(n_17), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_333), .B(n_18), .Y(n_373) );
OAI33xp33_ASAP7_75t_L g374 ( .A1(n_319), .A2(n_20), .A3(n_223), .B1(n_26), .B2(n_30), .B3(n_31), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_322), .B(n_150), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_333), .B(n_150), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_322), .B(n_345), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_355), .Y(n_378) );
AOI211xp5_ASAP7_75t_L g379 ( .A1(n_330), .A2(n_219), .B(n_192), .C(n_191), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_324), .A2(n_219), .B1(n_227), .B2(n_260), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_333), .B(n_260), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_329), .Y(n_382) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_347), .B(n_260), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_329), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_338), .B(n_34), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_345), .B(n_37), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_319), .B(n_38), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_348), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_321), .B(n_326), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_338), .B(n_41), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_321), .B(n_42), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_327), .B(n_43), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_327), .Y(n_393) );
OR2x6_ASAP7_75t_L g394 ( .A(n_347), .B(n_192), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_379), .A2(n_347), .B1(n_339), .B2(n_334), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_389), .B(n_350), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_389), .B(n_350), .Y(n_397) );
AOI21xp33_ASAP7_75t_SL g398 ( .A1(n_378), .A2(n_323), .B(n_346), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_363), .B(n_326), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_362), .A2(n_352), .B(n_346), .C(n_351), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_369), .B(n_349), .Y(n_401) );
AOI21xp33_ASAP7_75t_SL g402 ( .A1(n_360), .A2(n_346), .B(n_356), .Y(n_402) );
INVxp33_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_350), .B1(n_341), .B2(n_344), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_360), .A2(n_348), .B1(n_325), .B2(n_340), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_388), .B(n_327), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_358), .B(n_344), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_371), .A2(n_343), .B(n_348), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_370), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g413 ( .A1(n_359), .A2(n_325), .A3(n_331), .B1(n_337), .B2(n_335), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_381), .B(n_341), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_368), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_357), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_387), .A2(n_325), .B(n_337), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_367), .A2(n_343), .B1(n_331), .B2(n_340), .C(n_335), .Y(n_419) );
OAI21x1_ASAP7_75t_SL g420 ( .A1(n_361), .A2(n_336), .B(n_342), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_374), .A2(n_342), .B1(n_336), .B2(n_198), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
NAND2x1_ASAP7_75t_L g423 ( .A(n_394), .B(n_385), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_357), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_368), .B(n_342), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_409), .B(n_376), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_396), .B(n_372), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_415), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g429 ( .A1(n_423), .A2(n_385), .B1(n_390), .B2(n_394), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_397), .B(n_407), .Y(n_430) );
NAND2xp33_ASAP7_75t_SL g431 ( .A(n_403), .B(n_391), .Y(n_431) );
NOR4xp25_ASAP7_75t_SL g432 ( .A(n_398), .B(n_394), .C(n_383), .D(n_380), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_408), .B(n_387), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_399), .B(n_393), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_416), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_417), .Y(n_438) );
XOR2x2_ASAP7_75t_L g439 ( .A(n_395), .B(n_386), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_414), .B(n_372), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_412), .B(n_375), .Y(n_441) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_420), .B(n_394), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_401), .B(n_336), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_422), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_434), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g446 ( .A(n_439), .B(n_404), .Y(n_446) );
XOR2xp5_ASAP7_75t_L g447 ( .A(n_439), .B(n_411), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_430), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_436), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_444), .Y(n_450) );
AOI22xp5_ASAP7_75t_SL g451 ( .A1(n_438), .A2(n_424), .B1(n_412), .B2(n_405), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_440), .B(n_402), .Y(n_452) );
NOR2x1_ASAP7_75t_SL g453 ( .A(n_430), .B(n_425), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_437), .A2(n_406), .B1(n_400), .B2(n_413), .C(n_418), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_442), .A2(n_419), .B(n_421), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_433), .A2(n_392), .B(n_342), .Y(n_456) );
XOR2x2_ASAP7_75t_L g457 ( .A(n_429), .B(n_392), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_440), .B(n_364), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_443), .B(n_364), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_427), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_455), .A2(n_431), .B(n_441), .C(n_432), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_451), .A2(n_427), .B1(n_426), .B2(n_435), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_448), .B(n_454), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_452), .B(n_428), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_446), .A2(n_205), .B1(n_191), .B2(n_192), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_457), .A2(n_198), .B1(n_205), .B2(n_55), .Y(n_466) );
OAI211xp5_ASAP7_75t_SL g467 ( .A1(n_445), .A2(n_449), .B(n_460), .C(n_456), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g468 ( .A1(n_457), .A2(n_452), .B1(n_453), .B2(n_459), .C1(n_450), .C2(n_458), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_459), .A2(n_447), .B1(n_446), .B2(n_457), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_458), .A2(n_447), .B1(n_446), .B2(n_457), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_464), .Y(n_471) );
NAND2x1_ASAP7_75t_L g472 ( .A(n_462), .B(n_470), .Y(n_472) );
INVx4_ASAP7_75t_L g473 ( .A(n_471), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_472), .A2(n_469), .B1(n_463), .B2(n_468), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_473), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_474), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_475), .Y(n_477) );
XNOR2x1_ASAP7_75t_L g478 ( .A(n_477), .B(n_476), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_478), .A2(n_461), .B1(n_465), .B2(n_466), .C(n_467), .Y(n_479) );
endmodule