module fake_aes_3688_n_29 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_9), .B(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_0), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_1), .Y(n_18) );
OR2x2_ASAP7_75t_L g19 ( .A(n_13), .B(n_3), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_17), .B(n_18), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_14), .B1(n_19), .B2(n_16), .Y(n_22) );
OAI33xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .A3(n_14), .B1(n_19), .B2(n_15), .B3(n_21), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_0), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_26) );
AOI311xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_2), .A3(n_4), .B(n_5), .C(n_6), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_11), .C1(n_12), .C2(n_14), .Y(n_29) );
endmodule