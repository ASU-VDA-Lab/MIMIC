module fake_jpeg_22177_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_9),
.B1(n_13),
.B2(n_2),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_18),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_58),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_10),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_22),
.C(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_76),
.B1(n_31),
.B2(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_28),
.B1(n_15),
.B2(n_21),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_69),
.B(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_31),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_46),
.B1(n_17),
.B2(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_48),
.B1(n_59),
.B2(n_47),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_38),
.B1(n_37),
.B2(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_43),
.B1(n_56),
.B2(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_36),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_43),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_29),
.B1(n_26),
.B2(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_86),
.B1(n_88),
.B2(n_95),
.Y(n_101)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_78),
.B1(n_35),
.B2(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_89),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_51),
.B1(n_29),
.B2(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_36),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_58),
.B1(n_45),
.B2(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_96),
.B1(n_19),
.B2(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_37),
.B1(n_31),
.B2(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_69),
.B2(n_66),
.Y(n_102)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_52),
.B1(n_35),
.B2(n_32),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_27),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_27),
.B(n_24),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_67),
.C(n_63),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_106),
.C(n_119),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_110),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_116),
.B1(n_117),
.B2(n_105),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_80),
.B(n_71),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_91),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_100),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_76),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_115),
.B(n_81),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_74),
.C(n_64),
.Y(n_115)
);

CKINVDCx10_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_19),
.B1(n_93),
.B2(n_24),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_75),
.C(n_19),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_125),
.B(n_136),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_106),
.B(n_24),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_94),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_88),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_87),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_137),
.B1(n_105),
.B2(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_108),
.B(n_27),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_93),
.C(n_27),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_27),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_27),
.C(n_24),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_0),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_103),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_140),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_24),
.B1(n_9),
.B2(n_2),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_147),
.B1(n_144),
.B2(n_145),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_101),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_9),
.B1(n_13),
.B2(n_4),
.C(n_6),
.Y(n_157)
);

OAI322xp33_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_124),
.A3(n_136),
.B1(n_135),
.B2(n_133),
.C1(n_125),
.C2(n_126),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_157),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_130),
.B1(n_121),
.B2(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_139),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_10),
.B1(n_13),
.B2(n_6),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_0),
.CI(n_1),
.CON(n_163),
.SN(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_142),
.B1(n_152),
.B2(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_175),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_174),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_138),
.C(n_1),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_161),
.Y(n_175)
);

NAND4xp25_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_160),
.C(n_156),
.D(n_163),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_183),
.B(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_163),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_181),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_164),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_164),
.B(n_162),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_184),
.B(n_186),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_183),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_168),
.B(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_174),
.B1(n_8),
.B2(n_10),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_178),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_193),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_186),
.B(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_177),
.C(n_8),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_1),
.A3(n_8),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_192),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_14),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_198),
.Y(n_200)
);


endmodule