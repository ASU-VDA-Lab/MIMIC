module fake_jpeg_4158_n_98 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_31),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_26),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_52)
);

CKINVDCx12_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_19),
.B1(n_21),
.B2(n_14),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_7),
.C(n_11),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_43),
.C(n_51),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_14),
.B1(n_18),
.B2(n_21),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_40),
.B1(n_52),
.B2(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_16),
.C(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_50),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_20),
.B(n_16),
.C(n_22),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_6),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_23),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_35),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_67),
.B1(n_41),
.B2(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_39),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_48),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_46),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_59),
.C(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_50),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_76),
.C(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_53),
.B(n_50),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_69),
.C(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_75),
.B1(n_64),
.B2(n_59),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_71),
.B(n_62),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_84),
.B(n_85),
.Y(n_93)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_93),
.A3(n_85),
.B1(n_91),
.B2(n_88),
.C1(n_62),
.C2(n_66),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_93),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);


endmodule