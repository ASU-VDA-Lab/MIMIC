module fake_jpeg_16853_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_1),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_38),
.B1(n_31),
.B2(n_4),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_54),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_35),
.A3(n_38),
.B1(n_18),
.B2(n_20),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_16),
.B1(n_6),
.B2(n_10),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_35),
.C(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_11),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_67),
.C(n_12),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_60),
.B(n_66),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_58),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_68),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_71),
.B1(n_72),
.B2(n_69),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_69),
.A3(n_15),
.B1(n_21),
.B2(n_22),
.C1(n_24),
.C2(n_14),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_25),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_26),
.Y(n_82)
);

NOR2x1p5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_28),
.Y(n_83)
);


endmodule