module real_jpeg_18796_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AND2x2_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_39),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

NAND2x1_ASAP7_75t_SL g74 ( 
.A(n_0),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_0),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_0),
.B(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_5),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_5),
.B(n_62),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_5),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_6),
.B(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_99),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_97),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_65),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_13),
.B(n_65),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_36),
.C(n_50),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_14),
.B(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_24),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_16),
.A2(n_25),
.B(n_35),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_16),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_17),
.A2(n_18),
.B1(n_93),
.B2(n_96),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_31),
.B(n_33),
.Y(n_30)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_31),
.Y(n_33)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_20),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_20),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_25),
.A2(n_121),
.B(n_123),
.C(n_127),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_25),
.B(n_121),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_25),
.A2(n_34),
.B1(n_121),
.B2(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_31),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_36),
.A2(n_50),
.B1(n_51),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.C(n_47),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_42),
.B1(n_80),
.B2(n_86),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_41),
.A2(n_42),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_47),
.Y(n_105)
);

OR2x4_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_57),
.C(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_81),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_134),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_107),
.B(n_108),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_118),
.B(n_142),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_115),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_111),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_111),
.B1(n_112),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_131),
.B(n_141),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_128),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_121),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_124),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_137),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_136),
.B(n_140),
.Y(n_131)
);


endmodule