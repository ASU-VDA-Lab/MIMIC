module fake_netlist_1_3831_n_571 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_571);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_571;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_43), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_76), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_38), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_20), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_46), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_15), .Y(n_87) );
NOR2xp33_ASAP7_75t_L g88 ( .A(n_12), .B(n_7), .Y(n_88) );
BUFx10_ASAP7_75t_L g89 ( .A(n_70), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_31), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_53), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_62), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_44), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_28), .B(n_64), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_11), .Y(n_97) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_6), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_58), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_69), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_35), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_60), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_55), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_33), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_10), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_72), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_49), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_32), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_52), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_45), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_41), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_109), .B(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
NOR2xp67_ASAP7_75t_L g124 ( .A(n_121), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_90), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_92), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_86), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_91), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_109), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_85), .B(n_1), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_85), .B(n_2), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_100), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_93), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_100), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
INVx5_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_95), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_118), .B(n_3), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
BUFx8_ASAP7_75t_SL g146 ( .A(n_126), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
NOR2xp33_ASAP7_75t_R g148 ( .A(n_138), .B(n_112), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_123), .B(n_81), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_138), .B(n_89), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_130), .Y(n_153) );
OR2x6_ASAP7_75t_L g154 ( .A(n_133), .B(n_116), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g155 ( .A1(n_122), .A2(n_99), .B1(n_108), .B2(n_97), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_138), .B(n_80), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
BUFx8_ASAP7_75t_SL g158 ( .A(n_138), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
OR2x2_ASAP7_75t_L g160 ( .A(n_134), .B(n_117), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_123), .B(n_101), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_141), .B(n_102), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_141), .B(n_103), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_125), .B(n_120), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_154), .A2(n_134), .B1(n_129), .B2(n_142), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_152), .B(n_141), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_159), .B(n_141), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_146), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_148), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_152), .B(n_125), .Y(n_178) );
BUFx8_ASAP7_75t_SL g179 ( .A(n_158), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_152), .B(n_128), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_156), .B(n_128), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_151), .B(n_129), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_151), .B(n_136), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
NOR2xp67_ASAP7_75t_L g191 ( .A(n_159), .B(n_161), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_156), .B(n_136), .Y(n_192) );
NAND3xp33_ASAP7_75t_SL g193 ( .A(n_160), .B(n_97), .C(n_99), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_156), .B(n_139), .Y(n_194) );
NOR2xp33_ASAP7_75t_SL g195 ( .A(n_154), .B(n_82), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_160), .B(n_149), .Y(n_197) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_149), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_150), .A2(n_139), .B1(n_140), .B2(n_142), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_150), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_178), .A2(n_173), .B(n_194), .Y(n_205) );
OAI22x1_ASAP7_75t_L g206 ( .A1(n_172), .A2(n_108), .B1(n_116), .B2(n_88), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_202), .Y(n_207) );
INVx5_ASAP7_75t_L g208 ( .A(n_202), .Y(n_208) );
AOI222xp33_ASAP7_75t_L g209 ( .A1(n_200), .A2(n_155), .B1(n_143), .B2(n_131), .C1(n_140), .C2(n_83), .Y(n_209) );
NOR2x1_ASAP7_75t_SL g210 ( .A(n_183), .B(n_159), .Y(n_210) );
OAI22xp5_ASAP7_75t_SL g211 ( .A1(n_200), .A2(n_155), .B1(n_106), .B2(n_119), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_181), .A2(n_163), .B(n_164), .C(n_162), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_198), .B(n_162), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_202), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_198), .A2(n_170), .B1(n_166), .B2(n_157), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_183), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_178), .A2(n_163), .B(n_164), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_181), .A2(n_170), .B(n_166), .C(n_157), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_183), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_185), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_193), .B(n_159), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_197), .B(n_148), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_194), .A2(n_157), .B(n_87), .C(n_137), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_197), .B(n_161), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_180), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_SL g227 ( .A1(n_184), .A2(n_192), .B(n_195), .C(n_201), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_185), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_172), .A2(n_124), .B1(n_87), .B2(n_110), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_188), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_188), .Y(n_233) );
BUFx8_ASAP7_75t_SL g234 ( .A(n_179), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_196), .A2(n_96), .B(n_107), .C(n_105), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_193), .B(n_161), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_188), .Y(n_237) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_173), .A2(n_113), .B(n_115), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_227), .A2(n_96), .B(n_184), .C(n_192), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_218), .A2(n_197), .B(n_187), .C(n_189), .Y(n_241) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_205), .A2(n_165), .B(n_167), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_224), .A2(n_186), .B(n_203), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_208), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_211), .B(n_197), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_230), .Y(n_248) );
AOI31xp67_ASAP7_75t_L g249 ( .A1(n_223), .A2(n_168), .A3(n_167), .B(n_165), .Y(n_249) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_217), .A2(n_186), .B(n_203), .Y(n_250) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_238), .A2(n_168), .B(n_165), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_211), .A2(n_197), .B1(n_171), .B2(n_195), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_223), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_208), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_226), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_208), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_212), .A2(n_187), .B(n_189), .C(n_135), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_214), .A2(n_94), .B(n_113), .C(n_115), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_213), .A2(n_171), .B1(n_201), .B2(n_137), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_186), .B(n_203), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_209), .A2(n_199), .B1(n_177), .B2(n_124), .Y(n_261) );
OR2x6_ASAP7_75t_L g262 ( .A(n_216), .B(n_199), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_225), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_238), .A2(n_167), .B(n_168), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_215), .B(n_199), .Y(n_266) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_214), .A2(n_190), .B(n_182), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_252), .A2(n_215), .B1(n_222), .B2(n_208), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g269 ( .A1(n_261), .A2(n_209), .B1(n_235), .B2(n_236), .C(n_221), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_247), .B(n_231), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_263), .B(n_206), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_245), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_263), .A2(n_206), .B1(n_238), .B2(n_220), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_245), .Y(n_274) );
AND3x1_ASAP7_75t_L g275 ( .A(n_254), .B(n_234), .C(n_176), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_266), .A2(n_208), .B1(n_220), .B2(n_207), .Y(n_276) );
INVx4_ASAP7_75t_SL g277 ( .A(n_246), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_239), .A2(n_208), .B(n_210), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_241), .A2(n_225), .B1(n_237), .B2(n_229), .C(n_137), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_253), .B(n_228), .Y(n_282) );
INVx8_ASAP7_75t_L g283 ( .A(n_240), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_240), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_241), .A2(n_210), .B(n_182), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_248), .A2(n_228), .B1(n_232), .B2(n_216), .Y(n_286) );
NAND4xp25_ASAP7_75t_L g287 ( .A(n_257), .B(n_135), .C(n_132), .D(n_199), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_266), .A2(n_174), .B(n_182), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_255), .B(n_228), .Y(n_289) );
BUFx4f_ASAP7_75t_SL g290 ( .A(n_246), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_259), .A2(n_233), .B1(n_219), .B2(n_232), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_259), .A2(n_232), .B1(n_216), .B2(n_98), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_272), .B(n_255), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_281), .B(n_240), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_281), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_290), .Y(n_297) );
OR2x2_ASAP7_75t_SL g298 ( .A(n_271), .B(n_98), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_282), .B(n_240), .Y(n_302) );
NAND2xp33_ASAP7_75t_R g303 ( .A(n_270), .B(n_254), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_283), .Y(n_304) );
CKINVDCx14_ASAP7_75t_R g305 ( .A(n_275), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_284), .B(n_240), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_273), .B(n_240), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_286), .B(n_240), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_273), .B(n_257), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_251), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_279), .B(n_251), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_296), .B(n_251), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_295), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
AOI21x1_ASAP7_75t_L g322 ( .A1(n_313), .A2(n_242), .B(n_278), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_301), .B(n_251), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_295), .B(n_265), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_304), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_301), .B(n_265), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_300), .B(n_265), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_294), .Y(n_330) );
INVx5_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_306), .B(n_265), .Y(n_332) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_309), .B(n_254), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_311), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_311), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_312), .B(n_283), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_314), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_305), .A2(n_269), .B1(n_258), .B2(n_98), .C(n_287), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_306), .B(n_283), .Y(n_341) );
OAI31xp33_ASAP7_75t_L g342 ( .A1(n_304), .A2(n_268), .A3(n_291), .B(n_292), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_302), .B(n_264), .Y(n_343) );
AO21x2_ASAP7_75t_L g344 ( .A1(n_315), .A2(n_285), .B(n_242), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_302), .B(n_244), .Y(n_346) );
INVx3_ASAP7_75t_SL g347 ( .A(n_331), .Y(n_347) );
OAI33xp33_ASAP7_75t_L g348 ( .A1(n_335), .A2(n_132), .A3(n_135), .B1(n_293), .B2(n_276), .B3(n_110), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_345), .B(n_298), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_335), .B(n_315), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_326), .B(n_297), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_326), .B(n_316), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_326), .B(n_3), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_336), .B(n_308), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_340), .B(n_308), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_321), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_345), .B(n_298), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
OAI21xp33_ASAP7_75t_SL g363 ( .A1(n_337), .A2(n_299), .B(n_310), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_336), .B(n_308), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_345), .B(n_312), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_312), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_328), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_327), .B(n_307), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_338), .B(n_307), .Y(n_371) );
NAND4xp25_ASAP7_75t_L g372 ( .A(n_339), .B(n_303), .C(n_292), .D(n_310), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_340), .Y(n_373) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_320), .B(n_309), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_334), .B(n_98), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_337), .B(n_250), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_324), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_338), .B(n_98), .Y(n_380) );
OAI33xp33_ASAP7_75t_L g381 ( .A1(n_323), .A2(n_82), .A3(n_104), .B1(n_111), .B2(n_114), .B3(n_9), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_332), .B(n_250), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_323), .B(n_144), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_332), .B(n_250), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_329), .B(n_243), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_319), .Y(n_386) );
OR2x4_ASAP7_75t_L g387 ( .A(n_341), .B(n_318), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_337), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_353), .B(n_331), .Y(n_390) );
NOR2xp33_ASAP7_75t_SL g391 ( .A(n_375), .B(n_331), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_380), .B(n_329), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_380), .B(n_325), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_387), .A2(n_331), .B1(n_337), .B2(n_341), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_387), .A2(n_331), .B1(n_337), .B2(n_320), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_370), .B(n_343), .Y(n_399) );
OAI21xp5_ASAP7_75t_SL g400 ( .A1(n_389), .A2(n_339), .B(n_342), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_366), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_351), .B(n_325), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_370), .B(n_343), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_371), .B(n_331), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
OR2x6_ASAP7_75t_L g407 ( .A(n_375), .B(n_318), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_379), .B(n_344), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_351), .B(n_344), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_388), .B(n_344), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_389), .B(n_344), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_376), .B(n_342), .C(n_144), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_368), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_371), .B(n_322), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_358), .B(n_333), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_349), .B(n_352), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_349), .B(n_322), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_355), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_352), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_360), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_362), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_357), .B(n_333), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_357), .B(n_4), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_360), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_372), .A2(n_104), .B(n_111), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_350), .B(n_361), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_373), .B(n_144), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_359), .Y(n_429) );
NAND2x1_ASAP7_75t_L g430 ( .A(n_375), .B(n_254), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_369), .B(n_144), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g433 ( .A(n_386), .B(n_4), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_347), .B(n_246), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_367), .B(n_5), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_378), .B(n_144), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_383), .B(n_144), .C(n_145), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_350), .B(n_5), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_378), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_359), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_387), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_347), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_397), .B(n_381), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
BUFx12f_ASAP7_75t_L g445 ( .A(n_438), .Y(n_445) );
AOI221xp5_ASAP7_75t_SL g446 ( .A1(n_419), .A2(n_394), .B1(n_396), .B2(n_395), .C(n_441), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_400), .A2(n_361), .B1(n_347), .B2(n_383), .C(n_386), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_427), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_394), .A2(n_374), .B1(n_377), .B2(n_367), .Y(n_449) );
OAI21xp33_ASAP7_75t_SL g450 ( .A1(n_442), .A2(n_374), .B(n_365), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_399), .B(n_365), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_404), .B(n_377), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_433), .A2(n_377), .B1(n_364), .B2(n_382), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_405), .B(n_364), .Y(n_456) );
OAI322xp33_ASAP7_75t_L g457 ( .A1(n_408), .A2(n_384), .A3(n_382), .B1(n_385), .B2(n_348), .C1(n_114), .C2(n_169), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_403), .B(n_384), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_414), .B(n_385), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_391), .B(n_422), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_435), .A2(n_262), .B1(n_256), .B2(n_232), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_426), .B(n_256), .C(n_233), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_409), .A2(n_169), .B1(n_153), .B2(n_232), .C(n_13), .Y(n_463) );
AO22x1_ASAP7_75t_L g464 ( .A1(n_390), .A2(n_256), .B1(n_244), .B2(n_9), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_403), .B(n_6), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_424), .A2(n_256), .B(n_262), .C(n_219), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_409), .B(n_8), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_437), .B(n_243), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_420), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
NAND3xp33_ASAP7_75t_SL g473 ( .A(n_430), .B(n_8), .C(n_13), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_407), .A2(n_262), .B1(n_243), .B2(n_169), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_393), .B(n_14), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_416), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_439), .B(n_16), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_398), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_401), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_429), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_393), .B(n_16), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_392), .A2(n_262), .B1(n_169), .B2(n_244), .Y(n_484) );
OAI22x1_ASAP7_75t_L g485 ( .A1(n_411), .A2(n_434), .B1(n_410), .B2(n_412), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_415), .B(n_17), .Y(n_486) );
NAND4xp25_ASAP7_75t_L g487 ( .A(n_411), .B(n_17), .C(n_18), .D(n_19), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_402), .B(n_18), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g489 ( .A(n_428), .B(n_267), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_440), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_467), .B(n_413), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_443), .Y(n_492) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_453), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_469), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_471), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_478), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_459), .B(n_423), .Y(n_497) );
OAI21xp5_ASAP7_75t_SL g498 ( .A1(n_487), .A2(n_392), .B(n_428), .Y(n_498) );
NOR4xp25_ASAP7_75t_L g499 ( .A(n_444), .B(n_436), .C(n_432), .D(n_418), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_472), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_474), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_443), .A2(n_436), .B1(n_432), .B2(n_418), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_477), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_480), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_458), .B(n_19), .Y(n_505) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_446), .A2(n_169), .B1(n_288), .B2(n_153), .C(n_199), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_481), .Y(n_507) );
AOI211xp5_ASAP7_75t_L g508 ( .A1(n_450), .A2(n_169), .B(n_260), .C(n_191), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_473), .B(n_260), .C(n_190), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_447), .A2(n_262), .B1(n_169), .B2(n_267), .Y(n_510) );
OAI32xp33_ASAP7_75t_L g511 ( .A1(n_444), .A2(n_175), .A3(n_249), .B1(n_27), .B2(n_29), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_452), .B(n_153), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_486), .A2(n_153), .B1(n_190), .B2(n_174), .C(n_204), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_490), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_486), .A2(n_267), .B1(n_260), .B2(n_153), .Y(n_515) );
XOR2x2_ASAP7_75t_L g516 ( .A(n_473), .B(n_23), .Y(n_516) );
XNOR2x1_ASAP7_75t_L g517 ( .A(n_465), .B(n_24), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_L g518 ( .A1(n_460), .A2(n_249), .B(n_174), .C(n_161), .Y(n_518) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_460), .B(n_267), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_448), .Y(n_520) );
AOI21xp33_ASAP7_75t_L g521 ( .A1(n_468), .A2(n_30), .B(n_34), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g522 ( .A1(n_453), .A2(n_175), .B1(n_153), .B2(n_40), .C1(n_42), .C2(n_47), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_490), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_508), .B(n_485), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_491), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_492), .A2(n_488), .B(n_479), .C(n_483), .Y(n_526) );
NAND4xp75_ASAP7_75t_L g527 ( .A(n_506), .B(n_502), .C(n_519), .D(n_476), .Y(n_527) );
NOR3xp33_ASAP7_75t_SL g528 ( .A(n_506), .B(n_449), .C(n_457), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_493), .A2(n_464), .B(n_455), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_499), .B(n_451), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_498), .A2(n_445), .B1(n_454), .B2(n_461), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_520), .A2(n_462), .B1(n_456), .B2(n_463), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_512), .Y(n_533) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_517), .A2(n_462), .B(n_466), .Y(n_534) );
AOI322xp5_ASAP7_75t_L g535 ( .A1(n_497), .A2(n_482), .A3(n_484), .B1(n_470), .B2(n_475), .C1(n_466), .C2(n_489), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g536 ( .A1(n_505), .A2(n_470), .B(n_489), .Y(n_536) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_522), .A2(n_510), .B(n_509), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_522), .A2(n_153), .B(n_175), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_496), .A2(n_153), .B1(n_175), .B2(n_204), .Y(n_539) );
OAI21xp33_ASAP7_75t_SL g540 ( .A1(n_491), .A2(n_36), .B(n_39), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g541 ( .A(n_516), .B(n_48), .Y(n_541) );
AOI31xp33_ASAP7_75t_L g542 ( .A1(n_513), .A2(n_50), .A3(n_51), .B(n_54), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_515), .A2(n_191), .B1(n_204), .B2(n_61), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_533), .B(n_494), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_531), .A2(n_507), .B1(n_500), .B2(n_501), .C(n_503), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_535), .B(n_513), .C(n_521), .Y(n_546) );
AOI21xp33_ASAP7_75t_SL g547 ( .A1(n_524), .A2(n_521), .B(n_504), .Y(n_547) );
OAI211xp5_ASAP7_75t_L g548 ( .A1(n_534), .A2(n_511), .B(n_495), .C(n_523), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_525), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_530), .Y(n_550) );
AOI222xp33_ASAP7_75t_L g551 ( .A1(n_537), .A2(n_514), .B1(n_518), .B2(n_204), .C1(n_65), .C2(n_66), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_528), .B(n_204), .C(n_59), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_532), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_529), .A2(n_204), .B1(n_63), .B2(n_67), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_546), .A2(n_540), .B(n_527), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_553), .B(n_536), .Y(n_556) );
NOR2x1p5_ASAP7_75t_L g557 ( .A(n_550), .B(n_526), .Y(n_557) );
NAND3xp33_ASAP7_75t_SL g558 ( .A(n_547), .B(n_538), .C(n_539), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_544), .B(n_545), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_554), .A2(n_541), .B(n_542), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_556), .Y(n_561) );
OR2x4_ASAP7_75t_L g562 ( .A(n_558), .B(n_549), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g563 ( .A(n_555), .B(n_551), .C(n_548), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_563), .A2(n_559), .B(n_552), .Y(n_564) );
OAI22x1_ASAP7_75t_SL g565 ( .A1(n_561), .A2(n_557), .B1(n_560), .B2(n_544), .Y(n_565) );
OAI22xp5_ASAP7_75t_SL g566 ( .A1(n_564), .A2(n_562), .B1(n_543), .B2(n_538), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_565), .B(n_56), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_567), .A2(n_204), .B1(n_71), .B2(n_73), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_568), .Y(n_569) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_569), .A2(n_566), .B(n_74), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_570), .A2(n_68), .B1(n_75), .B2(n_77), .C(n_79), .Y(n_571) );
endmodule