module fake_jpeg_12585_n_165 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_79),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_1),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_88),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_52),
.B1(n_61),
.B2(n_69),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_66),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_52),
.B1(n_61),
.B2(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_100),
.Y(n_135)
);

AO22x2_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_53),
.B1(n_64),
.B2(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_106),
.B1(n_8),
.B2(n_13),
.Y(n_134)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_68),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_64),
.B(n_65),
.C(n_59),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_104),
.B(n_107),
.Y(n_119)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_58),
.B(n_56),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_50),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_117),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_47),
.B(n_46),
.C(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_2),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_3),
.B(n_4),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_4),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_134),
.B1(n_107),
.B2(n_17),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_29),
.C(n_11),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_140),
.B(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_107),
.B1(n_19),
.B2(n_22),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_128),
.B1(n_126),
.B2(n_132),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_149),
.B1(n_124),
.B2(n_36),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_16),
.B(n_23),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_133),
.B(n_136),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_25),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_28),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_150),
.C(n_35),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_43),
.B1(n_33),
.B2(n_34),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_32),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_147),
.B1(n_141),
.B2(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_159),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_155),
.B1(n_156),
.B2(n_149),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_145),
.Y(n_165)
);


endmodule