module fake_jpeg_1024_n_202 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_38),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_91),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_93),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_61),
.B1(n_72),
.B2(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_57),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_90),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_65),
.B(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_52),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_58),
.B1(n_59),
.B2(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_99),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_96),
.Y(n_124)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_106),
.Y(n_134)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_61),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_112),
.Y(n_115)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_57),
.B(n_82),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_0),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_105),
.B1(n_109),
.B2(n_104),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_122),
.B1(n_126),
.B2(n_131),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_68),
.B1(n_66),
.B2(n_71),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_125),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_51),
.B(n_55),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_67),
.B1(n_60),
.B2(n_56),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_68),
.B1(n_24),
.B2(n_25),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_0),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_48),
.B1(n_22),
.B2(n_27),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_143),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_142),
.C(n_149),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_146),
.C(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_134),
.B(n_1),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_2),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_3),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_4),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_7),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_29),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_4),
.CON(n_160),
.SN(n_160)
);

OAI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_12),
.B(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_17),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_172),
.B1(n_139),
.B2(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_10),
.B(n_11),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_173),
.B(n_14),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_36),
.B(n_47),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_141),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_164),
.B1(n_170),
.B2(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_177),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_164),
.B(n_34),
.C(n_46),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_32),
.C(n_45),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_173),
.C(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_15),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_183),
.B1(n_161),
.B2(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_187),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_167),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_190),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_189),
.B(n_166),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_168),
.Y(n_190)
);

NOR2x1_ASAP7_75t_SL g191 ( 
.A(n_190),
.B(n_177),
.Y(n_191)
);

NAND4xp25_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_158),
.C(n_185),
.D(n_186),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_160),
.B1(n_159),
.B2(n_171),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_196),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_188),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_197),
.C(n_193),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_199),
.A2(n_193),
.B(n_30),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_39),
.B(n_41),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_42),
.Y(n_202)
);


endmodule