module fake_jpeg_8862_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_31),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_50),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_22),
.B(n_27),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_17),
.B1(n_24),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_59),
.B1(n_17),
.B2(n_39),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_17),
.B1(n_24),
.B2(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_28),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_67),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_84),
.B1(n_61),
.B2(n_44),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_39),
.B(n_40),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_36),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_26),
.B1(n_19),
.B2(n_21),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_43),
.B1(n_44),
.B2(n_56),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_40),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_58),
.B(n_40),
.C(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_57),
.B1(n_55),
.B2(n_19),
.Y(n_93)
);

AOI22x1_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_59),
.B1(n_48),
.B2(n_41),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_73),
.Y(n_129)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_107),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_64),
.B1(n_67),
.B2(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_98),
.B1(n_103),
.B2(n_87),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_113),
.B1(n_85),
.B2(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_106),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_43),
.B1(n_64),
.B2(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_37),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_75),
.Y(n_114)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_111),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_41),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_110),
.C(n_95),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_38),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_75),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_129),
.B1(n_88),
.B2(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_132),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_81),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_126),
.C(n_37),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_133),
.B1(n_137),
.B2(n_37),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_70),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_42),
.B(n_20),
.Y(n_158)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_86),
.B1(n_80),
.B2(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_86),
.B1(n_83),
.B2(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_106),
.B1(n_109),
.B2(n_91),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_149),
.B1(n_119),
.B2(n_120),
.Y(n_171)
);

NOR4xp25_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_38),
.C(n_36),
.D(n_112),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_131),
.B(n_133),
.C(n_127),
.D(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_11),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_145),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_152),
.C(n_121),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_154),
.B1(n_129),
.B2(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_74),
.C(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_74),
.B1(n_21),
.B2(n_20),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_78),
.B1(n_63),
.B2(n_53),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_157),
.B1(n_42),
.B2(n_52),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_20),
.B1(n_42),
.B2(n_52),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_138),
.B(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_162),
.Y(n_173)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_29),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_164),
.B(n_165),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_175),
.C(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_176),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_131),
.B1(n_123),
.B2(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_182),
.B1(n_184),
.B2(n_143),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_148),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_116),
.B(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_29),
.B1(n_23),
.B2(n_2),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_29),
.C(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_162),
.C(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_192),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_183),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NOR4xp25_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_141),
.C(n_152),
.D(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_143),
.B(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_151),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_1),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_201),
.B1(n_207),
.B2(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_139),
.C(n_144),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_172),
.C(n_174),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_203),
.B(n_9),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_210),
.C(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_186),
.C(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_23),
.C(n_2),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_216),
.B1(n_207),
.B2(n_199),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_13),
.B(n_7),
.C(n_8),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_1),
.C(n_3),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_223),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_6),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_9),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_218),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_188),
.B(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_188),
.B(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_235),
.B1(n_236),
.B2(n_216),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_9),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_190),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_196),
.B(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_238),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_204),
.B1(n_196),
.B2(n_210),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_202),
.B1(n_200),
.B2(n_5),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_228),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_219),
.C(n_217),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_224),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_238),
.A2(n_234),
.B(n_235),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_237),
.B(n_230),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_247),
.B(n_232),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_6),
.C(n_10),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_225),
.CI(n_226),
.CON(n_255),
.SN(n_255)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_256),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_257),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_246),
.B1(n_248),
.B2(n_250),
.Y(n_259)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_262),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_13),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_253),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_256),
.B(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_263),
.C(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_269),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_255),
.B(n_12),
.C(n_13),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_268),
.C(n_4),
.Y(n_274)
);

NAND4xp25_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_264),
.C(n_260),
.D(n_12),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_272),
.B(n_3),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_275),
.B(n_3),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_3),
.B(n_5),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_5),
.Y(n_278)
);


endmodule