module real_aes_4989_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_577;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_1049;
wire n_466;
wire n_636;
wire n_976;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_755;
wire n_656;
wire n_284;
wire n_316;
wire n_532;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_303;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_366;
wire n_346;
wire n_727;
wire n_1056;
wire n_293;
wire n_358;
wire n_385;
wire n_397;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_1043;
wire n_850;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_473;
wire n_465;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_0), .A2(n_249), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_1), .A2(n_123), .B1(n_457), .B2(n_459), .Y(n_456) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_2), .Y(n_293) );
AND2x4_ASAP7_75t_L g765 ( .A(n_2), .B(n_273), .Y(n_765) );
AND2x4_ASAP7_75t_L g770 ( .A(n_2), .B(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_3), .A2(n_234), .B1(n_448), .B2(n_449), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_4), .A2(n_176), .B1(n_413), .B2(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g742 ( .A(n_5), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_6), .A2(n_62), .B1(n_391), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_7), .A2(n_40), .B1(n_436), .B2(n_438), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_8), .A2(n_18), .B1(n_431), .B2(n_433), .Y(n_668) );
AOI21xp33_ASAP7_75t_SL g657 ( .A1(n_9), .A2(n_391), .B(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g357 ( .A1(n_10), .A2(n_358), .B(n_359), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_11), .A2(n_121), .B1(n_404), .B2(n_513), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_12), .A2(n_196), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_13), .A2(n_129), .B1(n_454), .B2(n_455), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_14), .A2(n_673), .B(n_674), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_15), .A2(n_19), .B1(n_370), .B2(n_378), .Y(n_689) );
XNOR2x2_ASAP7_75t_L g736 ( .A(n_16), .B(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_16), .A2(n_87), .B1(n_774), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_17), .A2(n_155), .B1(n_404), .B2(n_585), .Y(n_1041) );
AO22x1_ASAP7_75t_L g558 ( .A1(n_20), .A2(n_22), .B1(n_559), .B2(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g792 ( .A(n_21), .Y(n_792) );
INVx1_ASAP7_75t_L g571 ( .A(n_23), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_24), .A2(n_88), .B1(n_377), .B2(n_381), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_25), .A2(n_74), .B1(n_431), .B2(n_459), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_26), .A2(n_1027), .B1(n_1028), .B2(n_1055), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_26), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_27), .A2(n_218), .B1(n_499), .B2(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_28), .A2(n_50), .B1(n_462), .B2(n_463), .C(n_464), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_29), .A2(n_84), .B1(n_762), .B2(n_766), .Y(n_761) );
INVx1_ASAP7_75t_SL g876 ( .A(n_30), .Y(n_876) );
INVx1_ASAP7_75t_SL g517 ( .A(n_31), .Y(n_517) );
INVx1_ASAP7_75t_L g586 ( .A(n_32), .Y(n_586) );
INVx1_ASAP7_75t_L g465 ( .A(n_33), .Y(n_465) );
INVx1_ASAP7_75t_L g700 ( .A(n_34), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_35), .A2(n_42), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_36), .A2(n_251), .B1(n_568), .B2(n_1001), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_37), .B(n_216), .Y(n_291) );
INVx1_ASAP7_75t_L g327 ( .A(n_37), .Y(n_327) );
INVxp67_ASAP7_75t_L g337 ( .A(n_37), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_38), .A2(n_95), .B1(n_769), .B2(n_781), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_39), .A2(n_77), .B1(n_419), .B2(n_438), .Y(n_1002) );
INVx1_ASAP7_75t_L g505 ( .A(n_41), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_43), .A2(n_57), .B1(n_374), .B2(n_375), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_44), .A2(n_149), .B1(n_344), .B2(n_626), .Y(n_699) );
INVx1_ASAP7_75t_L g628 ( .A(n_45), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_46), .A2(n_111), .B1(n_424), .B2(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_47), .B(n_311), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_48), .A2(n_244), .B1(n_431), .B2(n_433), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_49), .A2(n_119), .B1(n_1043), .B2(n_1045), .Y(n_1042) );
INVx1_ASAP7_75t_SL g508 ( .A(n_51), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_52), .A2(n_272), .B1(n_591), .B2(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_53), .A2(n_105), .B1(n_391), .B2(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g659 ( .A(n_54), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_55), .A2(n_281), .B1(n_778), .B2(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g583 ( .A(n_56), .Y(n_583) );
INVx1_ASAP7_75t_L g400 ( .A(n_58), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_59), .A2(n_221), .B1(n_330), .B2(n_369), .Y(n_624) );
INVxp67_ASAP7_75t_R g794 ( .A(n_60), .Y(n_794) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_61), .A2(n_626), .B(n_627), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_63), .A2(n_264), .B1(n_459), .B2(n_547), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_64), .A2(n_145), .B1(n_431), .B2(n_433), .Y(n_430) );
INVx1_ASAP7_75t_SL g515 ( .A(n_65), .Y(n_515) );
INVx1_ASAP7_75t_L g1018 ( .A(n_66), .Y(n_1018) );
INVx2_ASAP7_75t_L g288 ( .A(n_67), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_68), .A2(n_107), .B1(n_424), .B2(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g393 ( .A(n_69), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_70), .A2(n_183), .B1(n_340), .B2(n_344), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_71), .A2(n_127), .B1(n_451), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_72), .A2(n_140), .B1(n_424), .B2(n_610), .Y(n_740) );
INVx1_ASAP7_75t_L g764 ( .A(n_73), .Y(n_764) );
AND2x4_ASAP7_75t_L g767 ( .A(n_73), .B(n_288), .Y(n_767) );
INVx1_ASAP7_75t_SL g800 ( .A(n_73), .Y(n_800) );
INVx1_ASAP7_75t_SL g511 ( .A(n_75), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_76), .A2(n_86), .B1(n_530), .B2(n_533), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_78), .A2(n_104), .B1(n_330), .B2(n_340), .Y(n_694) );
INVx1_ASAP7_75t_L g588 ( .A(n_79), .Y(n_588) );
INVx1_ASAP7_75t_L g606 ( .A(n_80), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_81), .A2(n_194), .B1(n_715), .B2(n_718), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_82), .A2(n_210), .B1(n_774), .B2(n_799), .Y(n_810) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_83), .Y(n_311) );
XOR2x2_ASAP7_75t_L g989 ( .A(n_84), .B(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_84), .A2(n_1026), .B1(n_1056), .B2(n_1058), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_85), .A2(n_94), .B1(n_448), .B2(n_454), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_89), .B(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1014 ( .A(n_90), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_91), .A2(n_277), .B1(n_421), .B2(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g579 ( .A(n_92), .Y(n_579) );
INVx1_ASAP7_75t_L g711 ( .A(n_93), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g790 ( .A(n_96), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_97), .A2(n_180), .B1(n_769), .B2(n_772), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_98), .A2(n_248), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_99), .A2(n_125), .B1(n_377), .B2(n_381), .Y(n_690) );
INVx1_ASAP7_75t_L g312 ( .A(n_100), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_100), .B(n_215), .Y(n_334) );
OAI22x1_ASAP7_75t_L g663 ( .A1(n_101), .A2(n_664), .B1(n_669), .B2(n_680), .Y(n_663) );
NAND5xp2_ASAP7_75t_SL g664 ( .A(n_101), .B(n_665), .C(n_666), .D(n_667), .E(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g747 ( .A(n_102), .Y(n_747) );
XNOR2x1_ASAP7_75t_L g302 ( .A(n_103), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_106), .B(n_462), .Y(n_597) );
INVx1_ASAP7_75t_SL g540 ( .A(n_108), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_109), .A2(n_228), .B1(n_459), .B2(n_547), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_110), .A2(n_243), .B1(n_438), .B2(n_527), .Y(n_526) );
INVx2_ASAP7_75t_R g385 ( .A(n_112), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_113), .A2(n_212), .B1(n_424), .B2(n_485), .Y(n_1032) );
AOI21xp5_ASAP7_75t_L g1046 ( .A1(n_114), .A2(n_1047), .B(n_1049), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_115), .A2(n_138), .B1(n_601), .B2(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_116), .B(n_604), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_117), .A2(n_182), .B1(n_762), .B2(n_779), .Y(n_806) );
INVx1_ASAP7_75t_L g822 ( .A(n_118), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_120), .A2(n_242), .B1(n_438), .B2(n_451), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_122), .A2(n_199), .B1(n_436), .B2(n_438), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_124), .A2(n_250), .B1(n_377), .B2(n_378), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_126), .A2(n_604), .B(n_605), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_128), .A2(n_163), .B1(n_470), .B2(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_130), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_131), .B(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_132), .A2(n_198), .B1(n_599), .B2(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g481 ( .A(n_133), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_134), .A2(n_174), .B1(n_451), .B2(n_452), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_135), .A2(n_202), .B1(n_374), .B2(n_375), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_136), .A2(n_187), .B1(n_766), .B2(n_778), .Y(n_877) );
INVx1_ASAP7_75t_L g360 ( .A(n_137), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_139), .A2(n_256), .B1(n_424), .B2(n_485), .Y(n_665) );
INVx1_ASAP7_75t_L g1052 ( .A(n_141), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_142), .A2(n_235), .B1(n_419), .B2(n_452), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_143), .A2(n_156), .B1(n_615), .B2(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_144), .A2(n_209), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_146), .A2(n_262), .B1(n_369), .B2(n_370), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_147), .A2(n_278), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_148), .A2(n_188), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_150), .A2(n_181), .B1(n_470), .B2(n_601), .Y(n_753) );
INVx1_ASAP7_75t_L g675 ( .A(n_151), .Y(n_675) );
INVx1_ASAP7_75t_L g578 ( .A(n_152), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_153), .A2(n_225), .B1(n_340), .B2(n_344), .Y(n_339) );
INVx1_ASAP7_75t_L g998 ( .A(n_154), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_157), .A2(n_162), .B1(n_452), .B2(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_158), .A2(n_217), .B1(n_370), .B2(n_378), .Y(n_631) );
INVx1_ASAP7_75t_L g996 ( .A(n_159), .Y(n_996) );
AOI21xp33_ASAP7_75t_SL g1010 ( .A1(n_160), .A2(n_1011), .B(n_1013), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_161), .A2(n_208), .B1(n_419), .B2(n_421), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_164), .A2(n_270), .B1(n_547), .B2(n_566), .Y(n_616) );
INVx1_ASAP7_75t_L g507 ( .A(n_165), .Y(n_507) );
INVx1_ASAP7_75t_L g389 ( .A(n_166), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_167), .A2(n_252), .B1(n_802), .B2(n_803), .Y(n_811) );
INVx1_ASAP7_75t_L g825 ( .A(n_168), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_169), .A2(n_269), .B1(n_448), .B2(n_615), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_170), .A2(n_245), .B1(n_306), .B2(n_382), .Y(n_630) );
INVx1_ASAP7_75t_L g823 ( .A(n_171), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_172), .A2(n_189), .B1(n_496), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_173), .A2(n_253), .B1(n_306), .B2(n_382), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_175), .A2(n_271), .B1(n_560), .B2(n_615), .Y(n_614) );
XNOR2x1_ASAP7_75t_L g594 ( .A(n_177), .B(n_595), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_178), .Y(n_661) );
INVx1_ASAP7_75t_L g402 ( .A(n_179), .Y(n_402) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_184), .B(n_556), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_185), .A2(n_224), .B1(n_426), .B2(n_452), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_186), .B(n_1054), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_190), .A2(n_263), .B1(n_419), .B2(n_452), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_191), .A2(n_227), .B1(n_306), .B2(n_330), .Y(n_305) );
INVx1_ASAP7_75t_L g494 ( .A(n_192), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_193), .Y(n_827) );
OA22x2_ASAP7_75t_L g317 ( .A1(n_195), .A2(n_216), .B1(n_311), .B2(n_315), .Y(n_317) );
INVx1_ASAP7_75t_L g349 ( .A(n_195), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_197), .B(n_1009), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_200), .A2(n_231), .B1(n_599), .B2(n_656), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_201), .A2(n_236), .B1(n_491), .B2(n_492), .C(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g697 ( .A(n_203), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_204), .A2(n_257), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI221x1_ASAP7_75t_L g708 ( .A1(n_205), .A2(n_239), .B1(n_513), .B2(n_709), .C(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g1005 ( .A(n_206), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_207), .A2(n_211), .B1(n_436), .B2(n_438), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_213), .A2(n_254), .B1(n_431), .B2(n_1035), .Y(n_1034) );
CKINVDCx6p67_ASAP7_75t_R g788 ( .A(n_214), .Y(n_788) );
INVx1_ASAP7_75t_L g329 ( .A(n_215), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_215), .B(n_347), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g350 ( .A1(n_216), .A2(n_229), .B(n_338), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_219), .A2(n_280), .B1(n_769), .B2(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_220), .A2(n_255), .B1(n_436), .B2(n_438), .Y(n_435) );
INVx1_ASAP7_75t_SL g1021 ( .A(n_222), .Y(n_1021) );
INVx1_ASAP7_75t_SL g548 ( .A(n_223), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_226), .A2(n_241), .B1(n_498), .B2(n_499), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_229), .B(n_266), .Y(n_292) );
INVx1_ASAP7_75t_L g314 ( .A(n_229), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_230), .A2(n_261), .B1(n_374), .B2(n_375), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_232), .A2(n_354), .B(n_746), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_233), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_237), .B(n_492), .Y(n_652) );
INVx1_ASAP7_75t_L g618 ( .A(n_238), .Y(n_618) );
OAI21x1_ASAP7_75t_L g705 ( .A1(n_240), .A2(n_706), .B(n_729), .Y(n_705) );
INVx1_ASAP7_75t_L g732 ( .A(n_240), .Y(n_732) );
INVx1_ASAP7_75t_SL g1004 ( .A(n_246), .Y(n_1004) );
INVx1_ASAP7_75t_L g407 ( .A(n_247), .Y(n_407) );
INVx1_ASAP7_75t_SL g1016 ( .A(n_258), .Y(n_1016) );
INVx1_ASAP7_75t_SL g539 ( .A(n_259), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_260), .A2(n_276), .B1(n_391), .B2(n_404), .Y(n_500) );
INVx1_ASAP7_75t_L g575 ( .A(n_265), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_266), .B(n_322), .Y(n_321) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_267), .A2(n_369), .B(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_268), .A2(n_274), .B1(n_421), .B2(n_451), .Y(n_739) );
INVx1_ASAP7_75t_L g771 ( .A(n_273), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_275), .B(n_519), .Y(n_678) );
XNOR2x1_ASAP7_75t_L g444 ( .A(n_279), .B(n_445), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_294), .B(n_755), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx4_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .C(n_293), .Y(n_285) );
AND2x2_ASAP7_75t_L g984 ( .A(n_286), .B(n_985), .Y(n_984) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_286), .B(n_986), .Y(n_1057) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OA21x2_ASAP7_75t_L g1059 ( .A1(n_287), .A2(n_800), .B(n_1060), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g763 ( .A(n_288), .B(n_764), .Y(n_763) );
AND3x4_ASAP7_75t_L g799 ( .A(n_288), .B(n_770), .C(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_289), .B(n_986), .Y(n_985) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_290), .A2(n_364), .B(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g986 ( .A(n_293), .Y(n_986) );
XNOR2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_552), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_477), .Y(n_296) );
OAI22x1_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_442), .B2(n_476), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_383), .B1(n_384), .B2(n_441), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g441 ( .A(n_302), .Y(n_441) );
NOR2x1_ASAP7_75t_L g303 ( .A(n_304), .B(n_367), .Y(n_303) );
NAND4xp25_ASAP7_75t_L g304 ( .A(n_305), .B(n_339), .C(n_353), .D(n_357), .Y(n_304) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_318), .Y(n_306) );
AND2x4_ASAP7_75t_L g374 ( .A(n_307), .B(n_342), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_307), .B(n_351), .Y(n_375) );
AND2x4_ASAP7_75t_L g377 ( .A(n_307), .B(n_371), .Y(n_377) );
AND2x4_ASAP7_75t_L g425 ( .A(n_307), .B(n_379), .Y(n_425) );
AND2x4_ASAP7_75t_L g432 ( .A(n_307), .B(n_342), .Y(n_432) );
AND2x2_ASAP7_75t_L g434 ( .A(n_307), .B(n_351), .Y(n_434) );
AND2x4_ASAP7_75t_L g437 ( .A(n_307), .B(n_371), .Y(n_437) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_316), .Y(n_307) );
AND2x2_ASAP7_75t_L g356 ( .A(n_308), .B(n_317), .Y(n_356) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g341 ( .A(n_309), .B(n_317), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
NAND2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g315 ( .A(n_311), .Y(n_315) );
INVx3_ASAP7_75t_L g322 ( .A(n_311), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g328 ( .A(n_311), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_311), .Y(n_333) );
INVx1_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_312), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_314), .A2(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g335 ( .A(n_317), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g422 ( .A(n_318), .B(n_341), .Y(n_422) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g379 ( .A(n_319), .Y(n_379) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
AND2x2_ASAP7_75t_L g331 ( .A(n_320), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g342 ( .A(n_320), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
AND2x4_ASAP7_75t_L g371 ( .A(n_320), .B(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_322), .B(n_327), .Y(n_326) );
INVxp67_ASAP7_75t_L g347 ( .A(n_322), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g365 ( .A(n_323), .B(n_346), .C(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g343 ( .A(n_325), .Y(n_343) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_335), .Y(n_330) );
AND2x4_ASAP7_75t_L g414 ( .A(n_331), .B(n_335), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g358 ( .A(n_341), .B(n_351), .Y(n_358) );
AND2x4_ASAP7_75t_L g370 ( .A(n_341), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g378 ( .A(n_341), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g398 ( .A(n_341), .B(n_342), .Y(n_398) );
AND2x2_ASAP7_75t_L g411 ( .A(n_341), .B(n_351), .Y(n_411) );
AND2x2_ASAP7_75t_L g420 ( .A(n_341), .B(n_371), .Y(n_420) );
AND2x2_ASAP7_75t_L g574 ( .A(n_341), .B(n_371), .Y(n_574) );
AND2x4_ASAP7_75t_L g369 ( .A(n_342), .B(n_356), .Y(n_369) );
AND2x4_ASAP7_75t_L g392 ( .A(n_342), .B(n_356), .Y(n_392) );
AND2x4_ASAP7_75t_L g351 ( .A(n_343), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_351), .Y(n_344) );
AND2x4_ASAP7_75t_L g381 ( .A(n_345), .B(n_371), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_345), .B(n_379), .Y(n_382) );
AND2x4_ASAP7_75t_L g405 ( .A(n_345), .B(n_351), .Y(n_405) );
AND2x4_ASAP7_75t_L g428 ( .A(n_345), .B(n_379), .Y(n_428) );
AND2x4_ASAP7_75t_L g440 ( .A(n_345), .B(n_371), .Y(n_440) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x4_ASAP7_75t_L g355 ( .A(n_351), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g626 ( .A(n_351), .B(n_356), .Y(n_626) );
BUFx3_ASAP7_75t_L g585 ( .A(n_354), .Y(n_585) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g401 ( .A(n_355), .Y(n_401) );
BUFx8_ASAP7_75t_SL g462 ( .A(n_355), .Y(n_462) );
INVx2_ASAP7_75t_L g514 ( .A(n_355), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
INVx4_ASAP7_75t_L g496 ( .A(n_361), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_361), .B(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_361), .B(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_361), .B(n_711), .Y(n_710) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g698 ( .A(n_362), .Y(n_698) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_363), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g367 ( .A(n_368), .B(n_373), .C(n_376), .D(n_380), .Y(n_367) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
XNOR2x1_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_416), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_399), .C(n_406), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_393), .B2(n_394), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_390), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_390), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_577) );
INVx4_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx3_ASAP7_75t_L g601 ( .A(n_392), .Y(n_601) );
BUFx3_ASAP7_75t_L g673 ( .A(n_392), .Y(n_673) );
INVx1_ASAP7_75t_L g1012 ( .A(n_392), .Y(n_1012) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g509 ( .A(n_395), .Y(n_509) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g473 ( .A(n_396), .Y(n_473) );
INVx2_ASAP7_75t_L g581 ( .A(n_396), .Y(n_581) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g498 ( .A(n_397), .Y(n_498) );
INVx2_ASAP7_75t_L g717 ( .A(n_397), .Y(n_717) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_398), .Y(n_599) );
BUFx3_ASAP7_75t_L g677 ( .A(n_398), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_399) );
INVx3_ASAP7_75t_L g491 ( .A(n_401), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_403), .A2(n_511), .B1(n_512), .B2(n_515), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_403), .A2(n_583), .B1(n_584), .B2(n_586), .Y(n_582) );
INVx4_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g475 ( .A(n_405), .Y(n_475) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_405), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
INVx3_ASAP7_75t_SL g492 ( .A(n_410), .Y(n_492) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g521 ( .A(n_411), .Y(n_521) );
BUFx3_ASAP7_75t_L g604 ( .A(n_411), .Y(n_604) );
BUFx4f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx5_ASAP7_75t_L g471 ( .A(n_414), .Y(n_471) );
BUFx2_ASAP7_75t_L g591 ( .A(n_414), .Y(n_591) );
BUFx2_ASAP7_75t_L g1051 ( .A(n_414), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_429), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .Y(n_417) );
BUFx8_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_420), .Y(n_451) );
BUFx12f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_422), .Y(n_452) );
BUFx3_ASAP7_75t_L g542 ( .A(n_422), .Y(n_542) );
BUFx6f_ASAP7_75t_L g995 ( .A(n_422), .Y(n_995) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_425), .Y(n_448) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_425), .Y(n_532) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_425), .Y(n_560) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g449 ( .A(n_427), .Y(n_449) );
INVx2_ASAP7_75t_L g535 ( .A(n_427), .Y(n_535) );
INVx5_ASAP7_75t_L g610 ( .A(n_427), .Y(n_610) );
INVx1_ASAP7_75t_L g728 ( .A(n_427), .Y(n_728) );
INVx6_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_428), .Y(n_485) );
NAND2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_435), .Y(n_429) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g458 ( .A(n_432), .Y(n_458) );
BUFx12f_ASAP7_75t_L g547 ( .A(n_432), .Y(n_547) );
BUFx5_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_434), .Y(n_459) );
BUFx3_ASAP7_75t_L g566 ( .A(n_434), .Y(n_566) );
INVx1_ASAP7_75t_L g1037 ( .A(n_434), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx12f_ASAP7_75t_L g454 ( .A(n_437), .Y(n_454) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_437), .Y(n_615) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g455 ( .A(n_439), .Y(n_455) );
INVx1_ASAP7_75t_L g569 ( .A(n_439), .Y(n_569) );
INVx2_ASAP7_75t_L g612 ( .A(n_439), .Y(n_612) );
INVx1_ASAP7_75t_L g647 ( .A(n_439), .Y(n_647) );
INVx4_ASAP7_75t_L g751 ( .A(n_439), .Y(n_751) );
INVx8_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g476 ( .A(n_442), .Y(n_476) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_460), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_450), .C(n_453), .D(n_456), .Y(n_446) );
BUFx3_ASAP7_75t_L g538 ( .A(n_451), .Y(n_538) );
INVx1_ASAP7_75t_L g528 ( .A(n_454), .Y(n_528) );
BUFx12f_ASAP7_75t_L g568 ( .A(n_454), .Y(n_568) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g565 ( .A(n_458), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_458), .A2(n_549), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_L g549 ( .A(n_459), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_469), .C(n_472), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_466), .B(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g523 ( .A(n_468), .Y(n_523) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_468), .Y(n_607) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_468), .Y(n_660) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
INVx2_ASAP7_75t_L g651 ( .A(n_471), .Y(n_651) );
INVx3_ASAP7_75t_L g718 ( .A(n_471), .Y(n_718) );
INVx2_ASAP7_75t_L g1024 ( .A(n_471), .Y(n_1024) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g656 ( .A(n_475), .Y(n_656) );
OA22x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_501), .B2(n_502), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
XNOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .C(n_487), .D(n_488), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_497), .C(n_500), .Y(n_489) );
INVx2_ASAP7_75t_L g1017 ( .A(n_491), .Y(n_1017) );
INVx1_ASAP7_75t_L g589 ( .A(n_492), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_495), .B(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AO22x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_524), .B2(n_550), .Y(n_502) );
NOR4xp25_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .C(n_510), .D(n_516), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
NOR3xp33_ASAP7_75t_SL g551 ( .A(n_506), .B(n_510), .C(n_516), .Y(n_551) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g655 ( .A(n_514), .Y(n_655) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_522), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g709 ( .A(n_520), .Y(n_709) );
INVx2_ASAP7_75t_L g744 ( .A(n_520), .Y(n_744) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g622 ( .A(n_521), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_524), .B(n_551), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .C(n_543), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_532), .Y(n_1001) );
INVx1_ASAP7_75t_L g997 ( .A(n_533), .Y(n_997) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_535), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_541), .A2(n_571), .B1(n_572), .B2(n_575), .Y(n_570) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI22x1_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_545), .B1(n_548), .B2(n_549), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
XOR2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_636), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
XNOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_592), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_576), .Y(n_556) );
NOR3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .C(n_570), .Y(n_557) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
BUFx4f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx4f_ASAP7_75t_L g613 ( .A(n_574), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_582), .C(n_587), .Y(n_576) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_590), .Y(n_587) );
OA22x2_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_617), .B2(n_635), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_596), .B(n_608), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .C(n_600), .D(n_603), .Y(n_596) );
INVx3_ASAP7_75t_L g1022 ( .A(n_599), .Y(n_1022) );
BUFx3_ASAP7_75t_L g713 ( .A(n_602), .Y(n_713) );
INVx3_ASAP7_75t_L g1019 ( .A(n_602), .Y(n_1019) );
INVx1_ASAP7_75t_L g1048 ( .A(n_604), .Y(n_1048) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .C(n_614), .D(n_616), .Y(n_608) );
INVx2_ASAP7_75t_L g635 ( .A(n_617), .Y(n_635) );
AO21x2_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B(n_634), .Y(n_617) );
NOR3xp33_ASAP7_75t_SL g634 ( .A(n_618), .B(n_620), .C(n_629), .Y(n_634) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_629), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .C(n_624), .D(n_625), .Y(n_620) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_622), .Y(n_1009) );
NAND4xp25_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .C(n_632), .D(n_633), .Y(n_629) );
XNOR2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_701), .Y(n_636) );
XNOR2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_662), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
XNOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_661), .Y(n_640) );
NOR4xp75_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .C(n_649), .D(n_653), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_657), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_L g1054 ( .A(n_660), .Y(n_1054) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_684), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_665), .B(n_666), .C(n_668), .D(n_678), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_667), .B(n_679), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_678), .C(n_679), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g682 ( .A(n_671), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .Y(n_671) );
INVx2_ASAP7_75t_L g1044 ( .A(n_673), .Y(n_1044) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XOR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_700), .Y(n_685) );
NOR2xp67_ASAP7_75t_L g686 ( .A(n_687), .B(n_692), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .C(n_690), .D(n_691), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .C(n_695), .D(n_699), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
XOR2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_736), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_719), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .C(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g734 ( .A(n_708), .Y(n_734) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_712), .Y(n_735) );
INVx1_ASAP7_75t_L g731 ( .A(n_714), .Y(n_731) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_717), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g730 ( .A(n_721), .B(n_731), .C(n_732), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_725), .B(n_734), .C(n_735), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_732), .A2(n_787), .B1(n_789), .B2(n_876), .C(n_877), .Y(n_875) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .C(n_748), .D(n_752), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
OA21x2_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
OAI221xp5_ASAP7_75t_SL g755 ( .A1(n_756), .A2(n_981), .B1(n_983), .B2(n_987), .C(n_1025), .Y(n_755) );
O2A1O1Ixp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_848), .B(n_873), .C(n_878), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_782), .B(n_812), .C(n_831), .Y(n_757) );
INVx1_ASAP7_75t_L g932 ( .A(n_758), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_775), .Y(n_758) );
AND2x2_ASAP7_75t_L g829 ( .A(n_759), .B(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g859 ( .A(n_759), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_759), .B(n_874), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_759), .B(n_874), .Y(n_958) );
NOR3xp33_ASAP7_75t_L g977 ( .A(n_759), .B(n_864), .C(n_978), .Y(n_977) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g842 ( .A(n_760), .B(n_775), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_760), .B(n_835), .Y(n_902) );
AND2x2_ASAP7_75t_L g938 ( .A(n_760), .B(n_939), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_760), .B(n_775), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_760), .B(n_867), .Y(n_964) );
AND2x2_ASAP7_75t_L g975 ( .A(n_760), .B(n_776), .Y(n_975) );
AND2x4_ASAP7_75t_L g760 ( .A(n_761), .B(n_768), .Y(n_760) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
AND2x4_ASAP7_75t_L g769 ( .A(n_763), .B(n_770), .Y(n_769) );
AND2x4_ASAP7_75t_L g778 ( .A(n_763), .B(n_765), .Y(n_778) );
AND2x2_ASAP7_75t_L g802 ( .A(n_763), .B(n_765), .Y(n_802) );
AND2x4_ASAP7_75t_L g766 ( .A(n_765), .B(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g779 ( .A(n_765), .B(n_767), .Y(n_779) );
AND2x2_ASAP7_75t_L g803 ( .A(n_765), .B(n_767), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_765), .Y(n_1060) );
INVx2_ASAP7_75t_L g795 ( .A(n_766), .Y(n_795) );
BUFx2_ASAP7_75t_L g982 ( .A(n_766), .Y(n_982) );
AND2x4_ASAP7_75t_L g774 ( .A(n_767), .B(n_770), .Y(n_774) );
AND2x4_ASAP7_75t_L g781 ( .A(n_767), .B(n_770), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_767), .B(n_770), .Y(n_789) );
INVx3_ASAP7_75t_L g787 ( .A(n_769), .Y(n_787) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx3_ASAP7_75t_L g856 ( .A(n_775), .Y(n_856) );
AND2x2_ASAP7_75t_L g860 ( .A(n_775), .B(n_785), .Y(n_860) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g867 ( .A(n_776), .B(n_785), .Y(n_867) );
AND2x2_ASAP7_75t_L g897 ( .A(n_776), .B(n_830), .Y(n_897) );
OR2x2_ASAP7_75t_L g907 ( .A(n_776), .B(n_785), .Y(n_907) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
INVx3_ASAP7_75t_L g793 ( .A(n_778), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_796), .Y(n_782) );
INVx2_ASAP7_75t_L g885 ( .A(n_783), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_SL g942 ( .A1(n_783), .A2(n_814), .B(n_943), .C(n_945), .Y(n_942) );
BUFx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_784), .B(n_833), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_784), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g892 ( .A(n_784), .Y(n_892) );
AND2x2_ASAP7_75t_L g925 ( .A(n_784), .B(n_903), .Y(n_925) );
O2A1O1Ixp33_ASAP7_75t_L g929 ( .A1(n_784), .A2(n_930), .B(n_931), .C(n_932), .Y(n_929) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx3_ASAP7_75t_L g830 ( .A(n_785), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_785), .B(n_819), .Y(n_872) );
OR2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_791), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_789), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_791) );
AND2x2_ASAP7_75t_L g818 ( .A(n_796), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g895 ( .A(n_796), .Y(n_895) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_804), .Y(n_796) );
CKINVDCx6p67_ASAP7_75t_R g815 ( .A(n_797), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_797), .B(n_809), .Y(n_833) );
INVx1_ASAP7_75t_L g840 ( .A(n_797), .Y(n_840) );
AND2x2_ASAP7_75t_L g852 ( .A(n_797), .B(n_853), .Y(n_852) );
OR2x2_ASAP7_75t_L g922 ( .A(n_797), .B(n_809), .Y(n_922) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .Y(n_797) );
INVx1_ASAP7_75t_L g821 ( .A(n_799), .Y(n_821) );
INVx1_ASAP7_75t_L g828 ( .A(n_802), .Y(n_828) );
INVx1_ASAP7_75t_L g826 ( .A(n_803), .Y(n_826) );
AND2x2_ASAP7_75t_SL g948 ( .A(n_804), .B(n_815), .Y(n_948) );
AND2x2_ASAP7_75t_L g955 ( .A(n_804), .B(n_884), .Y(n_955) );
OR2x2_ASAP7_75t_L g961 ( .A(n_804), .B(n_853), .Y(n_961) );
INVxp33_ASAP7_75t_L g968 ( .A(n_804), .Y(n_968) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
INVx1_ASAP7_75t_L g817 ( .A(n_805), .Y(n_817) );
AND2x2_ASAP7_75t_L g845 ( .A(n_805), .B(n_809), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_L g816 ( .A(n_808), .B(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_808), .B(n_839), .Y(n_919) );
OAI222xp33_ASAP7_75t_L g952 ( .A1(n_808), .A2(n_936), .B1(n_941), .B2(n_953), .C1(n_954), .C2(n_956), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g853 ( .A(n_809), .B(n_817), .Y(n_853) );
AOI322xp5_ASAP7_75t_L g901 ( .A1(n_809), .A2(n_856), .A3(n_858), .B1(n_892), .B2(n_902), .C1(n_903), .C2(n_905), .Y(n_901) );
AND2x4_ASAP7_75t_SL g809 ( .A(n_810), .B(n_811), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_818), .B(n_829), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
AND2x2_ASAP7_75t_L g846 ( .A(n_815), .B(n_847), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_815), .B(n_845), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_815), .B(n_819), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_815), .B(n_861), .Y(n_866) );
AND2x2_ASAP7_75t_L g888 ( .A(n_815), .B(n_817), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_815), .A2(n_894), .B1(n_895), .B2(n_896), .Y(n_893) );
AND2x2_ASAP7_75t_L g913 ( .A(n_815), .B(n_853), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_815), .B(n_891), .Y(n_933) );
AND2x2_ASAP7_75t_L g883 ( .A(n_816), .B(n_884), .Y(n_883) );
AND2x2_ASAP7_75t_L g891 ( .A(n_816), .B(n_819), .Y(n_891) );
INVx1_ASAP7_75t_L g906 ( .A(n_816), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_817), .B(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g871 ( .A(n_817), .B(n_839), .Y(n_871) );
INVx1_ASAP7_75t_L g900 ( .A(n_817), .Y(n_900) );
INVx1_ASAP7_75t_L g836 ( .A(n_819), .Y(n_836) );
CKINVDCx6p67_ASAP7_75t_R g847 ( .A(n_819), .Y(n_847) );
AND2x2_ASAP7_75t_L g909 ( .A(n_819), .B(n_830), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_819), .B(n_838), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_819), .B(n_830), .Y(n_973) );
OR2x6_ASAP7_75t_SL g819 ( .A(n_820), .B(n_824), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_830), .B(n_842), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_830), .B(n_859), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_830), .B(n_944), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_830), .B(n_847), .Y(n_979) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_834), .B(n_841), .C(n_843), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_837), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_835), .B(n_852), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_835), .B(n_897), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_835), .B(n_968), .Y(n_967) );
INVx3_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g884 ( .A(n_839), .B(n_847), .Y(n_884) );
AND2x2_ASAP7_75t_L g890 ( .A(n_839), .B(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_839), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_841), .A2(n_874), .B1(n_925), .B2(n_926), .C(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g861 ( .A(n_845), .Y(n_861) );
AND2x2_ASAP7_75t_L g903 ( .A(n_845), .B(n_904), .Y(n_903) );
AND2x2_ASAP7_75t_L g944 ( .A(n_845), .B(n_884), .Y(n_944) );
INVxp67_ASAP7_75t_L g962 ( .A(n_846), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_847), .B(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_847), .B(n_867), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_847), .B(n_897), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_847), .B(n_913), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_847), .B(n_919), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g923 ( .A(n_847), .B(n_907), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_855), .B1(n_857), .B2(n_861), .C(n_862), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_854), .Y(n_850) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_851), .A2(n_963), .B1(n_970), .B2(n_974), .C(n_976), .Y(n_969) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
OAI21xp33_ASAP7_75t_L g920 ( .A1(n_852), .A2(n_921), .B(n_923), .Y(n_920) );
INVx1_ASAP7_75t_L g864 ( .A(n_853), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_853), .B(n_909), .Y(n_908) );
OAI321xp33_ASAP7_75t_L g959 ( .A1(n_854), .A2(n_960), .A3(n_962), .B1(n_963), .B2(n_964), .C(n_965), .Y(n_959) );
INVx3_ASAP7_75t_L g869 ( .A(n_856), .Y(n_869) );
INVx1_ASAP7_75t_L g956 ( .A(n_856), .Y(n_956) );
O2A1O1Ixp33_ASAP7_75t_SL g898 ( .A1(n_857), .A2(n_899), .B(n_901), .C(n_910), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_860), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_858), .B(n_947), .Y(n_946) );
INVx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g894 ( .A(n_860), .Y(n_894) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_860), .B(n_871), .C(n_902), .Y(n_965) );
O2A1O1Ixp33_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_866), .B(n_867), .C(n_868), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
INVx1_ASAP7_75t_L g904 ( .A(n_865), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_866), .B(n_883), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_869), .B(n_910), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_869), .B(n_874), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
CKINVDCx16_ASAP7_75t_R g980 ( .A(n_873), .Y(n_980) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx3_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g910 ( .A(n_875), .Y(n_910) );
NAND5xp2_ASAP7_75t_L g878 ( .A(n_879), .B(n_924), .C(n_937), .D(n_949), .E(n_966), .Y(n_878) );
AOI211xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B(n_898), .C(n_911), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_885), .B1(n_886), .B2(n_887), .C(n_889), .Y(n_881) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_892), .B(n_893), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_892), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g936 ( .A(n_897), .Y(n_936) );
INVx1_ASAP7_75t_L g972 ( .A(n_900), .Y(n_972) );
OAI21xp33_ASAP7_75t_SL g905 ( .A1(n_906), .A2(n_907), .B(n_908), .Y(n_905) );
INVx1_ASAP7_75t_L g939 ( .A(n_907), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_909), .B(n_948), .Y(n_947) );
CKINVDCx16_ASAP7_75t_R g930 ( .A(n_910), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_910), .B(n_936), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_914), .B1(n_915), .B2(n_917), .C(n_920), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_913), .B(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g950 ( .A(n_927), .Y(n_950) );
OAI21xp33_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_933), .B(n_934), .Y(n_928) );
AOI211xp5_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_940), .B(n_942), .C(n_946), .Y(n_937) );
A2O1A1Ixp33_ASAP7_75t_L g966 ( .A1(n_938), .A2(n_967), .B(n_969), .C(n_980), .Y(n_966) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g951 ( .A(n_945), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_951), .B1(n_952), .B2(n_957), .C(n_959), .Y(n_949) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVxp67_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
BUFx6f_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_1006), .Y(n_990) );
NOR3xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_999), .C(n_1003), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
BUFx3_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
NAND2xp5_ASAP7_75t_SL g999 ( .A(n_1000), .B(n_1002), .Y(n_999) );
NOR3xp33_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1015), .C(n_1020), .Y(n_1006) );
NAND2xp5_ASAP7_75t_SL g1007 ( .A(n_1008), .B(n_1010), .Y(n_1007) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1017), .B1(n_1018), .B2(n_1019), .Y(n_1015) );
OAI21xp5_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1022), .B(n_1023), .Y(n_1020) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1028), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1039), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND4xp25_ASAP7_75t_SL g1031 ( .A(n_1032), .B(n_1033), .C(n_1034), .D(n_1038), .Y(n_1031) );
BUFx6f_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .C(n_1046), .Y(n_1040) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
OAI21xp5_ASAP7_75t_SL g1049 ( .A1(n_1050), .A2(n_1052), .B(n_1053), .Y(n_1049) );
INVxp67_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
endmodule