module real_aes_12327_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_18;
wire n_7;
wire n_8;
wire n_10;
INVx1_ASAP7_75t_L g19 ( .A(n_0), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g8 ( .A(n_1), .B(n_9), .Y(n_8) );
INVx3_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_15), .Y(n_14) );
BUFx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
INVx1_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
O2A1O1Ixp33_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_12), .B(n_13), .C(n_17), .Y(n_7) );
INVx2_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_12), .B(n_14), .Y(n_13) );
INVx2_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
endmodule