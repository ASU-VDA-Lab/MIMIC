module fake_jpeg_5592_n_69 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_0),
.B(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_20),
.Y(n_26)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_16),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_27),
.C(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_21),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_31),
.Y(n_40)
);

AOI221xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B1(n_35),
.B2(n_8),
.C(n_11),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_29),
.C(n_32),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_44),
.B(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_15),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_11),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_50),
.B(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_32),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_38),
.B1(n_24),
.B2(n_45),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AO221x1_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_32),
.B1(n_24),
.B2(n_25),
.C(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_25),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_29),
.C(n_38),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_56),
.Y(n_58)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_51),
.B1(n_25),
.B2(n_24),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_14),
.C(n_12),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_7),
.C(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_59),
.B1(n_60),
.B2(n_12),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_6),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_65),
.B(n_10),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_0),
.B(n_3),
.C(n_10),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_14),
.Y(n_69)
);


endmodule