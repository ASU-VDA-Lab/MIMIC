module fake_netlist_1_8199_n_697 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_64), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_41), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_20), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_35), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_32), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_12), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_14), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_61), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_57), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_53), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_80), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_5), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_7), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_36), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_11), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_9), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_8), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_9), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_49), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_78), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_4), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_75), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_26), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_12), .B(n_59), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_74), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_45), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_18), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_23), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_46), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_62), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_14), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_27), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_38), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_51), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_31), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_67), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_30), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_117), .B(n_0), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_112), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_97), .B(n_0), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_94), .B(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_91), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_105), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
CKINVDCx6p67_ASAP7_75t_R g141 ( .A(n_114), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_112), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_121), .B(n_2), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_95), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_128), .B(n_3), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_93), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_90), .B(n_5), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_89), .B(n_6), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_83), .B(n_6), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_86), .B(n_7), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_88), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_103), .Y(n_157) );
CKINVDCx6p67_ASAP7_75t_R g158 ( .A(n_106), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_104), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_110), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_118), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_147), .A2(n_131), .B1(n_143), .B2(n_151), .Y(n_164) );
BUFx10_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_141), .B(n_101), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_133), .B(n_125), .Y(n_172) );
INVx6_ASAP7_75t_L g173 ( .A(n_131), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_141), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_131), .B(n_90), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
AND2x6_ASAP7_75t_L g182 ( .A(n_143), .B(n_96), .Y(n_182) );
AND2x6_ASAP7_75t_L g183 ( .A(n_147), .B(n_96), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_133), .B(n_134), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_134), .A2(n_123), .B1(n_99), .B2(n_119), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_135), .B(n_107), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_135), .B(n_120), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_132), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_144), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_142), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_137), .B(n_120), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_137), .B(n_116), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
AOI22xp33_ASAP7_75t_SL g199 ( .A1(n_138), .A2(n_100), .B1(n_101), .B2(n_115), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_138), .B(n_109), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_132), .B(n_100), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_144), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_149), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_140), .B(n_116), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_129), .B(n_109), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_152), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_146), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_159), .B(n_85), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_157), .B(n_85), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_203), .B(n_192), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_213), .B(n_157), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_217), .B(n_153), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_183), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_187), .A2(n_163), .B(n_162), .C(n_161), .Y(n_225) );
AO22x1_ASAP7_75t_L g226 ( .A1(n_209), .A2(n_158), .B1(n_87), .B2(n_108), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_195), .B(n_157), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_205), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_206), .Y(n_230) );
AND2x2_ASAP7_75t_SL g231 ( .A(n_212), .B(n_158), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_190), .B(n_159), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_167), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_168), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_179), .B(n_154), .Y(n_235) );
NAND2xp33_ASAP7_75t_SL g236 ( .A(n_174), .B(n_108), .Y(n_236) );
BUFx4f_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_190), .B(n_161), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_183), .A2(n_163), .B1(n_162), .B2(n_145), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_183), .A2(n_87), .B1(n_145), .B2(n_102), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_190), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_191), .B(n_163), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
AND2x6_ASAP7_75t_L g246 ( .A(n_164), .B(n_145), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_165), .B(n_162), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_212), .B(n_145), .Y(n_248) );
AND3x1_ASAP7_75t_L g249 ( .A(n_189), .B(n_130), .C(n_155), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_216), .B(n_130), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_165), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_SL g254 ( .A1(n_218), .A2(n_113), .B(n_111), .C(n_98), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_174), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_183), .B(n_84), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_187), .B(n_160), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_195), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_191), .B(n_156), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_173), .Y(n_260) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_218), .B(n_8), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_168), .Y(n_262) );
INVx5_ASAP7_75t_L g263 ( .A(n_178), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g264 ( .A(n_166), .B(n_160), .C(n_156), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_196), .B(n_160), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_178), .A2(n_160), .B1(n_156), .B2(n_152), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_196), .B(n_210), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_210), .B(n_160), .Y(n_268) );
NOR2x1_ASAP7_75t_R g269 ( .A(n_199), .B(n_152), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_179), .B(n_160), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_219), .B(n_156), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_200), .Y(n_272) );
O2A1O1Ixp5_ASAP7_75t_L g273 ( .A1(n_172), .A2(n_156), .B(n_152), .C(n_52), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_179), .B(n_156), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_181), .B(n_152), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_181), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_170), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_181), .B(n_10), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_169), .B(n_50), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_173), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_178), .A2(n_10), .B1(n_11), .B2(n_15), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_244), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_251), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_255), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_246), .A2(n_178), .B1(n_182), .B2(n_173), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_243), .Y(n_286) );
INVxp67_ASAP7_75t_SL g287 ( .A(n_251), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_267), .A2(n_180), .B(n_186), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_241), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_245), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_278), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_237), .A2(n_180), .B1(n_189), .B2(n_200), .Y(n_293) );
OAI21x1_ASAP7_75t_SL g294 ( .A1(n_267), .A2(n_186), .B(n_178), .Y(n_294) );
AO32x1_ASAP7_75t_L g295 ( .A1(n_248), .A2(n_186), .A3(n_194), .B1(n_177), .B2(n_175), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_258), .A2(n_172), .B(n_200), .C(n_170), .Y(n_297) );
BUFx2_ASAP7_75t_SL g298 ( .A(n_263), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_263), .B(n_182), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_223), .B(n_182), .Y(n_300) );
AND2x2_ASAP7_75t_SL g301 ( .A(n_237), .B(n_182), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_220), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_232), .Y(n_303) );
NAND2x1_ASAP7_75t_L g304 ( .A(n_276), .B(n_182), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_246), .A2(n_193), .B1(n_214), .B2(n_211), .Y(n_305) );
INVx6_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_236), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_226), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_251), .B(n_193), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_276), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_229), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_253), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_231), .B(n_15), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_253), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_232), .A2(n_214), .B1(n_211), .B2(n_198), .C(n_215), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_238), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_230), .Y(n_317) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_253), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g319 ( .A1(n_272), .A2(n_215), .B1(n_208), .B2(n_204), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_254), .A2(n_198), .B(n_175), .C(n_177), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g321 ( .A(n_240), .B(n_215), .C(n_208), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_224), .B(n_17), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_256), .B(n_208), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_222), .B(n_215), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_274), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_238), .B(n_194), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_222), .B(n_184), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_294), .A2(n_273), .B(n_279), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_282), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_292), .B(n_246), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_286), .Y(n_333) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_321), .A2(n_261), .B(n_281), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_311), .B(n_246), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_291), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_297), .A2(n_242), .B(n_225), .C(n_259), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_320), .A2(n_278), .B(n_265), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_288), .A2(n_268), .B(n_271), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_291), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_324), .A2(n_249), .B(n_257), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_295), .A2(n_249), .B(n_257), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_311), .B(n_256), .Y(n_343) );
OR2x6_ASAP7_75t_L g344 ( .A(n_299), .B(n_280), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_295), .A2(n_228), .B(n_239), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_247), .B(n_270), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_296), .Y(n_347) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_305), .A2(n_264), .B(n_250), .Y(n_348) );
CKINVDCx14_ASAP7_75t_R g349 ( .A(n_284), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_296), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_290), .B(n_250), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_317), .B(n_235), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_293), .A2(n_260), .B1(n_227), .B2(n_235), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_295), .A2(n_266), .B(n_264), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_295), .A2(n_184), .B(n_262), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_304), .A2(n_277), .B(n_234), .Y(n_357) );
AO31x2_ASAP7_75t_L g358 ( .A1(n_337), .A2(n_325), .A3(n_289), .B(n_275), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_351), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_356), .A2(n_309), .B(n_283), .Y(n_360) );
BUFx6f_ASAP7_75t_SL g361 ( .A(n_331), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_333), .Y(n_362) );
AOI211xp5_ASAP7_75t_L g363 ( .A1(n_330), .A2(n_313), .B(n_328), .C(n_308), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_333), .A2(n_309), .B(n_285), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_343), .A2(n_319), .B1(n_301), .B2(n_308), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_333), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_356), .A2(n_283), .B(n_312), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_351), .B(n_303), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_330), .A2(n_302), .B(n_284), .C(n_307), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_332), .B(n_316), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_342), .A2(n_315), .B(n_327), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_325), .B(n_327), .C(n_323), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_343), .A2(n_301), .B1(n_322), .B2(n_307), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_341), .A2(n_342), .B(n_345), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_331), .B(n_298), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_331), .A2(n_310), .B1(n_322), .B2(n_326), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_332), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_347), .A2(n_322), .B(n_287), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_331), .A2(n_310), .B1(n_326), .B2(n_299), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_336), .B(n_299), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_383), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_362), .B(n_347), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_362), .B(n_336), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_369), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_378), .B(n_350), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_366), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_366), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_365), .A2(n_349), .B1(n_350), .B2(n_355), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_380), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_378), .B(n_355), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_378), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_366), .B(n_357), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_368), .B(n_342), .Y(n_402) );
AND2x4_ASAP7_75t_SL g403 ( .A(n_377), .B(n_344), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_368), .B(n_341), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_367), .B(n_357), .Y(n_405) );
INVx3_ASAP7_75t_SL g406 ( .A(n_377), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_383), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_377), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_367), .B(n_335), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_359), .A2(n_335), .B1(n_353), .B2(n_334), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_374), .A2(n_341), .B(n_345), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_358), .B(n_334), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_360), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_388), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_417), .A2(n_371), .B1(n_363), .B2(n_376), .C(n_375), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_386), .B(n_358), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_417), .B(n_415), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_386), .B(n_358), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_395), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_388), .Y(n_426) );
AOI21xp5_ASAP7_75t_SL g427 ( .A1(n_408), .A2(n_374), .B(n_361), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_415), .B(n_379), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
AO221x1_ASAP7_75t_L g430 ( .A1(n_409), .A2(n_361), .B1(n_283), .B2(n_312), .C(n_314), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_386), .B(n_358), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_389), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_391), .Y(n_433) );
AND2x4_ASAP7_75t_SL g434 ( .A(n_414), .B(n_344), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_390), .B(n_358), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_389), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
NOR2x1p5_ASAP7_75t_L g439 ( .A(n_414), .B(n_352), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_406), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_390), .B(n_373), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_390), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_393), .A2(n_382), .B1(n_352), .B2(n_344), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_385), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_385), .B(n_364), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_385), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_396), .B(n_373), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_406), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_396), .B(n_373), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_393), .B(n_381), .C(n_346), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_406), .A2(n_344), .B1(n_312), .B2(n_314), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_416), .A2(n_334), .B1(n_204), .B2(n_197), .C(n_208), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_409), .A2(n_334), .B1(n_344), .B2(n_348), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_403), .B(n_314), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_411), .A2(n_318), .B(n_338), .C(n_339), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_408), .A2(n_348), .B1(n_338), .B2(n_339), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_414), .B(n_345), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_397), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_403), .A2(n_339), .B1(n_354), .B2(n_356), .C1(n_329), .C2(n_233), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_416), .B(n_348), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g463 ( .A1(n_397), .A2(n_19), .A3(n_21), .B1(n_22), .B2(n_24), .B3(n_28), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_394), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_408), .B(n_329), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_384), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g468 ( .A1(n_403), .A2(n_354), .B1(n_329), .B2(n_204), .C1(n_197), .C2(n_188), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_416), .B(n_348), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_384), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_404), .B(n_354), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_464), .B(n_404), .Y(n_472) );
NOR2x1p5_ASAP7_75t_L g473 ( .A(n_440), .B(n_414), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_419), .Y(n_475) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_456), .B(n_384), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_429), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_464), .B(n_436), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_422), .A2(n_420), .B1(n_428), .B2(n_455), .C(n_436), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_421), .B(n_402), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_421), .B(n_402), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_424), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_424), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_423), .B(n_402), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_463), .B(n_407), .C(n_412), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_432), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_444), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_431), .A2(n_412), .B1(n_410), .B2(n_407), .C(n_413), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_442), .B(n_410), .Y(n_491) );
OR2x4_ASAP7_75t_L g492 ( .A(n_450), .B(n_413), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_427), .A2(n_407), .B(n_400), .Y(n_493) );
OAI21x1_ASAP7_75t_L g494 ( .A1(n_458), .A2(n_418), .B(n_391), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_440), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_446), .B(n_407), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_423), .B(n_410), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_426), .B(n_399), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_426), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_462), .B(n_410), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_462), .B(n_410), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_469), .B(n_418), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_441), .B(n_399), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_437), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_451), .B(n_391), .C(n_392), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_437), .B(n_400), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_466), .B(n_405), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_460), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_466), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_439), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_467), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_466), .B(n_433), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_456), .B(n_405), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_469), .B(n_401), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_461), .B(n_413), .C(n_405), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_438), .B(n_401), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_441), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_453), .Y(n_520) );
INVx6_ASAP7_75t_L g521 ( .A(n_448), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_471), .B(n_418), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_471), .B(n_405), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_447), .B(n_405), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_449), .B(n_394), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_453), .B(n_413), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_443), .A2(n_392), .B1(n_398), .B2(n_413), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_470), .B(n_392), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_465), .B(n_413), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_434), .Y(n_531) );
NAND5xp2_ASAP7_75t_SL g532 ( .A(n_454), .B(n_29), .C(n_33), .D(n_34), .E(n_37), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_445), .B(n_398), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_433), .B(n_413), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_433), .B(n_398), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_479), .B(n_459), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_501), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_480), .A2(n_430), .B1(n_434), .B2(n_435), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_523), .B(n_435), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_479), .B(n_435), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_523), .B(n_468), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_484), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_481), .B(n_398), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_519), .B(n_427), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_481), .B(n_398), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_474), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_512), .B(n_457), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_473), .B(n_430), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_477), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_510), .B(n_452), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_521), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_482), .B(n_188), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_488), .B(n_188), .Y(n_555) );
NOR2xp67_ASAP7_75t_SL g556 ( .A(n_521), .B(n_306), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_509), .B(n_43), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_483), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_496), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_482), .B(n_188), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
NAND2xp67_ASAP7_75t_L g562 ( .A(n_535), .B(n_44), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_485), .B(n_47), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_485), .B(n_176), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_501), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_502), .B(n_176), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_513), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_495), .B(n_48), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_521), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_502), .B(n_176), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_506), .Y(n_571) );
NOR2x1p5_ASAP7_75t_SL g572 ( .A(n_518), .B(n_54), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_472), .B(n_176), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_484), .B(n_55), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_505), .B(n_56), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_515), .A2(n_204), .B1(n_197), .B2(n_306), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_503), .B(n_499), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_475), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_475), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_503), .B(n_197), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_490), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_490), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_509), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_472), .B(n_58), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_520), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_505), .B(n_60), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_499), .B(n_63), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_524), .B(n_65), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_524), .B(n_66), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_504), .B(n_68), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_498), .B(n_69), .Y(n_592) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_498), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_558), .Y(n_594) );
OAI211xp5_ASAP7_75t_L g595 ( .A1(n_538), .A2(n_515), .B(n_527), .C(n_531), .Y(n_595) );
INVxp67_ASAP7_75t_SL g596 ( .A(n_558), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_542), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_548), .B(n_486), .C(n_517), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_549), .A2(n_492), .B(n_493), .Y(n_599) );
OAI21xp5_ASAP7_75t_SL g600 ( .A1(n_549), .A2(n_476), .B(n_509), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_541), .A2(n_514), .B1(n_511), .B2(n_528), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_541), .A2(n_514), .B1(n_511), .B2(n_528), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_546), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_567), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_548), .A2(n_590), .B1(n_544), .B2(n_589), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_583), .B(n_542), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_556), .B(n_507), .C(n_489), .Y(n_607) );
BUFx2_ASAP7_75t_L g608 ( .A(n_593), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_547), .Y(n_609) );
AOI222xp33_ASAP7_75t_L g610 ( .A1(n_551), .A2(n_497), .B1(n_504), .B2(n_522), .C1(n_525), .C2(n_511), .Y(n_610) );
INVx3_ASAP7_75t_L g611 ( .A(n_583), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_550), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_590), .A2(n_476), .B1(n_491), .B2(n_492), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_577), .B(n_522), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_563), .A2(n_514), .B1(n_535), .B2(n_525), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_577), .B(n_533), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_552), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_557), .A2(n_491), .B1(n_500), .B2(n_508), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_553), .Y(n_619) );
NOR2xp33_ASAP7_75t_SL g620 ( .A(n_569), .B(n_532), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_568), .A2(n_534), .B1(n_529), .B2(n_520), .C(n_526), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_559), .A2(n_530), .B1(n_526), .B2(n_534), .C(n_529), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_571), .Y(n_624) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_555), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_536), .B(n_530), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_578), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_568), .A2(n_306), .B1(n_494), .B2(n_73), .C(n_76), .Y(n_628) );
INVx3_ASAP7_75t_SL g629 ( .A(n_553), .Y(n_629) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_583), .A2(n_494), .B(n_71), .C(n_77), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_557), .A2(n_592), .B(n_574), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_540), .B(n_70), .Y(n_632) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_588), .A2(n_79), .B(n_306), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_539), .B(n_575), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_626), .B(n_545), .Y(n_635) );
NAND2xp33_ASAP7_75t_L g636 ( .A(n_629), .B(n_591), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_608), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_601), .B(n_539), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_614), .B(n_545), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_603), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_609), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_610), .B(n_582), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_619), .B(n_562), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_623), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_627), .B(n_579), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_612), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_597), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_617), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_624), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_606), .B(n_543), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_604), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_600), .A2(n_586), .B1(n_576), .B2(n_557), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_598), .A2(n_561), .B1(n_565), .B2(n_560), .C(n_573), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_598), .A2(n_591), .B1(n_584), .B2(n_587), .C(n_554), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_596), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_622), .B(n_581), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_616), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_625), .Y(n_659) );
OAI22xp33_ASAP7_75t_SL g660 ( .A1(n_599), .A2(n_592), .B1(n_574), .B2(n_564), .Y(n_660) );
AOI221x1_ASAP7_75t_L g661 ( .A1(n_643), .A2(n_607), .B1(n_631), .B2(n_606), .C(n_613), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_646), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_646), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_636), .A2(n_607), .B1(n_602), .B2(n_605), .C(n_595), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_660), .A2(n_621), .B(n_618), .C(n_620), .Y(n_665) );
NAND4xp75_ASAP7_75t_L g666 ( .A(n_643), .B(n_572), .C(n_632), .D(n_615), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_659), .B(n_634), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_638), .Y(n_668) );
OAI311xp33_ASAP7_75t_L g669 ( .A1(n_655), .A2(n_628), .A3(n_611), .B1(n_580), .C1(n_554), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_648), .A2(n_611), .B1(n_630), .B2(n_580), .Y(n_670) );
OAI21xp33_ASAP7_75t_SL g671 ( .A1(n_651), .A2(n_566), .B(n_570), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_655), .A2(n_633), .B(n_566), .C(n_570), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_653), .A2(n_537), .B1(n_585), .B2(n_639), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_637), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_649), .Y(n_675) );
AND3x1_ASAP7_75t_L g676 ( .A(n_665), .B(n_644), .C(n_654), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_664), .A2(n_657), .B(n_656), .C(n_652), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_661), .A2(n_657), .B(n_642), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_671), .A2(n_664), .B(n_673), .C(n_668), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_674), .B(n_641), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_670), .B(n_645), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_675), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_662), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_680), .Y(n_684) );
NOR2xp33_ASAP7_75t_R g685 ( .A(n_680), .B(n_667), .Y(n_685) );
NOR3xp33_ASAP7_75t_SL g686 ( .A(n_679), .B(n_666), .C(n_669), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_677), .B(n_678), .C(n_681), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_684), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_687), .B(n_672), .C(n_683), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_685), .Y(n_690) );
NAND2x1_ASAP7_75t_L g691 ( .A(n_690), .B(n_686), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_688), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_691), .A2(n_676), .B1(n_689), .B2(n_682), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_693), .B(n_692), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_663), .B1(n_647), .B2(n_650), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_695), .B(n_658), .C(n_640), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_537), .B1(n_635), .B2(n_585), .Y(n_697) );
endmodule