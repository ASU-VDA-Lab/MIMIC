module fake_jpeg_6214_n_133 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_28),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_1),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_2),
.C(n_3),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_14),
.C(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_26),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_41),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_25),
.B1(n_22),
.B2(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_61),
.B1(n_40),
.B2(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_33),
.C(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_26),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_36),
.B1(n_45),
.B2(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_48),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_53),
.B(n_49),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_50),
.C(n_60),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_88),
.C(n_68),
.Y(n_91)
);

AOI21x1_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_26),
.B(n_16),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_45),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_70),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_57),
.B1(n_17),
.B2(n_26),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_17),
.B1(n_26),
.B2(n_16),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_80),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_94),
.C(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_67),
.B(n_33),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_96),
.B(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_77),
.C(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_99),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

XOR2x2_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_33),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_84),
.B(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_101),
.B1(n_103),
.B2(n_107),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_107),
.C(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_110),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_27),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_4),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_16),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

AOI31xp33_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_112),
.A3(n_116),
.B(n_16),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_11),
.B(n_8),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.C(n_123),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_6),
.B(n_9),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_127),
.B(n_10),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_10),
.C(n_11),
.Y(n_132)
);


endmodule