module fake_jpeg_1718_n_563 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_563);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_563;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_98),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_65),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_19),
.B(n_18),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_66),
.B(n_123),
.Y(n_210)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_71),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_90),
.Y(n_135)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_76),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_77),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_79),
.Y(n_207)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_81),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_84),
.Y(n_208)
);

CKINVDCx9p33_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_33),
.B(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

CKINVDCx9p33_ASAP7_75t_R g97 ( 
.A(n_28),
.Y(n_97)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_32),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_103),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_100),
.Y(n_196)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_32),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_108),
.Y(n_150)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_125),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_50),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_20),
.B1(n_54),
.B2(n_55),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_136),
.A2(n_168),
.B1(n_184),
.B2(n_185),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_66),
.B(n_39),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_141),
.B(n_153),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_55),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_149),
.B(n_166),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_67),
.B(n_39),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_65),
.B(n_49),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_155),
.B(n_159),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_49),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_59),
.B(n_22),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_162),
.B(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_22),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_71),
.A2(n_56),
.B1(n_24),
.B2(n_27),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_24),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_57),
.B1(n_45),
.B2(n_53),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_112),
.A2(n_57),
.B1(n_45),
.B2(n_53),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_34),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_114),
.A2(n_27),
.B1(n_48),
.B2(n_31),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_188),
.A2(n_191),
.B1(n_212),
.B2(n_213),
.Y(n_274)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_73),
.Y(n_190)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_71),
.A2(n_56),
.B1(n_48),
.B2(n_31),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_63),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_192),
.B(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_78),
.B(n_34),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_123),
.B(n_54),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_77),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_204),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_88),
.A2(n_20),
.B1(n_47),
.B2(n_57),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_203),
.A2(n_16),
.B(n_3),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_81),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_92),
.A2(n_56),
.B1(n_47),
.B2(n_52),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_47),
.B1(n_52),
.B2(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_216),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_128),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_218),
.B(n_223),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_136),
.A2(n_110),
.B1(n_82),
.B2(n_106),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_219),
.A2(n_237),
.B1(n_288),
.B2(n_211),
.Y(n_314)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_210),
.A2(n_89),
.B1(n_104),
.B2(n_72),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_165),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_108),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_224),
.B(n_235),
.C(n_240),
.Y(n_327)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_129),
.A2(n_72),
.B1(n_107),
.B2(n_102),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_229),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_230),
.B(n_236),
.Y(n_339)
);

INVx6_ASAP7_75t_SL g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_232),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_139),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_234),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_131),
.B(n_108),
.C(n_91),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_203),
.A2(n_83),
.B1(n_47),
.B2(n_52),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_140),
.Y(n_239)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_239),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_145),
.B(n_52),
.C(n_3),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_241),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_130),
.B(n_16),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_242),
.A2(n_256),
.B(n_275),
.Y(n_329)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_244),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_150),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_147),
.B(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_248),
.B(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_154),
.Y(n_249)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_181),
.B(n_132),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_SL g291 ( 
.A(n_252),
.B(n_208),
.C(n_143),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_157),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_254),
.Y(n_292)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_158),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_262),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_134),
.B(n_16),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_149),
.B(n_1),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_257),
.B(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_135),
.B(n_3),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_259),
.B(n_281),
.Y(n_300)
);

BUFx4f_ASAP7_75t_SL g262 ( 
.A(n_187),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_129),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_264),
.A2(n_269),
.B1(n_286),
.B2(n_287),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_127),
.B(n_6),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_148),
.B(n_6),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_266),
.B(n_270),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_172),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_272),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_209),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_268),
.A2(n_189),
.B1(n_248),
.B2(n_283),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_208),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_175),
.B(n_10),
.Y(n_270)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_174),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_142),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_201),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_273),
.A2(n_268),
.B1(n_234),
.B2(n_220),
.Y(n_340)
);

OR2x2_ASAP7_75t_SL g275 ( 
.A(n_201),
.B(n_12),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_277),
.Y(n_310)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_165),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_137),
.A2(n_12),
.B(n_13),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_284),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_13),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_144),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_160),
.B(n_16),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_157),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_171),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_160),
.B(n_142),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_212),
.A2(n_168),
.B1(n_191),
.B2(n_167),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g381 ( 
.A(n_291),
.B(n_330),
.C(n_335),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_293),
.B(n_251),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_257),
.A2(n_169),
.B(n_151),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g361 ( 
.A1(n_294),
.A2(n_329),
.B(n_256),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_238),
.A2(n_167),
.B1(n_199),
.B2(n_198),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_295),
.A2(n_318),
.B1(n_321),
.B2(n_334),
.Y(n_364)
);

AO22x2_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_178),
.B1(n_171),
.B2(n_143),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_231),
.A2(n_178),
.B1(n_206),
.B2(n_174),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_307),
.A2(n_311),
.B1(n_295),
.B2(n_321),
.Y(n_369)
);

OA22x2_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_302),
.B1(n_326),
.B2(n_299),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_245),
.A2(n_196),
.B(n_197),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_253),
.B(n_285),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_258),
.A2(n_206),
.B1(n_199),
.B2(n_198),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_250),
.A2(n_183),
.B1(n_146),
.B2(n_205),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_260),
.A2(n_187),
.B1(n_189),
.B2(n_176),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_328),
.A2(n_340),
.B1(n_343),
.B2(n_215),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_252),
.A2(n_187),
.B(n_189),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_237),
.A2(n_183),
.B1(n_172),
.B2(n_176),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_341),
.B1(n_242),
.B2(n_240),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_247),
.A2(n_256),
.B(n_217),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_224),
.B(n_249),
.C(n_239),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_286),
.C(n_226),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_235),
.A2(n_266),
.B1(n_270),
.B2(n_288),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_232),
.A2(n_282),
.B1(n_280),
.B2(n_255),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_344),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_243),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_354),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_346),
.A2(n_348),
.B1(n_358),
.B2(n_383),
.Y(n_392)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_312),
.Y(n_347)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_314),
.A2(n_242),
.B1(n_278),
.B2(n_265),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_298),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_349),
.B(n_377),
.Y(n_414)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_352),
.A2(n_369),
.B(n_376),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_361),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_339),
.Y(n_354)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_324),
.B(n_275),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_357),
.B(n_362),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_306),
.A2(n_246),
.B1(n_271),
.B2(n_227),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_382),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_263),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_306),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_365),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_256),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_330),
.A2(n_216),
.B(n_225),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_367),
.A2(n_303),
.B(n_297),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_261),
.C(n_221),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_289),
.C(n_290),
.Y(n_391)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_373),
.C(n_374),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_327),
.B(n_254),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_229),
.C(n_241),
.Y(n_374)
);

AOI22x1_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_244),
.B1(n_277),
.B2(n_262),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_355),
.B1(n_369),
.B2(n_383),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_302),
.A2(n_233),
.B1(n_262),
.B2(n_299),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_324),
.B(n_335),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_322),
.B(n_300),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_380),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_293),
.B(n_334),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_318),
.C(n_290),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_311),
.B(n_294),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_313),
.B(n_292),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_297),
.A2(n_333),
.B1(n_300),
.B2(n_315),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_316),
.B(n_310),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_384),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_296),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_385),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_388),
.A2(n_348),
.B1(n_375),
.B2(n_363),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_391),
.B(n_353),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_396),
.C(n_397),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_325),
.C(n_289),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_336),
.C(n_331),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_399),
.A2(n_409),
.B(n_379),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_355),
.A2(n_297),
.B1(n_315),
.B2(n_303),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_399),
.B(n_409),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_336),
.C(n_331),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_301),
.C(n_305),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_367),
.A2(n_297),
.B(n_317),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_346),
.A2(n_319),
.B1(n_338),
.B2(n_309),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_410),
.A2(n_413),
.B1(n_356),
.B2(n_317),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_355),
.A2(n_319),
.B1(n_338),
.B2(n_309),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_364),
.A2(n_317),
.B1(n_305),
.B2(n_301),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_401),
.B1(n_394),
.B2(n_388),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_380),
.A2(n_384),
.B(n_381),
.C(n_353),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_357),
.B(n_375),
.C(n_365),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_372),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_427),
.C(n_434),
.Y(n_469)
);

AO21x1_ASAP7_75t_L g456 ( 
.A1(n_421),
.A2(n_430),
.B(n_440),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_422),
.A2(n_447),
.B1(n_448),
.B2(n_407),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_349),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_382),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_425),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_351),
.Y(n_426)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_377),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_347),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g431 ( 
.A(n_418),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_431),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_358),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_433),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_389),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_396),
.B(n_352),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_366),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_437),
.Y(n_470)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_414),
.B(n_359),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_438),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_444),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_371),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_445),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_364),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_449),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_443),
.B(n_398),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_397),
.B(n_353),
.C(n_350),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_446),
.A2(n_415),
.B1(n_413),
.B2(n_401),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_386),
.B(n_323),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_368),
.Y(n_449)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_451),
.B(n_461),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_422),
.A2(n_392),
.B1(n_398),
.B2(n_410),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_452),
.A2(n_460),
.B1(n_465),
.B2(n_472),
.Y(n_477)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

AO22x1_ASAP7_75t_L g455 ( 
.A1(n_431),
.A2(n_398),
.B1(n_394),
.B2(n_416),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_473),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_448),
.A2(n_392),
.B1(n_406),
.B2(n_393),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_402),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_395),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_469),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_440),
.A2(n_393),
.B1(n_416),
.B2(n_419),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_433),
.A2(n_419),
.B1(n_405),
.B2(n_403),
.Y(n_468)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_431),
.A2(n_411),
.B1(n_387),
.B2(n_403),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_426),
.A2(n_411),
.B1(n_368),
.B2(n_323),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_444),
.B1(n_436),
.B2(n_446),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_475),
.A2(n_449),
.B1(n_434),
.B2(n_435),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_454),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_494),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_482),
.A2(n_489),
.B1(n_495),
.B2(n_463),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_471),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_483),
.B(n_487),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_427),
.C(n_439),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_484),
.B(n_492),
.C(n_490),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_456),
.A2(n_421),
.B(n_430),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_456),
.A2(n_428),
.B(n_443),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_486),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_465),
.A2(n_432),
.B(n_441),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_445),
.Y(n_488)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_488),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_452),
.A2(n_424),
.B1(n_460),
.B2(n_476),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_464),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_457),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_457),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_463),
.B(n_451),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_497),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_470),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_476),
.A2(n_455),
.B1(n_475),
.B2(n_466),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_458),
.Y(n_496)
);

INVx13_ASAP7_75t_L g507 ( 
.A(n_496),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_462),
.A2(n_455),
.B(n_472),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_501),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_491),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_477),
.A2(n_466),
.B1(n_462),
.B2(n_467),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_478),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_459),
.Y(n_509)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_509),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_511),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_470),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_498),
.B(n_474),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_512),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_467),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_505),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_520),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_480),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_522),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_491),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_521),
.B(n_527),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_510),
.C(n_482),
.Y(n_522)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_524),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_493),
.C(n_480),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_525),
.B(n_499),
.C(n_513),
.Y(n_536)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_509),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_526),
.A2(n_479),
.B1(n_506),
.B2(n_502),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_499),
.A2(n_497),
.B(n_485),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_523),
.B(n_508),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_529),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_523),
.B(n_481),
.C(n_504),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_535),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_518),
.A2(n_481),
.B1(n_506),
.B2(n_502),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_536),
.B(n_530),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_477),
.C(n_489),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_538),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_495),
.C(n_478),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_541),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_522),
.C(n_525),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_520),
.C(n_515),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_545),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_527),
.Y(n_543)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_543),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_531),
.B(n_516),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_524),
.C(n_487),
.Y(n_547)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_547),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g548 ( 
.A(n_539),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_496),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_540),
.A2(n_546),
.B(n_544),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_553),
.A2(n_544),
.B(n_534),
.Y(n_554)
);

AOI21xp33_ASAP7_75t_L g558 ( 
.A1(n_554),
.A2(n_555),
.B(n_556),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_552),
.B(n_537),
.C(n_494),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_551),
.B(n_486),
.C(n_496),
.Y(n_557)
);

OAI221xp5_ASAP7_75t_L g559 ( 
.A1(n_557),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.C(n_507),
.Y(n_559)
);

O2A1O1Ixp33_ASAP7_75t_SL g560 ( 
.A1(n_559),
.A2(n_458),
.B(n_507),
.C(n_453),
.Y(n_560)
);

BUFx24_ASAP7_75t_SL g561 ( 
.A(n_560),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_561),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_558),
.Y(n_563)
);


endmodule