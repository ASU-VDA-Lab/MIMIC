module real_aes_3820_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_17;
wire n_13;
wire n_6;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_5;
wire n_15;
wire n_9;
wire n_20;
wire n_18;
wire n_7;
wire n_8;
wire n_10;
INVx2_ASAP7_75t_L g6 ( .A(n_0), .Y(n_6) );
AND2x4_ASAP7_75t_L g5 ( .A(n_1), .B(n_6), .Y(n_5) );
INVx1_ASAP7_75t_L g19 ( .A(n_1), .Y(n_19) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
AND2x4_ASAP7_75t_L g12 ( .A(n_2), .B(n_13), .Y(n_12) );
AND2x4_ASAP7_75t_L g20 ( .A(n_2), .B(n_3), .Y(n_20) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
AOI211xp5_ASAP7_75t_SL g4 ( .A1(n_5), .A2(n_7), .B(n_9), .C(n_14), .Y(n_4) );
AND2x4_ASAP7_75t_L g11 ( .A(n_5), .B(n_12), .Y(n_11) );
AND2x2_ASAP7_75t_L g18 ( .A(n_6), .B(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
INVx2_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx2_ASAP7_75t_SL g10 ( .A(n_11), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_18), .B(n_20), .Y(n_17) );
endmodule