module fake_jpeg_3645_n_546 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_546);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_65),
.Y(n_107)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g148 ( 
.A(n_54),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_69),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_88),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_61),
.A2(n_67),
.B1(n_43),
.B2(n_42),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_19),
.B(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_18),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_2),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_94),
.Y(n_136)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_87),
.Y(n_129)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_28),
.B(n_4),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_100),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_102),
.Y(n_159)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_51),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_104),
.B(n_163),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_28),
.B1(n_39),
.B2(n_37),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_111),
.A2(n_139),
.B1(n_150),
.B2(n_73),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_26),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_112),
.B(n_115),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_50),
.B1(n_37),
.B2(n_39),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_113),
.A2(n_120),
.B1(n_124),
.B2(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_26),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_52),
.A2(n_25),
.B1(n_23),
.B2(n_31),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_118),
.A2(n_137),
.B1(n_146),
.B2(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_50),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_96),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_102),
.B1(n_95),
.B2(n_92),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_55),
.A2(n_46),
.B1(n_23),
.B2(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_26),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_127),
.B(n_143),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_62),
.A2(n_25),
.B1(n_46),
.B2(n_35),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_59),
.A2(n_46),
.B1(n_35),
.B2(n_31),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_60),
.A2(n_35),
.B1(n_25),
.B2(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_40),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_75),
.A2(n_49),
.B1(n_48),
.B2(n_36),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_66),
.A2(n_49),
.B1(n_48),
.B2(n_24),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_71),
.B(n_43),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_154),
.B(n_7),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_85),
.A2(n_48),
.B1(n_40),
.B2(n_43),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_73),
.B1(n_44),
.B2(n_33),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_88),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_109),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_58),
.A2(n_42),
.B1(n_36),
.B2(n_32),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_54),
.A2(n_32),
.B(n_30),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_77),
.A2(n_32),
.B1(n_30),
.B2(n_44),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_103),
.B1(n_101),
.B2(n_99),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_167),
.A2(n_181),
.B1(n_189),
.B2(n_199),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_171),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_172),
.B(n_180),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_97),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_173),
.B(n_187),
.C(n_156),
.Y(n_242)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_177),
.Y(n_227)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_83),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_91),
.B1(n_81),
.B2(n_96),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_70),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_182),
.B(n_184),
.Y(n_240)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_204),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_109),
.B(n_70),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_112),
.A2(n_30),
.B1(n_44),
.B2(n_33),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_190),
.B(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_192),
.A2(n_203),
.B1(n_212),
.B2(n_17),
.Y(n_273)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_142),
.B1(n_130),
.B2(n_144),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_123),
.Y(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_44),
.B1(n_33),
.B2(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_200),
.B(n_202),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_114),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_201),
.B(n_209),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_133),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_113),
.A2(n_44),
.B1(n_33),
.B2(n_7),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_128),
.B(n_5),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_205),
.B(n_206),
.Y(n_278)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_208),
.Y(n_279)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_138),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_135),
.B(n_6),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_210),
.B(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_140),
.A2(n_44),
.B1(n_33),
.B2(n_9),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_213),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_215),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_114),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_122),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_224),
.B1(n_126),
.B2(n_162),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_110),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_145),
.B(n_8),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_220),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_138),
.Y(n_220)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_223),
.Y(n_262)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_122),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_224)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_131),
.B1(n_158),
.B2(n_145),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_231),
.A2(n_257),
.B1(n_267),
.B2(n_217),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_235),
.A2(n_236),
.B1(n_253),
.B2(n_256),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_126),
.B1(n_162),
.B2(n_116),
.Y(n_236)
);

NAND2x1p5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_179),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_237),
.B(n_273),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_242),
.B(n_207),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_SL g285 ( 
.A1(n_243),
.A2(n_245),
.B(n_263),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_169),
.B(n_105),
.C(n_156),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_268),
.C(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_142),
.B(n_130),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_245),
.A2(n_263),
.B(n_249),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_105),
.B(n_152),
.C(n_121),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_246),
.B(n_189),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_185),
.A2(n_116),
.B1(n_165),
.B2(n_152),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_175),
.A2(n_165),
.B1(n_153),
.B2(n_131),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_197),
.A2(n_153),
.B1(n_11),
.B2(n_12),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_222),
.A2(n_194),
.B(n_166),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_173),
.B(n_10),
.CI(n_11),
.CON(n_266),
.SN(n_266)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_203),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_222),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_182),
.B(n_12),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_14),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_196),
.A2(n_17),
.B(n_15),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_209),
.B(n_205),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_190),
.B(n_15),
.C(n_16),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_276),
.C(n_220),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_187),
.B(n_15),
.C(n_16),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_193),
.B(n_16),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_224),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_280),
.B(n_287),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_184),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g365 ( 
.A1(n_283),
.A2(n_292),
.B(n_296),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_300),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_295),
.B1(n_303),
.B2(n_305),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_286),
.A2(n_304),
.B1(n_314),
.B2(n_318),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_227),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_178),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_288),
.B(n_294),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_297),
.Y(n_363)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_174),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_239),
.A2(n_192),
.B1(n_195),
.B2(n_200),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_261),
.B(n_230),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_240),
.B(n_168),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_187),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_SL g302 ( 
.A1(n_239),
.A2(n_181),
.B(n_199),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_302),
.A2(n_276),
.B(n_253),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_228),
.A2(n_167),
.B1(n_198),
.B2(n_183),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_216),
.B1(n_201),
.B2(n_226),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_228),
.A2(n_218),
.B1(n_176),
.B2(n_171),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_238),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_313),
.Y(n_357)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_322),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_237),
.B(n_170),
.C(n_208),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_319),
.C(n_321),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_206),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_310),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_311),
.A2(n_325),
.B(n_327),
.Y(n_343)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_176),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_264),
.A2(n_218),
.B1(n_202),
.B2(n_213),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_232),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_316),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_246),
.A2(n_177),
.B(n_225),
.C(n_223),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_317),
.A2(n_229),
.B(n_233),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_252),
.A2(n_202),
.B1(n_221),
.B2(n_207),
.Y(n_318)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_242),
.B(n_207),
.C(n_17),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_230),
.B(n_254),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_231),
.Y(n_323)
);

NAND2x1_ASAP7_75t_SL g336 ( 
.A(n_323),
.B(n_243),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_265),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_234),
.C(n_247),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_249),
.A2(n_248),
.B(n_265),
.Y(n_325)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_342),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_235),
.B1(n_256),
.B2(n_267),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_335),
.A2(n_347),
.B1(n_355),
.B2(n_286),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_336),
.A2(n_337),
.B(n_340),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_259),
.B(n_277),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_346),
.Y(n_394)
);

XOR2x2_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_268),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_289),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_318),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_257),
.B1(n_236),
.B2(n_243),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_309),
.B(n_266),
.CI(n_244),
.CON(n_349),
.SN(n_349)
);

AOI21xp33_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_298),
.B(n_303),
.Y(n_396)
);

OA22x2_ASAP7_75t_L g350 ( 
.A1(n_307),
.A2(n_243),
.B1(n_229),
.B2(n_269),
.Y(n_350)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_301),
.A2(n_266),
.B1(n_269),
.B2(n_250),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_321),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_360),
.A2(n_362),
.B(n_274),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_311),
.A2(n_278),
.B(n_279),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_270),
.C(n_272),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_289),
.C(n_325),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_405),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_377),
.C(n_379),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_324),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_287),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_380),
.B(n_381),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_368),
.B(n_291),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_339),
.B(n_308),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_383),
.B(n_386),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_357),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_401),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_328),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_387),
.C(n_389),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_368),
.B(n_306),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_315),
.C(n_299),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_343),
.A2(n_317),
.B(n_323),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_393),
.B(n_397),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_295),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_337),
.B1(n_338),
.B2(n_367),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_323),
.C(n_274),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_395),
.C(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_343),
.A2(n_283),
.B(n_284),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_314),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g422 ( 
.A(n_396),
.B(n_355),
.CI(n_349),
.CON(n_422),
.SN(n_422)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_365),
.B(n_250),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_403),
.Y(n_437)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_345),
.B(n_234),
.C(n_247),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_320),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_360),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_407),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_329),
.B(n_305),
.C(n_282),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_408),
.A2(n_409),
.B1(n_415),
.B2(n_417),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_384),
.B1(n_392),
.B2(n_394),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_372),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_410),
.B(n_427),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_374),
.A2(n_332),
.B1(n_347),
.B2(n_330),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_394),
.A2(n_332),
.B1(n_329),
.B2(n_338),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_393),
.A2(n_334),
.B1(n_335),
.B2(n_346),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_418),
.A2(n_425),
.B1(n_358),
.B2(n_354),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

INVx3_ASAP7_75t_SL g460 ( 
.A(n_419),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_404),
.A2(n_334),
.B1(n_369),
.B2(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

AOI221xp5_ASAP7_75t_L g444 ( 
.A1(n_422),
.A2(n_376),
.B1(n_373),
.B2(n_375),
.C(n_385),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_336),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_372),
.A2(n_361),
.B1(n_352),
.B2(n_340),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_361),
.B1(n_356),
.B2(n_336),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_405),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_387),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_429),
.B(n_434),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_344),
.B1(n_350),
.B2(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_391),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_378),
.A2(n_350),
.B1(n_359),
.B2(n_342),
.Y(n_438)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_375),
.A2(n_350),
.B1(n_349),
.B2(n_354),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_402),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_440),
.B(n_445),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_377),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_456),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_444),
.A2(n_459),
.B1(n_411),
.B2(n_422),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_379),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_406),
.Y(n_446)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_446),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_413),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_447),
.B(n_418),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_378),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_448),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_397),
.B(n_399),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_414),
.B(n_424),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_401),
.C(n_398),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_461),
.C(n_420),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_423),
.B(n_382),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_454),
.B(n_426),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_382),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_455),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_358),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_428),
.B(n_353),
.C(n_331),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_353),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_428),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_331),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_433),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_478),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_476),
.C(n_479),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_472),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_471),
.A2(n_474),
.B(n_453),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_449),
.A2(n_424),
.B(n_413),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_439),
.C(n_438),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_461),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_432),
.C(n_408),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_443),
.B(n_425),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_483),
.Y(n_495)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

OA21x2_ASAP7_75t_SL g483 ( 
.A1(n_441),
.A2(n_422),
.B(n_411),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_451),
.Y(n_497)
);

A2O1A1O1Ixp25_ASAP7_75t_L g486 ( 
.A1(n_458),
.A2(n_413),
.B(n_415),
.C(n_421),
.D(n_430),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_486),
.A2(n_457),
.B(n_455),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_431),
.B1(n_430),
.B2(n_419),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_465),
.B1(n_459),
.B2(n_466),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_494),
.B1(n_504),
.B2(n_505),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_446),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_501),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_466),
.B1(n_450),
.B2(n_462),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_454),
.C(n_462),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_498),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_473),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_477),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_499),
.A2(n_474),
.B(n_448),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_457),
.C(n_451),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_500),
.B(n_472),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_453),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_468),
.Y(n_506)
);

INVx11_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_480),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_509),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_470),
.C(n_476),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_508),
.B(n_510),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_495),
.A2(n_484),
.B1(n_487),
.B2(n_488),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_479),
.C(n_475),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_518),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_484),
.B1(n_463),
.B2(n_460),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_512),
.A2(n_514),
.B1(n_504),
.B2(n_498),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_489),
.Y(n_522)
);

OAI21x1_ASAP7_75t_SL g515 ( 
.A1(n_503),
.A2(n_471),
.B(n_431),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_515),
.A2(n_517),
.B(n_501),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_490),
.B(n_460),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_460),
.C(n_333),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_519),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_524),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_523),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_508),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_497),
.C(n_500),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_499),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_509),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_527),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_529),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_528),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_519),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_534),
.A2(n_528),
.B(n_525),
.Y(n_538)
);

AOI21xp33_ASAP7_75t_L g541 ( 
.A1(n_536),
.A2(n_537),
.B(n_538),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_532),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_520),
.C(n_507),
.Y(n_539)
);

AO221x1_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_520),
.B1(n_535),
.B2(n_533),
.C(n_514),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_505),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_543),
.B(n_489),
.C(n_502),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_541),
.A2(n_492),
.B1(n_494),
.B2(n_491),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_333),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_290),
.Y(n_546)
);


endmodule