module fake_jpeg_30365_n_188 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_0),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_30),
.B1(n_17),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_68),
.B1(n_71),
.B2(n_1),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_55),
.B(n_60),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_17),
.C(n_29),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_20),
.C(n_19),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_17),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_16),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_26),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_25),
.B1(n_29),
.B2(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_25),
.B1(n_28),
.B2(n_15),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_16),
.B1(n_2),
.B2(n_4),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_72),
.B1(n_85),
.B2(n_80),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_76),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_26),
.B(n_18),
.C(n_20),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_28),
.B1(n_18),
.B2(n_16),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_63),
.B1(n_50),
.B2(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_92),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_16),
.B1(n_2),
.B2(n_4),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_97),
.B1(n_6),
.B2(n_7),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_67),
.C(n_61),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_58),
.B1(n_50),
.B2(n_48),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_118),
.B1(n_120),
.B2(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_58),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_64),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_59),
.C(n_7),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_93),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_125),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_89),
.B1(n_96),
.B2(n_94),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_130),
.B1(n_137),
.B2(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_74),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_120),
.B1(n_103),
.B2(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_124),
.B1(n_126),
.B2(n_130),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_137),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_124),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_113),
.B(n_116),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_147),
.B(n_150),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_103),
.B(n_110),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_101),
.B(n_109),
.C(n_115),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_131),
.B(n_138),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_108),
.B(n_74),
.C(n_59),
.D(n_91),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_124),
.B1(n_126),
.B2(n_129),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_155),
.B1(n_143),
.B2(n_147),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_146),
.B(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_139),
.C(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_108),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_162),
.B(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_168),
.B1(n_8),
.B2(n_9),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_165),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_8),
.B(n_9),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_150),
.B1(n_74),
.B2(n_10),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_161),
.B1(n_156),
.B2(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_168),
.B1(n_166),
.B2(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_157),
.C(n_160),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

NOR4xp25_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_164),
.C(n_12),
.D(n_10),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_R g183 ( 
.A(n_178),
.B(n_12),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_172),
.B1(n_171),
.B2(n_176),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_180),
.B(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_182),
.B(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_167),
.C(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_10),
.Y(n_188)
);


endmodule