module fake_ibex_441_n_1347 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1347);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1347;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_377;
wire n_647;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_339;
wire n_276;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_245;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1277;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_138),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_99),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_146),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_8),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_51),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_97),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_144),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_148),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_28),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_200),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_104),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_61),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_142),
.B(n_87),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_156),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_177),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_145),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_113),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_129),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_163),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_46),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_162),
.B(n_149),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_65),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_223),
.Y(n_283)
);

INVx4_ASAP7_75t_R g284 ( 
.A(n_128),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_160),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_36),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_132),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_20),
.B(n_158),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_77),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_126),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_174),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_94),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_75),
.Y(n_295)
);

BUFx2_ASAP7_75t_SL g296 ( 
.A(n_181),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_201),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_166),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_60),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_35),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_38),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_196),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_78),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_27),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_107),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_152),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_16),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_213),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_164),
.B(n_244),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_0),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_60),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_11),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_9),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_161),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_66),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_76),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_239),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_176),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_159),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_116),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_112),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_7),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_168),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_38),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_217),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_230),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_117),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_153),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_143),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_194),
.B(n_77),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_188),
.B(n_219),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_236),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_130),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_205),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_72),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_135),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_110),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_212),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_67),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_231),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_61),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_169),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_127),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_137),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_72),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_184),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_220),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_179),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_170),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_195),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_23),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_105),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_78),
.B(n_218),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_180),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_211),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_42),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_35),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_91),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_109),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_121),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_84),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_183),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_125),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_178),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_147),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_51),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_224),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_92),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_30),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_228),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_93),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_206),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_9),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_58),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_70),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_30),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_102),
.B(n_155),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_167),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_11),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_151),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_7),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_12),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_16),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_45),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_68),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_31),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_45),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_95),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_242),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_89),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_70),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_165),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_237),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_225),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_32),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_141),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_34),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_172),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_240),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_221),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_171),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_25),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_26),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_85),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_186),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_215),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_120),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_226),
.B(n_139),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_123),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_136),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_235),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_111),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_76),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_187),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_122),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_134),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_50),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_66),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_190),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_124),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_6),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_173),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_191),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_29),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_54),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_73),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_29),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_22),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_131),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_175),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_28),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_305),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_300),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_248),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_252),
.B(n_0),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_288),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_248),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_300),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_245),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_315),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_305),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_315),
.A2(n_88),
.B(n_86),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_399),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_330),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g450 ( 
.A1(n_330),
.A2(n_338),
.B(n_332),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_288),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_303),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_260),
.B(n_4),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_277),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_245),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_332),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_277),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_339),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_421),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_245),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_256),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_363),
.B(n_5),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_338),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_363),
.B(n_8),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_339),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_355),
.B(n_10),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_355),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_245),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_255),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_388),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_274),
.B(n_10),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_428),
.B(n_267),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_428),
.Y(n_482)
);

INVx6_ASAP7_75t_L g483 ( 
.A(n_255),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_362),
.B(n_13),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_264),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_246),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_247),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_249),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_283),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_253),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_431),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_255),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_251),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_327),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_255),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_434),
.B(n_14),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_254),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_325),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_327),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_418),
.B(n_90),
.Y(n_505)
);

NAND2x1_ASAP7_75t_L g506 ( 
.A(n_284),
.B(n_431),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_316),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_257),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_431),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_316),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_420),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_323),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_323),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_325),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_325),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_261),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_296),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_258),
.B(n_19),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_263),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_250),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_325),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_278),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_352),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_266),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_268),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_269),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_450),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_501),
.B(n_270),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_447),
.A2(n_276),
.B(n_272),
.Y(n_529)
);

INVxp33_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_505),
.B(n_381),
.Y(n_531)
);

INVxp33_ASAP7_75t_SL g532 ( 
.A(n_465),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_473),
.A2(n_487),
.B1(n_490),
.B2(n_489),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_446),
.B(n_436),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_446),
.A2(n_348),
.B1(n_353),
.B2(n_331),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_491),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_491),
.A2(n_348),
.B1(n_353),
.B2(n_331),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_450),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_489),
.B(n_281),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_460),
.B(n_273),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_490),
.B(n_496),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_456),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_456),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_460),
.B(n_398),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_512),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_460),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_485),
.Y(n_549)
);

NOR2x1p5_ASAP7_75t_L g550 ( 
.A(n_465),
.B(n_328),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_481),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_455),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_517),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_444),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_520),
.B(n_282),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_459),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_462),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_506),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_398),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_496),
.A2(n_280),
.B1(n_287),
.B2(n_285),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_462),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_507),
.A2(n_406),
.B1(n_345),
.B2(n_291),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_447),
.A2(n_294),
.B(n_286),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_481),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_511),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_469),
.Y(n_569)
);

AND3x2_ASAP7_75t_L g570 ( 
.A(n_480),
.B(n_289),
.C(n_290),
.Y(n_570)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_470),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_464),
.Y(n_572)
);

INVxp33_ASAP7_75t_L g573 ( 
.A(n_466),
.Y(n_573)
);

NOR2x1p5_ASAP7_75t_L g574 ( 
.A(n_511),
.B(n_295),
.Y(n_574)
);

INVxp33_ASAP7_75t_SL g575 ( 
.A(n_466),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_464),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_522),
.Y(n_577)
);

AND3x1_ASAP7_75t_L g578 ( 
.A(n_507),
.B(n_306),
.C(n_302),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_502),
.B(n_297),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_502),
.B(n_298),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_463),
.A2(n_517),
.B1(n_468),
.B2(n_439),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_464),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_438),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_438),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_476),
.Y(n_587)
);

INVx6_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_441),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_441),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_512),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_463),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_505),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_480),
.Y(n_595)
);

NOR2x1p5_ASAP7_75t_L g596 ( 
.A(n_513),
.B(n_479),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_484),
.B(n_326),
.C(n_312),
.Y(n_597)
);

NOR2x1p5_ASAP7_75t_L g598 ( 
.A(n_513),
.B(n_309),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_508),
.A2(n_358),
.B1(n_402),
.B2(n_374),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_510),
.B(n_313),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_508),
.B(n_299),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_519),
.A2(n_318),
.B1(n_319),
.B2(n_314),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_445),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_519),
.B(n_421),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_524),
.A2(n_343),
.B1(n_361),
.B2(n_349),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_478),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_451),
.B(n_301),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_479),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_505),
.B(n_352),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_449),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_524),
.B(n_525),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_458),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_518),
.B(n_358),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_448),
.A2(n_329),
.B1(n_402),
.B2(n_374),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_516),
.B(n_378),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_478),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_516),
.B(n_307),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

INVxp33_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_500),
.Y(n_622)
);

OAI22x1_ASAP7_75t_L g623 ( 
.A1(n_510),
.A2(n_412),
.B1(n_406),
.B2(n_345),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_500),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_453),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_467),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_437),
.B(n_317),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_471),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_471),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_454),
.A2(n_321),
.B(n_320),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_475),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_495),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_500),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_R g636 ( 
.A(n_437),
.B(n_329),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_499),
.B(n_322),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_486),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_515),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_443),
.B(n_324),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_443),
.B(n_380),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_488),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_504),
.B(n_352),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_497),
.A2(n_498),
.B1(n_472),
.B2(n_474),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_495),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_515),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_504),
.B(n_461),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_498),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_515),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_461),
.B(n_385),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_495),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_521),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_521),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_521),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_472),
.B(n_360),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_474),
.A2(n_336),
.B(n_333),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_521),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_537),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_567),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_621),
.B(n_477),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_534),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_531),
.A2(n_341),
.B(n_337),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_551),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_554),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_527),
.A2(n_346),
.B(n_344),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_575),
.A2(n_424),
.B1(n_365),
.B2(n_377),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_595),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_604),
.B(n_424),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_553),
.B(n_259),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_575),
.A2(n_386),
.B1(n_390),
.B2(n_389),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_551),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_548),
.B(n_482),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_593),
.B(n_482),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_588),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_536),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_262),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_559),
.B(n_271),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_569),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_621),
.B(n_275),
.Y(n_680)
);

BUFx8_ASAP7_75t_L g681 ( 
.A(n_549),
.Y(n_681)
);

AOI221xp5_ASAP7_75t_L g682 ( 
.A1(n_530),
.A2(n_492),
.B1(n_422),
.B2(n_425),
.C(n_429),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_546),
.B(n_304),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_599),
.B(n_430),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_569),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_571),
.B(n_435),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_636),
.A2(n_373),
.B1(n_383),
.B2(n_379),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_638),
.B(n_292),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_571),
.B(n_435),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_561),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_559),
.B(n_308),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_634),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_566),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_566),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_651),
.A2(n_334),
.B1(n_351),
.B2(n_347),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_533),
.B(n_359),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_578),
.A2(n_391),
.B1(n_395),
.B2(n_387),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_594),
.B(n_340),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_581),
.B(n_342),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_577),
.B(n_364),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_651),
.A2(n_367),
.B1(n_376),
.B2(n_375),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_582),
.B(n_382),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_L g703 ( 
.A(n_597),
.B(n_493),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_538),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_544),
.B(n_310),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_560),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_545),
.B(n_563),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_564),
.B(n_615),
.C(n_616),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_558),
.B(n_350),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_556),
.B(n_354),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_550),
.B(n_357),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_648),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_609),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_552),
.B(n_356),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_557),
.B(n_366),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_573),
.B(n_368),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_SL g718 ( 
.A(n_568),
.B(n_408),
.C(n_407),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_574),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_631),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_586),
.Y(n_722)
);

O2A1O1Ixp5_ASAP7_75t_L g723 ( 
.A1(n_528),
.A2(n_384),
.B(n_396),
.C(n_394),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_656),
.B(n_417),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_609),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_535),
.A2(n_409),
.B1(n_400),
.B2(n_405),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_627),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_617),
.B(n_289),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_584),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_588),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_585),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_543),
.B(n_410),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_543),
.B(n_411),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_564),
.B(n_625),
.C(n_592),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_596),
.B(n_265),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_589),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_535),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_600),
.A2(n_415),
.B1(n_423),
.B2(n_414),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_570),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_590),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_598),
.B(n_279),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_532),
.B(n_641),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_632),
.B(n_293),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_591),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_603),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_601),
.B(n_404),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_547),
.B(n_413),
.C(n_416),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_539),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_427),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_539),
.B(n_311),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_SL g751 ( 
.A(n_610),
.B(n_433),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_613),
.B(n_311),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_657),
.B(n_335),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_613),
.B(n_493),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_562),
.B(n_493),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_601),
.B(n_369),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_611),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_614),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_541),
.A2(n_494),
.B1(n_509),
.B2(n_483),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_607),
.B(n_369),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_607),
.B(n_369),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_540),
.B(n_495),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_626),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_630),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_623),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_633),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_541),
.B(n_503),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_579),
.A2(n_371),
.B1(n_372),
.B2(n_392),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_643),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_579),
.B(n_503),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_629),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_562),
.B(n_371),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_580),
.B(n_503),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_637),
.Y(n_775)
);

AND2x4_ASAP7_75t_SL g776 ( 
.A(n_600),
.B(n_392),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_600),
.A2(n_483),
.B1(n_457),
.B2(n_397),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_619),
.A2(n_397),
.B1(n_483),
.B2(n_457),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_619),
.B(n_503),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_649),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_602),
.A2(n_457),
.B1(n_397),
.B2(n_514),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_529),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_640),
.B(n_21),
.Y(n_783)
);

OAI221xp5_ASAP7_75t_L g784 ( 
.A1(n_602),
.A2(n_514),
.B1(n_523),
.B2(n_521),
.C(n_25),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_640),
.B(n_514),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_637),
.B(n_514),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_605),
.A2(n_514),
.B1(n_523),
.B2(n_24),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_529),
.B(n_523),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_565),
.B(n_523),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_652),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_645),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_652),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_646),
.B(n_27),
.Y(n_793)
);

AND2x6_ASAP7_75t_SL g794 ( 
.A(n_644),
.B(n_31),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_646),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_612),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_612),
.B(n_33),
.Y(n_797)
);

AND2x2_ASAP7_75t_SL g798 ( 
.A(n_583),
.B(n_33),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_555),
.B(n_34),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_583),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_583),
.B(n_98),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_555),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_659),
.B(n_662),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_737),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_708),
.A2(n_658),
.B(n_655),
.C(n_654),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_659),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_665),
.B(n_36),
.Y(n_807)
);

BUFx12f_ASAP7_75t_L g808 ( 
.A(n_681),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_742),
.B(n_37),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_686),
.A2(n_689),
.B(n_677),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_734),
.B(n_576),
.C(n_572),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_698),
.B(n_773),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_773),
.A2(n_622),
.B1(n_650),
.B2(n_647),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_663),
.A2(n_653),
.B(n_642),
.C(n_639),
.Y(n_814)
);

CKINVDCx6p67_ASAP7_75t_R g815 ( 
.A(n_665),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_737),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_698),
.B(n_668),
.Y(n_817)
);

XOR2x2_ASAP7_75t_L g818 ( 
.A(n_667),
.B(n_39),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_669),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_661),
.B(n_40),
.Y(n_820)
);

OA22x2_ASAP7_75t_L g821 ( 
.A1(n_684),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_737),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_661),
.B(n_41),
.Y(n_823)
);

NOR2x1_ASAP7_75t_L g824 ( 
.A(n_718),
.B(n_642),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_724),
.B(n_43),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_681),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_696),
.A2(n_620),
.B1(n_635),
.B2(n_628),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_675),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_728),
.B(n_43),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_721),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_707),
.B(n_48),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_666),
.A2(n_624),
.B(n_620),
.C(n_618),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_748),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_738),
.A2(n_618),
.B(n_606),
.C(n_50),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_719),
.B(n_48),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_695),
.B(n_49),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_776),
.B(n_735),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_684),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_692),
.B(n_587),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_746),
.B(n_683),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_684),
.B(n_49),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_716),
.B(n_52),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_696),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_739),
.B(n_53),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_692),
.B(n_56),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_777),
.B(n_56),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_715),
.B(n_710),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_748),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_676),
.B(n_57),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_671),
.B(n_57),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_666),
.A2(n_58),
.B(n_59),
.C(n_62),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_687),
.B(n_59),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_692),
.B(n_62),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_798),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_664),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_692),
.B(n_63),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_705),
.B(n_64),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_703),
.B(n_67),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_701),
.B(n_68),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_747),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_704),
.A2(n_697),
.B1(n_712),
.B2(n_673),
.Y(n_861)
);

O2A1O1Ixp5_ASAP7_75t_L g862 ( 
.A1(n_743),
.A2(n_699),
.B(n_751),
.C(n_723),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_680),
.B(n_74),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_726),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_80),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_783),
.A2(n_731),
.B(n_736),
.C(n_729),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_674),
.B(n_80),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_740),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_672),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_744),
.A2(n_758),
.B(n_759),
.C(n_745),
.Y(n_870)
);

AND2x2_ASAP7_75t_SL g871 ( 
.A(n_749),
.B(n_82),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_770),
.A2(n_84),
.B1(n_100),
.B2(n_101),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_755),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_722),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_697),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_730),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_693),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_792),
.Y(n_878)
);

CKINVDCx10_ASAP7_75t_R g879 ( 
.A(n_766),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_694),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_682),
.B(n_118),
.C(n_119),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_670),
.A2(n_691),
.B(n_678),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_764),
.A2(n_765),
.B1(n_780),
.B2(n_767),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_688),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_712),
.B(n_140),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_791),
.B(n_157),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_732),
.A2(n_733),
.B1(n_775),
.B2(n_711),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_794),
.Y(n_888)
);

BUFx5_ASAP7_75t_L g889 ( 
.A(n_714),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_777),
.B(n_185),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_741),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_891)
);

OA22x2_ASAP7_75t_L g892 ( 
.A1(n_741),
.A2(n_238),
.B1(n_199),
.B2(n_202),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_781),
.B(n_197),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_732),
.A2(n_733),
.B1(n_752),
.B2(n_700),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_743),
.A2(n_204),
.B1(n_207),
.B2(n_209),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_754),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_781),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_754),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_792),
.B(n_234),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_792),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_702),
.A2(n_787),
.B1(n_679),
.B2(n_685),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_757),
.A2(n_785),
.B(n_727),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_795),
.A2(n_768),
.B(n_771),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_750),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_660),
.B(n_709),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_720),
.B(n_725),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_774),
.A2(n_802),
.B(n_779),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_796),
.B(n_784),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_750),
.A2(n_793),
.B1(n_786),
.B2(n_762),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_799),
.A2(n_760),
.B(n_761),
.C(n_790),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_796),
.B(n_778),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_797),
.B(n_769),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_801),
.B(n_800),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_798),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_756),
.Y(n_915)
);

AO22x1_ASAP7_75t_L g916 ( 
.A1(n_681),
.A2(n_599),
.B1(n_536),
.B2(n_538),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_772),
.B(n_713),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_659),
.B(n_536),
.Y(n_918)
);

AOI221xp5_ASAP7_75t_L g919 ( 
.A1(n_708),
.A2(n_564),
.B1(n_530),
.B2(n_697),
.C(n_578),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_763),
.A2(n_531),
.B(n_690),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_713),
.A2(n_575),
.B1(n_773),
.B2(n_533),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_713),
.A2(n_575),
.B1(n_773),
.B2(n_533),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_706),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_659),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_659),
.B(n_530),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_662),
.B(n_530),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_763),
.A2(n_531),
.B(n_690),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_772),
.B(n_713),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_772),
.B(n_713),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_663),
.A2(n_666),
.B(n_772),
.C(n_690),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_772),
.B(n_713),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_763),
.A2(n_531),
.B(n_690),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_808),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_917),
.B(n_928),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_925),
.B(n_803),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_914),
.A2(n_922),
.B1(n_921),
.B2(n_929),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_918),
.B(n_810),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_915),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_861),
.B(n_926),
.Y(n_939)
);

OAI22xp33_ASAP7_75t_L g940 ( 
.A1(n_914),
.A2(n_919),
.B1(n_846),
.B2(n_826),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_815),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_804),
.Y(n_942)
);

CKINVDCx8_ASAP7_75t_R g943 ( 
.A(n_879),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_897),
.A2(n_846),
.B1(n_831),
.B2(n_829),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_832),
.A2(n_903),
.B(n_870),
.Y(n_945)
);

OAI22x1_ASAP7_75t_L g946 ( 
.A1(n_831),
.A2(n_841),
.B1(n_838),
.B2(n_916),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_SL g947 ( 
.A(n_817),
.B(n_878),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_804),
.Y(n_948)
);

NOR4xp25_ASAP7_75t_L g949 ( 
.A(n_843),
.B(n_851),
.C(n_866),
.D(n_834),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_816),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_850),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_SL g952 ( 
.A(n_893),
.B(n_871),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_887),
.A2(n_898),
.B(n_896),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_846),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_907),
.A2(n_908),
.B(n_862),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_884),
.B(n_809),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_893),
.A2(n_840),
.B1(n_886),
.B2(n_820),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_819),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_819),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_893),
.Y(n_960)
);

AO21x2_ASAP7_75t_L g961 ( 
.A1(n_902),
.A2(n_812),
.B(n_908),
.Y(n_961)
);

BUFx8_ASAP7_75t_L g962 ( 
.A(n_837),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_818),
.B(n_849),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_825),
.B(n_847),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_852),
.B(n_836),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_883),
.A2(n_823),
.B(n_901),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_828),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_878),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_855),
.B(n_869),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_813),
.A2(n_811),
.B(n_814),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_877),
.B(n_880),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_821),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_888),
.B(n_844),
.Y(n_973)
);

OAI22x1_ASAP7_75t_L g974 ( 
.A1(n_860),
.A2(n_858),
.B1(n_875),
.B2(n_857),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_858),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_807),
.B(n_885),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_912),
.A2(n_899),
.B(n_839),
.Y(n_977)
);

AO31x2_ASAP7_75t_L g978 ( 
.A1(n_910),
.A2(n_827),
.A3(n_872),
.B(n_913),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_835),
.B(n_904),
.Y(n_979)
);

CKINVDCx16_ASAP7_75t_R g980 ( 
.A(n_890),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_865),
.B(n_842),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_867),
.B(n_859),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_878),
.B(n_900),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_900),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_909),
.A2(n_881),
.B(n_882),
.Y(n_985)
);

CKINVDCx11_ASAP7_75t_R g986 ( 
.A(n_868),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_900),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_906),
.B(n_923),
.Y(n_988)
);

NAND3x1_ASAP7_75t_L g989 ( 
.A(n_891),
.B(n_824),
.C(n_895),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_845),
.A2(n_856),
.B(n_853),
.C(n_911),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_905),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_822),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_833),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_892),
.A2(n_830),
.B1(n_874),
.B2(n_876),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_848),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_889),
.B(n_917),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_L g997 ( 
.A1(n_812),
.A2(n_753),
.B(n_863),
.C(n_862),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_920),
.A2(n_531),
.B(n_927),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_917),
.B(n_928),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_917),
.B(n_928),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_917),
.B(n_928),
.Y(n_1001)
);

AO31x2_ASAP7_75t_L g1002 ( 
.A1(n_866),
.A2(n_782),
.A3(n_789),
.B(n_788),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_806),
.B(n_659),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_917),
.B(n_928),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_920),
.A2(n_531),
.B(n_927),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_925),
.B(n_659),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_804),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_914),
.A2(n_921),
.B1(n_922),
.B2(n_917),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_920),
.A2(n_932),
.B(n_927),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_808),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_806),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_808),
.Y(n_1012)
);

BUFx4f_ASAP7_75t_L g1013 ( 
.A(n_808),
.Y(n_1013)
);

CKINVDCx11_ASAP7_75t_R g1014 ( 
.A(n_808),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_808),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_918),
.B(n_659),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_806),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_808),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_804),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_924),
.B(n_917),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_917),
.B(n_928),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_920),
.A2(n_932),
.B(n_927),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_806),
.B(n_659),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_806),
.B(n_659),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_840),
.A2(n_929),
.B(n_928),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_924),
.B(n_917),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_930),
.A2(n_840),
.B(n_805),
.C(n_857),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_SL g1028 ( 
.A1(n_893),
.A2(n_846),
.B(n_930),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_917),
.B(n_928),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_920),
.A2(n_932),
.B(n_927),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_806),
.B(n_659),
.Y(n_1031)
);

AOI211x1_ASAP7_75t_L g1032 ( 
.A1(n_894),
.A2(n_921),
.B(n_922),
.C(n_927),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_866),
.A2(n_782),
.A3(n_789),
.B(n_788),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_806),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_925),
.B(n_659),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_917),
.B(n_928),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_920),
.A2(n_932),
.B(n_927),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_808),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_917),
.B(n_928),
.Y(n_1039)
);

INVx3_ASAP7_75t_SL g1040 ( 
.A(n_815),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_917),
.B(n_928),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_930),
.A2(n_840),
.B(n_805),
.C(n_857),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_914),
.A2(n_921),
.B1(n_922),
.B2(n_917),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_808),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_917),
.B(n_928),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_914),
.A2(n_708),
.B1(n_919),
.B2(n_886),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_920),
.A2(n_932),
.B(n_927),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_866),
.A2(n_782),
.A3(n_789),
.B(n_788),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_930),
.A2(n_928),
.B(n_931),
.C(n_929),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_918),
.B(n_659),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_918),
.B(n_659),
.Y(n_1051)
);

AO32x2_ASAP7_75t_L g1052 ( 
.A1(n_854),
.A2(n_864),
.A3(n_873),
.B1(n_922),
.B2(n_921),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_808),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_806),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_957),
.A2(n_944),
.B1(n_954),
.B2(n_960),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_984),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_954),
.A2(n_1046),
.B1(n_980),
.B2(n_1008),
.Y(n_1057)
);

OR3x4_ASAP7_75t_SL g1058 ( 
.A(n_943),
.B(n_1014),
.C(n_1013),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_955),
.A2(n_1022),
.B(n_1009),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_1053),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1040),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_974),
.A2(n_940),
.B(n_952),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_993),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_1054),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1054),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_952),
.B(n_994),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_1030),
.A2(n_1047),
.B(n_1037),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1006),
.B(n_1035),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_1011),
.Y(n_1069)
);

AOI21xp33_ASAP7_75t_SL g1070 ( 
.A1(n_941),
.A2(n_933),
.B(n_946),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1042),
.A2(n_1005),
.B(n_998),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_1017),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_935),
.B(n_934),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_1012),
.B(n_1015),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_993),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1020),
.B(n_1026),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_1013),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_999),
.B(n_1000),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1001),
.B(n_1004),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_1028),
.B(n_959),
.Y(n_1080)
);

CKINVDCx11_ASAP7_75t_R g1081 ( 
.A(n_1018),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_939),
.A2(n_1046),
.B1(n_937),
.B2(n_936),
.Y(n_1082)
);

OAI21xp33_ASAP7_75t_SL g1083 ( 
.A1(n_953),
.A2(n_966),
.B(n_996),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_SL g1084 ( 
.A1(n_1043),
.A2(n_972),
.B1(n_963),
.B2(n_1051),
.Y(n_1084)
);

AO21x2_ASAP7_75t_L g1085 ( 
.A1(n_945),
.A2(n_970),
.B(n_985),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_1012),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_938),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_1012),
.B(n_1015),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_965),
.A2(n_1016),
.B1(n_1050),
.B2(n_986),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_968),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_981),
.A2(n_964),
.B(n_990),
.C(n_997),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1029),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1036),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_1010),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1039),
.A2(n_1045),
.B(n_1041),
.C(n_956),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_951),
.B(n_1032),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_961),
.A2(n_949),
.B(n_977),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1024),
.B(n_1031),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_949),
.B(n_1034),
.C(n_1023),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1015),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_991),
.A2(n_976),
.B(n_969),
.C(n_971),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_983),
.A2(n_995),
.B(n_989),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_988),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_976),
.A2(n_992),
.B(n_950),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_973),
.B(n_975),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_987),
.A2(n_1048),
.B(n_1033),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_1002),
.A2(n_1048),
.B(n_1033),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1002),
.B(n_1048),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_1002),
.A2(n_1033),
.B(n_978),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_968),
.A2(n_1052),
.B(n_967),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_947),
.A2(n_978),
.B(n_1052),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_978),
.B(n_979),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_1010),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1052),
.A2(n_942),
.A3(n_948),
.B(n_1019),
.Y(n_1114)
);

BUFx8_ASAP7_75t_L g1115 ( 
.A(n_1038),
.Y(n_1115)
);

OA21x2_ASAP7_75t_L g1116 ( 
.A1(n_1007),
.A2(n_1019),
.B(n_958),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_962),
.B(n_1044),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1044),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_962),
.B(n_1046),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1027),
.A2(n_1042),
.B(n_927),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_1012),
.B(n_808),
.Y(n_1121)
);

NAND2x1p5_ASAP7_75t_L g1122 ( 
.A(n_954),
.B(n_914),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_960),
.B(n_808),
.Y(n_1123)
);

INVxp33_ASAP7_75t_L g1124 ( 
.A(n_1003),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_1027),
.B(n_1042),
.C(n_1032),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_952),
.B(n_994),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1040),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1049),
.A2(n_1025),
.B(n_982),
.C(n_1021),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_952),
.B(n_994),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1006),
.B(n_1035),
.Y(n_1130)
);

CKINVDCx8_ASAP7_75t_R g1131 ( 
.A(n_1012),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1027),
.B(n_1042),
.C(n_1032),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1076),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1116),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1103),
.B(n_1073),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1096),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1067),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1065),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1082),
.A2(n_1084),
.B1(n_1055),
.B2(n_1101),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1080),
.B(n_1104),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1065),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1084),
.A2(n_1057),
.B1(n_1082),
.B2(n_1062),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_SL g1143 ( 
.A(n_1131),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1116),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1078),
.B(n_1079),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1064),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1059),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1104),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1083),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_1071),
.A2(n_1110),
.B(n_1120),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1072),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1080),
.B(n_1102),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1114),
.Y(n_1153)
);

INVx4_ASAP7_75t_SL g1154 ( 
.A(n_1080),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_1081),
.Y(n_1155)
);

AO21x2_ASAP7_75t_L g1156 ( 
.A1(n_1071),
.A2(n_1120),
.B(n_1125),
.Y(n_1156)
);

AO21x2_ASAP7_75t_L g1157 ( 
.A1(n_1125),
.A2(n_1132),
.B(n_1111),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1087),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1106),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1119),
.B(n_1092),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_1090),
.Y(n_1161)
);

CKINVDCx14_ASAP7_75t_R g1162 ( 
.A(n_1061),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1068),
.B(n_1130),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1108),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1055),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1146),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1156),
.B(n_1107),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1152),
.B(n_1107),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1156),
.B(n_1109),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1156),
.B(n_1109),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1157),
.B(n_1149),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1161),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1138),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1160),
.B(n_1093),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1152),
.B(n_1097),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1152),
.B(n_1066),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1164),
.Y(n_1177)
);

AND2x2_ASAP7_75t_SL g1178 ( 
.A(n_1149),
.B(n_1112),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1164),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1138),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1159),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1154),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1139),
.A2(n_1057),
.B1(n_1062),
.B2(n_1119),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1147),
.B(n_1085),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1144),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1139),
.A2(n_1126),
.B1(n_1129),
.B2(n_1066),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1165),
.B(n_1099),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1136),
.B(n_1095),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1165),
.B(n_1136),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1152),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1161),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1191),
.B(n_1168),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1190),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1189),
.B(n_1148),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1172),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1167),
.B(n_1150),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1181),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1185),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1167),
.B(n_1150),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1188),
.B(n_1141),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1181),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1188),
.B(n_1141),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1173),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1167),
.B(n_1150),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1172),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1169),
.B(n_1153),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1183),
.A2(n_1142),
.B1(n_1126),
.B2(n_1129),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1172),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_1182),
.B(n_1134),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1192),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1189),
.B(n_1173),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1192),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_1180),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1192),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1170),
.B(n_1184),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1194),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1213),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1209),
.B(n_1210),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1199),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1198),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1218),
.B(n_1180),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1198),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_1199),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1218),
.B(n_1171),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1193),
.B(n_1175),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1212),
.B(n_1176),
.Y(n_1229)
);

NOR2x1_ASAP7_75t_L g1230 ( 
.A(n_1206),
.B(n_1121),
.Y(n_1230)
);

NAND2x1_ASAP7_75t_SL g1231 ( 
.A(n_1212),
.B(n_1182),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1218),
.B(n_1177),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1209),
.B(n_1171),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1202),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1210),
.B(n_1197),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1207),
.B(n_1177),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1214),
.B(n_1187),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1214),
.B(n_1187),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1207),
.B(n_1179),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1197),
.B(n_1171),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1197),
.B(n_1200),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1202),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1223),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1223),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1228),
.B(n_1196),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1225),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1219),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1225),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1230),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1221),
.B(n_1174),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1234),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1234),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1222),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1221),
.B(n_1195),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1226),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1224),
.A2(n_1183),
.B1(n_1174),
.B2(n_1208),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1219),
.Y(n_1257)
);

AOI21xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1229),
.A2(n_1088),
.B(n_1074),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1242),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1242),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1220),
.B(n_1201),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1254),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1243),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1249),
.A2(n_1229),
.B1(n_1211),
.B2(n_1196),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1261),
.B(n_1235),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1244),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1246),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1247),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1261),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1256),
.A2(n_1228),
.B1(n_1232),
.B2(n_1240),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1250),
.B(n_1241),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1248),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1250),
.A2(n_1163),
.B1(n_1135),
.B2(n_1145),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1251),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1255),
.B(n_1235),
.Y(n_1275)
);

AOI322xp5_ASAP7_75t_L g1276 ( 
.A1(n_1255),
.A2(n_1241),
.A3(n_1227),
.B1(n_1233),
.B2(n_1240),
.C1(n_1205),
.C2(n_1200),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1245),
.A2(n_1228),
.B1(n_1239),
.B2(n_1236),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1252),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1245),
.B(n_1233),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1253),
.B(n_1237),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1270),
.A2(n_1253),
.B1(n_1227),
.B2(n_1205),
.Y(n_1281)
);

AOI32xp33_ASAP7_75t_L g1282 ( 
.A1(n_1264),
.A2(n_1213),
.A3(n_1217),
.B1(n_1215),
.B2(n_1211),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1280),
.Y(n_1283)
);

OAI21xp33_ASAP7_75t_L g1284 ( 
.A1(n_1276),
.A2(n_1238),
.B(n_1237),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1263),
.B(n_1260),
.Y(n_1285)
);

AOI221xp5_ASAP7_75t_L g1286 ( 
.A1(n_1269),
.A2(n_1258),
.B1(n_1070),
.B2(n_1201),
.C(n_1203),
.Y(n_1286)
);

OAI321xp33_ASAP7_75t_L g1287 ( 
.A1(n_1269),
.A2(n_1229),
.A3(n_1238),
.B1(n_1088),
.B2(n_1074),
.C(n_1216),
.Y(n_1287)
);

AO22x1_ASAP7_75t_L g1288 ( 
.A1(n_1265),
.A2(n_1115),
.B1(n_1182),
.B2(n_1196),
.Y(n_1288)
);

OAI211xp5_ASAP7_75t_L g1289 ( 
.A1(n_1273),
.A2(n_1162),
.B(n_1089),
.C(n_1231),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1279),
.B(n_1229),
.Y(n_1290)
);

OAI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_1273),
.A2(n_1089),
.B1(n_1186),
.B2(n_1203),
.C(n_1216),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1287),
.A2(n_1277),
.B1(n_1275),
.B2(n_1271),
.Y(n_1292)
);

NOR3xp33_ASAP7_75t_L g1293 ( 
.A(n_1289),
.B(n_1117),
.C(n_1100),
.Y(n_1293)
);

OAI211xp5_ASAP7_75t_L g1294 ( 
.A1(n_1286),
.A2(n_1117),
.B(n_1127),
.C(n_1086),
.Y(n_1294)
);

AOI211xp5_ASAP7_75t_L g1295 ( 
.A1(n_1288),
.A2(n_1118),
.B(n_1058),
.C(n_1265),
.Y(n_1295)
);

AOI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1284),
.A2(n_1262),
.B1(n_1274),
.B2(n_1272),
.C(n_1278),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1283),
.A2(n_1143),
.B1(n_1267),
.B2(n_1266),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1281),
.A2(n_1211),
.B(n_1215),
.Y(n_1298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1299 ( 
.A1(n_1291),
.A2(n_1155),
.B(n_1204),
.C(n_1143),
.D(n_1158),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1282),
.B(n_1285),
.C(n_1115),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1285),
.B(n_1077),
.C(n_1099),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1290),
.B(n_1268),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1289),
.A2(n_1200),
.B1(n_1205),
.B2(n_1178),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1283),
.B(n_1268),
.Y(n_1304)
);

AOI211xp5_ASAP7_75t_L g1305 ( 
.A1(n_1292),
.A2(n_1118),
.B(n_1155),
.C(n_1105),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1300),
.A2(n_1095),
.B(n_1204),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1293),
.B(n_1118),
.Y(n_1307)
);

NAND4xp25_ASAP7_75t_L g1308 ( 
.A(n_1295),
.B(n_1186),
.C(n_1182),
.D(n_1128),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1296),
.B(n_1259),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1304),
.Y(n_1310)
);

NAND4xp25_ASAP7_75t_SL g1311 ( 
.A(n_1294),
.B(n_1155),
.C(n_1217),
.D(n_1187),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1301),
.B(n_1257),
.Y(n_1312)
);

AOI221xp5_ASAP7_75t_L g1313 ( 
.A1(n_1297),
.A2(n_1298),
.B1(n_1303),
.B2(n_1302),
.C(n_1299),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1296),
.B(n_1257),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1305),
.B(n_1069),
.C(n_1056),
.Y(n_1315)
);

NOR2x1_ASAP7_75t_L g1316 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1316)
);

NOR3xp33_ASAP7_75t_L g1317 ( 
.A(n_1313),
.B(n_1075),
.C(n_1063),
.Y(n_1317)
);

NAND4xp75_ASAP7_75t_L g1318 ( 
.A(n_1306),
.B(n_1094),
.C(n_1113),
.D(n_1163),
.Y(n_1318)
);

NOR3xp33_ASAP7_75t_L g1319 ( 
.A(n_1308),
.B(n_1075),
.C(n_1063),
.Y(n_1319)
);

NOR3xp33_ASAP7_75t_L g1320 ( 
.A(n_1314),
.B(n_1309),
.C(n_1310),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1312),
.B(n_1247),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1307),
.B(n_1123),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1310),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1320),
.B(n_1151),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1318),
.B(n_1060),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1323),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1321),
.B(n_1166),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_L g1328 ( 
.A(n_1317),
.B(n_1315),
.C(n_1316),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1319),
.Y(n_1329)
);

NOR2x1p5_ASAP7_75t_L g1330 ( 
.A(n_1322),
.B(n_1056),
.Y(n_1330)
);

NOR3xp33_ASAP7_75t_SL g1331 ( 
.A(n_1322),
.B(n_1091),
.C(n_1098),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1320),
.B(n_1151),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1327),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1329),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1325),
.B(n_1123),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1328),
.A2(n_1123),
.B(n_1122),
.Y(n_1336)
);

AND3x4_ASAP7_75t_L g1337 ( 
.A(n_1331),
.B(n_1140),
.C(n_1133),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1335),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1334),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1333),
.B(n_1326),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1339),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1341),
.A2(n_1338),
.B1(n_1340),
.B2(n_1337),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1341),
.Y(n_1343)
);

NOR2x1_ASAP7_75t_L g1344 ( 
.A(n_1343),
.B(n_1336),
.Y(n_1344)
);

AOI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1344),
.A2(n_1342),
.B1(n_1330),
.B2(n_1056),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1345),
.A2(n_1332),
.B(n_1324),
.Y(n_1346)
);

AOI21xp33_ASAP7_75t_L g1347 ( 
.A1(n_1346),
.A2(n_1124),
.B(n_1098),
.Y(n_1347)
);


endmodule