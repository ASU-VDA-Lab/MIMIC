module fake_jpeg_31439_n_167 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_44),
.Y(n_47)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_10),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_23),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_84),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_32),
.B(n_39),
.C(n_15),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_87),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_34),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_72),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_45),
.B1(n_22),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_19),
.B1(n_16),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_16),
.B1(n_29),
.B2(n_30),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_28),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_25),
.B1(n_17),
.B2(n_28),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_25),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_17),
.B1(n_63),
.B2(n_53),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_30),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_72),
.B1(n_84),
.B2(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_76),
.B1(n_87),
.B2(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_105),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_77),
.B1(n_73),
.B2(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_49),
.C(n_82),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_106),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_101),
.A3(n_91),
.B1(n_10),
.B2(n_9),
.C1(n_108),
.C2(n_103),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_9),
.C(n_2),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_70),
.B1(n_67),
.B2(n_64),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_108),
.B1(n_92),
.B2(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_82),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_29),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_131),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_109),
.B(n_95),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_110),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_105),
.B(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_133),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_116),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_113),
.B1(n_121),
.B2(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_134),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_112),
.B1(n_114),
.B2(n_121),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_113),
.B1(n_109),
.B2(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_142),
.A2(n_144),
.B1(n_124),
.B2(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_150),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_125),
.B(n_129),
.C(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_96),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_107),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_138),
.B(n_143),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_149),
.Y(n_157)
);

OAI221xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_154),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_56),
.B1(n_16),
.B2(n_3),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_1),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_1),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_159),
.C(n_64),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_4),
.B1(n_7),
.B2(n_161),
.C(n_153),
.Y(n_167)
);


endmodule