module fake_jpeg_16388_n_265 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_28),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_23),
.B1(n_25),
.B2(n_22),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_35),
.B1(n_50),
.B2(n_55),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_42),
.B(n_27),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_37),
.B1(n_23),
.B2(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_46),
.B1(n_51),
.B2(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_23),
.B1(n_25),
.B2(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_22),
.B2(n_14),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_24),
.C(n_28),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_31),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_18),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_30),
.A2(n_19),
.B1(n_22),
.B2(n_14),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_66),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_67),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_71),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_32),
.B(n_39),
.C(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_19),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_30),
.B1(n_34),
.B2(n_15),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_58),
.B1(n_51),
.B2(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_40),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_41),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_88),
.B1(n_63),
.B2(n_16),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_56),
.B1(n_54),
.B2(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_47),
.B1(n_40),
.B2(n_34),
.Y(n_88)
);

AO21x2_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_40),
.B(n_46),
.Y(n_90)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_59),
.B1(n_68),
.B2(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_71),
.B1(n_78),
.B2(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_40),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_104),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_33),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_67),
.B(n_73),
.C(n_65),
.D(n_46),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_75),
.C(n_64),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_122),
.C(n_89),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_65),
.B(n_41),
.C(n_66),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_70),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_64),
.A3(n_68),
.B1(n_17),
.B2(n_20),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_85),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_105),
.B1(n_82),
.B2(n_91),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_111),
.B(n_118),
.C(n_113),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_124),
.B1(n_96),
.B2(n_101),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_125),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_29),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_63),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_28),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_90),
.B1(n_103),
.B2(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_138),
.B1(n_145),
.B2(n_146),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_89),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_142),
.C(n_150),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_90),
.B(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_148),
.B(n_43),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_85),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_60),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_106),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_99),
.B1(n_83),
.B2(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_83),
.B(n_28),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_26),
.B(n_16),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_121),
.C(n_124),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_119),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_48),
.C(n_43),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_76),
.C(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_24),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_162),
.C(n_164),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_159),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_149),
.B1(n_114),
.B2(n_145),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_170),
.B1(n_173),
.B2(n_26),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_117),
.C(n_128),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_117),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_172),
.C(n_27),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_140),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_118),
.B1(n_115),
.B2(n_15),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_153),
.B1(n_146),
.B2(n_138),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_27),
.B(n_29),
.C(n_24),
.D(n_28),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_169),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_17),
.B1(n_20),
.B2(n_2),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_48),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_161),
.B(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_152),
.B1(n_148),
.B2(n_132),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_188),
.B1(n_194),
.B2(n_18),
.Y(n_210)
);

OAI321xp33_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_132),
.A3(n_26),
.B1(n_16),
.B2(n_18),
.C(n_10),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_193),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_162),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_29),
.B1(n_26),
.B2(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_12),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_176),
.B1(n_169),
.B2(n_157),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_209),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_208),
.B1(n_187),
.B2(n_183),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_168),
.C(n_176),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_212),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_186),
.B(n_178),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_172),
.C(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_197),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_154),
.C(n_24),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_211),
.C(n_184),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_13),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_0),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_18),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_210),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_27),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_179),
.B1(n_181),
.B2(n_178),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_211),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_224),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.C(n_220),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_192),
.C(n_24),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_192),
.Y(n_220)
);

XOR2x1_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_12),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_205),
.C(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_0),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_11),
.C(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_234),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_11),
.C(n_9),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_27),
.C(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.C(n_246),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_221),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_216),
.B(n_222),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_232),
.B(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_218),
.C(n_219),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_232),
.C(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_248),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_251),
.B1(n_8),
.B2(n_6),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_3),
.B(n_4),
.Y(n_250)
);

NOR3xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_253),
.C(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_242),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_4),
.C(n_5),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_238),
.C(n_244),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_254),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_255),
.A2(n_6),
.B(n_7),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_7),
.B(n_8),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_8),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_261),
.B(n_256),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_7),
.B(n_262),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);


endmodule