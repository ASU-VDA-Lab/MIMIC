module fake_jpeg_2121_n_194 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_71),
.Y(n_77)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_0),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_61),
.B1(n_43),
.B2(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_75),
.B1(n_67),
.B2(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_43),
.B1(n_60),
.B2(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_44),
.B1(n_62),
.B2(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_1),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_64),
.B1(n_44),
.B2(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_76),
.B1(n_83),
.B2(n_80),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_90),
.B1(n_92),
.B2(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_54),
.B1(n_58),
.B2(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_56),
.B1(n_48),
.B2(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_93),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_58),
.B1(n_70),
.B2(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_72),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_48),
.B(n_57),
.C(n_52),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_80),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_77),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_7),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_2),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_R g115 ( 
.A(n_85),
.B(n_57),
.Y(n_115)
);

XNOR2x2_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_35),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_87),
.B1(n_96),
.B2(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_3),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_137),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_52),
.B(n_4),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_131),
.B(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_52),
.B(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_134),
.B1(n_13),
.B2(n_14),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_7),
.B(n_9),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_106),
.C(n_110),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_151),
.C(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_10),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_11),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_153),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_102),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_114),
.C(n_20),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_12),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_156),
.B1(n_134),
.B2(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_16),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_122),
.B1(n_156),
.B2(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_165),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_126),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_142),
.C(n_149),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_170),
.B(n_171),
.Y(n_178)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_176),
.C(n_161),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_149),
.B(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_131),
.C(n_114),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_183),
.Y(n_184)
);

OAI322xp33_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_161),
.A3(n_159),
.B1(n_163),
.B2(n_166),
.C1(n_170),
.C2(n_28),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_166),
.B1(n_174),
.B2(n_178),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_179),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_179),
.A3(n_176),
.B1(n_175),
.B2(n_18),
.C(n_19),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_18),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_187),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_22),
.C(n_23),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_26),
.Y(n_194)
);


endmodule