module fake_jpeg_2529_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_48),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_19),
.B(n_15),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_55),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_53),
.B(n_59),
.Y(n_126)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_10),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_10),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_63),
.B(n_66),
.Y(n_127)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_7),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_32),
.B(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_40),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_20),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_40),
.B1(n_29),
.B2(n_35),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_89),
.A2(n_97),
.B1(n_101),
.B2(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_95),
.B(n_103),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_0),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_40),
.B1(n_29),
.B2(n_45),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_29),
.B1(n_41),
.B2(n_44),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_41),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_44),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_105),
.B(n_123),
.Y(n_179)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_108),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_13),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_31),
.C(n_39),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_108),
.C(n_114),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_35),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_76),
.A2(n_28),
.B1(n_39),
.B2(n_27),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_31),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_121),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_28),
.B1(n_20),
.B2(n_43),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_43),
.B1(n_21),
.B2(n_33),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_43),
.B1(n_21),
.B2(n_33),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_47),
.A2(n_43),
.B1(n_21),
.B2(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_61),
.A2(n_43),
.B1(n_21),
.B2(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_50),
.A2(n_87),
.B1(n_86),
.B2(n_85),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_104),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_69),
.A2(n_43),
.B1(n_21),
.B2(n_3),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_79),
.A2(n_21),
.B1(n_2),
.B2(n_4),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_162),
.Y(n_195)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_145),
.B(n_154),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_67),
.B1(n_54),
.B2(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_146),
.A2(n_152),
.B1(n_120),
.B2(n_111),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_12),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_91),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_11),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_158),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_13),
.B1(n_14),
.B2(n_0),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_175),
.B1(n_178),
.B2(n_137),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_90),
.A2(n_13),
.B(n_14),
.C(n_5),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_164),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_186),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_88),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_167),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_116),
.B(n_98),
.CI(n_139),
.CON(n_168),
.SN(n_168)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_92),
.B(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_134),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_92),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_187),
.Y(n_191)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_113),
.B(n_133),
.C(n_111),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_134),
.B1(n_111),
.B2(n_119),
.Y(n_207)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_93),
.B(n_113),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_183),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_122),
.B1(n_115),
.B2(n_128),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_107),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_185),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_115),
.C(n_137),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_208),
.B1(n_209),
.B2(n_214),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_204),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_117),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_100),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_221),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_174),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_146),
.A2(n_100),
.B1(n_119),
.B2(n_120),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_163),
.A2(n_111),
.B1(n_171),
.B2(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_151),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_182),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_147),
.A2(n_165),
.B1(n_156),
.B2(n_171),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_179),
.B1(n_167),
.B2(n_157),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_172),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_232),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_168),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_227),
.C(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_163),
.B(n_158),
.C(n_174),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g269 ( 
.A1(n_226),
.A2(n_215),
.B(n_188),
.C(n_211),
.D(n_193),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_170),
.C(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_230),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_149),
.B1(n_181),
.B2(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_236),
.B1(n_237),
.B2(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_197),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_161),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_239),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_183),
.B1(n_173),
.B2(n_180),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_178),
.B1(n_160),
.B2(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_153),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_144),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_245),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_196),
.A2(n_144),
.B1(n_143),
.B2(n_176),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_195),
.B(n_202),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_203),
.B(n_220),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_207),
.B(n_196),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_207),
.B(n_197),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_247),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_202),
.A3(n_195),
.B1(n_190),
.B2(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_190),
.B1(n_189),
.B2(n_209),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_234),
.B1(n_223),
.B2(n_246),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_269),
.B(n_256),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_192),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_263),
.C(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_239),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_268),
.B(n_226),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_208),
.B1(n_220),
.B2(n_218),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_266),
.B1(n_238),
.B2(n_225),
.Y(n_274)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_218),
.B1(n_210),
.B2(n_211),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_215),
.B(n_188),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_230),
.B1(n_234),
.B2(n_232),
.C(n_245),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_249),
.B1(n_262),
.B2(n_257),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_278),
.B1(n_285),
.B2(n_261),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_274),
.A2(n_267),
.B1(n_265),
.B2(n_264),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_282),
.C(n_284),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_243),
.A3(n_223),
.B1(n_247),
.B2(n_235),
.C1(n_228),
.C2(n_241),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_280),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_281),
.C(n_255),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_226),
.B1(n_236),
.B2(n_233),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_222),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_222),
.B(n_237),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_252),
.B(n_253),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_257),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_193),
.B1(n_213),
.B2(n_259),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_295),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_259),
.B1(n_269),
.B2(n_266),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_291),
.B(n_213),
.C(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.C(n_296),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_252),
.C(n_253),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_261),
.C(n_267),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_272),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_274),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_283),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_284),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_287),
.C(n_290),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_304),
.Y(n_313)
);

AOI321xp33_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_275),
.A3(n_280),
.B1(n_270),
.B2(n_291),
.C(n_279),
.Y(n_304)
);

AOI321xp33_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_279),
.A3(n_282),
.B1(n_272),
.B2(n_283),
.C(n_285),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_308),
.B1(n_288),
.B2(n_287),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_315),
.B1(n_308),
.B2(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_301),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_302),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_290),
.B1(n_297),
.B2(n_300),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_313),
.B1(n_310),
.B2(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_305),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_311),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_312),
.C(n_315),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_324),
.B1(n_318),
.B2(n_325),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_327),
.Y(n_328)
);


endmodule