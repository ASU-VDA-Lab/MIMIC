module fake_jpeg_9878_n_248 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_18),
.B1(n_14),
.B2(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_48),
.B1(n_33),
.B2(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_18),
.B1(n_26),
.B2(n_17),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_56),
.B1(n_33),
.B2(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_23),
.B1(n_17),
.B2(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_23),
.B1(n_28),
.B2(n_19),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_34),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_37),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_67),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_32),
.C(n_36),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_51),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_55),
.B1(n_50),
.B2(n_49),
.Y(n_88)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_66),
.B1(n_75),
.B2(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_59),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_57),
.B1(n_64),
.B2(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_100),
.B1(n_102),
.B2(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_64),
.C(n_67),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_104),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_65),
.B1(n_45),
.B2(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_107),
.B1(n_95),
.B2(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_47),
.B1(n_74),
.B2(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_110),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_63),
.B1(n_74),
.B2(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_60),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_67),
.B(n_36),
.Y(n_132)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_60),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_77),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_114),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_68),
.B1(n_44),
.B2(n_67),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_124),
.C(n_125),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_133),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_123),
.B(n_132),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_77),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_88),
.B1(n_92),
.B2(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_130),
.B1(n_44),
.B2(n_37),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_106),
.B1(n_115),
.B2(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_94),
.B1(n_91),
.B2(n_84),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_95),
.B1(n_81),
.B2(n_53),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_67),
.B(n_38),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_37),
.B(n_1),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_109),
.B(n_103),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_103),
.C(n_98),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_146),
.C(n_153),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_80),
.C(n_30),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_80),
.B1(n_95),
.B2(n_68),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_150),
.B1(n_155),
.B2(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_136),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_68),
.B(n_25),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_128),
.B1(n_120),
.B2(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_120),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_162),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_165),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_166),
.C(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_147),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_132),
.C(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_37),
.B1(n_52),
.B2(n_30),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_171),
.B1(n_52),
.B2(n_37),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_170),
.B(n_172),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_37),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_145),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_183),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_143),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_24),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_155),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_143),
.B(n_138),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_189),
.B(n_8),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_149),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_188),
.C(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_165),
.B1(n_157),
.B2(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_30),
.C(n_24),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_11),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_163),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_160),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_194),
.A2(n_205),
.B(n_5),
.C(n_8),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_25),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_177),
.B1(n_176),
.B2(n_189),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_172),
.C(n_30),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_19),
.C(n_2),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_9),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_11),
.B(n_13),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_11),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_176),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_24),
.CI(n_21),
.CON(n_204),
.SN(n_204)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_178),
.B1(n_24),
.B2(n_27),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_205),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_211),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_214),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_217),
.C(n_195),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_215),
.A2(n_6),
.B1(n_7),
.B2(n_5),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_198),
.C(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_221),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_206),
.Y(n_221)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_203),
.B(n_209),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_212),
.B(n_5),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_204),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_227),
.A2(n_212),
.B(n_217),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_234),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_232),
.B(n_25),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_6),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_7),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_228),
.B(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_0),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_232),
.C(n_231),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_0),
.C(n_2),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_2),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_3),
.B(n_4),
.C(n_199),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_246),
.B(n_3),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_4),
.Y(n_248)
);


endmodule