module real_aes_16962_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1146 ( .A1(n_0), .A2(n_196), .B1(n_1123), .B2(n_1134), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_1), .A2(n_6), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_1), .A2(n_227), .B1(n_522), .B2(n_523), .Y(n_521) );
OAI22xp33_ASAP7_75t_SL g730 ( .A1(n_2), .A2(n_124), .B1(n_562), .B2(n_576), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g741 ( .A1(n_2), .A2(n_26), .B1(n_301), .B2(n_742), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_3), .A2(n_27), .B1(n_354), .B2(n_634), .Y(n_775) );
OAI22xp5_ASAP7_75t_SL g783 ( .A1(n_3), .A2(n_127), .B1(n_301), .B2(n_339), .Y(n_783) );
INVx1_ASAP7_75t_L g1350 ( .A(n_4), .Y(n_1350) );
INVx1_ASAP7_75t_L g875 ( .A(n_5), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_6), .A2(n_231), .B1(n_432), .B2(n_522), .Y(n_533) );
INVx1_ASAP7_75t_L g1093 ( .A(n_7), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_8), .A2(n_248), .B1(n_523), .B2(n_548), .Y(n_547) );
INVxp33_ASAP7_75t_SL g600 ( .A(n_8), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_9), .A2(n_59), .B1(n_1123), .B2(n_1134), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_10), .Y(n_778) );
INVx1_ASAP7_75t_L g672 ( .A(n_11), .Y(n_672) );
INVx1_ASAP7_75t_L g859 ( .A(n_12), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_13), .Y(n_749) );
INVx1_ASAP7_75t_L g280 ( .A(n_14), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_14), .B(n_290), .Y(n_413) );
INVx1_ASAP7_75t_L g489 ( .A(n_15), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_15), .A2(n_39), .B1(n_322), .B2(n_507), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_16), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g704 ( .A(n_17), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_18), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_19), .A2(n_222), .B1(n_405), .B2(n_819), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_19), .A2(n_65), .B1(n_836), .B2(n_837), .Y(n_835) );
OAI222xp33_ASAP7_75t_L g796 ( .A1(n_20), .A2(n_202), .B1(n_355), .B2(n_493), .C1(n_797), .C2(n_798), .Y(n_796) );
OAI222xp33_ASAP7_75t_L g825 ( .A1(n_20), .A2(n_145), .B1(n_202), .B2(n_322), .C1(n_826), .C2(n_827), .Y(n_825) );
INVx1_ASAP7_75t_L g499 ( .A(n_21), .Y(n_499) );
INVx2_ASAP7_75t_L g1115 ( .A(n_22), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_22), .B(n_110), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_22), .B(n_1116), .Y(n_1130) );
OAI22xp33_ASAP7_75t_L g1332 ( .A1(n_23), .A2(n_180), .B1(n_282), .B2(n_562), .Y(n_1332) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_23), .A2(n_180), .B1(n_582), .B2(n_1057), .Y(n_1379) );
OAI22xp33_ASAP7_75t_SL g1340 ( .A1(n_24), .A2(n_25), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
OAI22xp33_ASAP7_75t_L g1383 ( .A1(n_24), .A2(n_25), .B1(n_597), .B2(n_1066), .Y(n_1383) );
OAI22xp33_ASAP7_75t_SL g727 ( .A1(n_26), .A2(n_235), .B1(n_354), .B2(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_27), .B(n_336), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_28), .A2(n_43), .B1(n_1128), .B2(n_1129), .Y(n_1159) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_29), .A2(n_207), .B1(n_301), .B2(n_877), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_29), .A2(n_260), .B1(n_354), .B2(n_636), .Y(n_886) );
INVx1_ASAP7_75t_L g1362 ( .A(n_30), .Y(n_1362) );
INVx1_ASAP7_75t_L g668 ( .A(n_31), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_32), .A2(n_200), .B1(n_916), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_32), .A2(n_225), .B1(n_433), .B2(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g810 ( .A(n_33), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_33), .A2(n_222), .B1(n_837), .B2(n_845), .Y(n_844) );
XOR2xp5_ASAP7_75t_L g699 ( .A(n_34), .B(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_34), .A2(n_123), .B1(n_1128), .B2(n_1129), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_35), .A2(n_163), .B1(n_562), .B2(n_633), .Y(n_1044) );
OAI22xp33_ASAP7_75t_L g1046 ( .A1(n_35), .A2(n_257), .B1(n_301), .B2(n_742), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_36), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_37), .A2(n_141), .B1(n_354), .B2(n_636), .Y(n_635) );
OAI22xp33_ASAP7_75t_SL g638 ( .A1(n_37), .A2(n_141), .B1(n_301), .B2(n_639), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_38), .Y(n_762) );
INVx1_ASAP7_75t_L g495 ( .A(n_39), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_40), .A2(n_195), .B1(n_354), .B2(n_485), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_40), .A2(n_105), .B1(n_301), .B2(n_742), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_41), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_42), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_44), .A2(n_115), .B1(n_556), .B2(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g614 ( .A(n_44), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_45), .A2(n_107), .B1(n_1123), .B2(n_1125), .Y(n_1122) );
INVx1_ASAP7_75t_L g299 ( .A(n_46), .Y(n_299) );
INVx1_ASAP7_75t_L g1004 ( .A(n_47), .Y(n_1004) );
OAI211xp5_ASAP7_75t_L g1009 ( .A1(n_47), .A2(n_641), .B(n_1010), .C(n_1013), .Y(n_1009) );
INVx1_ASAP7_75t_L g1083 ( .A(n_48), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_49), .A2(n_101), .B1(n_1123), .B2(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g500 ( .A(n_50), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_51), .Y(n_1031) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_52), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_53), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_54), .A2(n_148), .B1(n_322), .B2(n_328), .Y(n_321) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_54), .Y(n_366) );
INVx1_ASAP7_75t_L g630 ( .A(n_55), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_56), .A2(n_84), .B1(n_916), .B2(n_918), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g930 ( .A1(n_56), .A2(n_96), .B1(n_426), .B2(n_543), .Y(n_930) );
INVx1_ASAP7_75t_L g305 ( .A(n_57), .Y(n_305) );
INVx1_ASAP7_75t_L g320 ( .A(n_57), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_58), .A2(n_136), .B1(n_582), .B2(n_1057), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_58), .A2(n_136), .B1(n_282), .B2(n_562), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_60), .A2(n_130), .B1(n_1123), .B2(n_1155), .Y(n_1168) );
INVx1_ASAP7_75t_L g900 ( .A(n_61), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_61), .A2(n_109), .B1(n_328), .B2(n_671), .C(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_62), .A2(n_80), .B1(n_464), .B2(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g520 ( .A(n_62), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_63), .Y(n_752) );
XOR2x2_ASAP7_75t_L g295 ( .A(n_64), .B(n_296), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_64), .A2(n_218), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
INVx1_ASAP7_75t_L g811 ( .A(n_65), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_66), .A2(n_81), .B1(n_403), .B2(n_405), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_66), .A2(n_236), .B1(n_432), .B2(n_446), .Y(n_445) );
XOR2xp5_ASAP7_75t_L g846 ( .A(n_67), .B(n_847), .Y(n_846) );
OAI211xp5_ASAP7_75t_L g1000 ( .A1(n_68), .A2(n_627), .B(n_1001), .C(n_1002), .Y(n_1000) );
INVx1_ASAP7_75t_L g1014 ( .A(n_68), .Y(n_1014) );
INVx1_ASAP7_75t_L g273 ( .A(n_69), .Y(n_273) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_70), .A2(n_212), .B1(n_575), .B2(n_577), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_70), .A2(n_212), .B1(n_596), .B2(n_597), .Y(n_595) );
INVx2_ASAP7_75t_L g307 ( .A(n_71), .Y(n_307) );
INVx1_ASAP7_75t_L g852 ( .A(n_72), .Y(n_852) );
INVx1_ASAP7_75t_L g1363 ( .A(n_73), .Y(n_1363) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_74), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g367 ( .A1(n_74), .A2(n_148), .B1(n_368), .B2(n_372), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g963 ( .A1(n_75), .A2(n_253), .B1(n_336), .B2(n_339), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_75), .A2(n_253), .B1(n_633), .B2(n_634), .Y(n_969) );
INVx1_ASAP7_75t_L g553 ( .A(n_76), .Y(n_553) );
OAI22xp33_ASAP7_75t_SL g957 ( .A1(n_77), .A2(n_263), .B1(n_301), .B2(n_742), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_77), .A2(n_263), .B1(n_354), .B2(n_636), .Y(n_965) );
INVx1_ASAP7_75t_L g483 ( .A(n_78), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_79), .A2(n_105), .B1(n_562), .B2(n_576), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1015 ( .A1(n_79), .A2(n_195), .B1(n_336), .B2(n_339), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_80), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_81), .A2(n_91), .B1(n_432), .B2(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g657 ( .A(n_82), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_83), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_84), .A2(n_185), .B1(n_426), .B2(n_925), .Y(n_924) );
XOR2xp5_ASAP7_75t_L g788 ( .A(n_85), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g941 ( .A(n_86), .Y(n_941) );
INVx1_ASAP7_75t_L g571 ( .A(n_87), .Y(n_571) );
INVx1_ASAP7_75t_L g629 ( .A(n_88), .Y(n_629) );
INVx1_ASAP7_75t_L g725 ( .A(n_89), .Y(n_725) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_89), .A2(n_588), .B(n_734), .C(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g938 ( .A(n_90), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_91), .A2(n_236), .B1(n_400), .B2(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g491 ( .A(n_92), .Y(n_491) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_93), .B(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g1135 ( .A1(n_94), .A2(n_126), .B1(n_1128), .B2(n_1129), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_95), .A2(n_112), .B1(n_1123), .B2(n_1134), .Y(n_1151) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_96), .A2(n_185), .B1(n_479), .B2(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g973 ( .A(n_97), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_98), .A2(n_175), .B1(n_633), .B2(n_634), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_98), .A2(n_175), .B1(n_336), .B2(n_339), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g871 ( .A1(n_99), .A2(n_260), .B1(n_336), .B2(n_742), .C(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g884 ( .A(n_99), .Y(n_884) );
INVx1_ASAP7_75t_L g1089 ( .A(n_100), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_102), .A2(n_203), .B1(n_633), .B2(n_634), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_102), .A2(n_203), .B1(n_336), .B2(n_339), .Y(n_909) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_103), .Y(n_275) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_103), .B(n_273), .Y(n_1113) );
OAI211xp5_ASAP7_75t_L g791 ( .A1(n_104), .A2(n_792), .B(n_793), .C(n_802), .Y(n_791) );
INVx1_ASAP7_75t_L g831 ( .A(n_104), .Y(n_831) );
INVx1_ASAP7_75t_L g854 ( .A(n_106), .Y(n_854) );
INVx1_ASAP7_75t_L g1338 ( .A(n_108), .Y(n_1338) );
INVx1_ASAP7_75t_L g902 ( .A(n_109), .Y(n_902) );
INVx1_ASAP7_75t_L g1116 ( .A(n_110), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_110), .B(n_1115), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_111), .A2(n_171), .B1(n_1128), .B2(n_1129), .Y(n_1167) );
INVx1_ASAP7_75t_L g855 ( .A(n_113), .Y(n_855) );
INVx1_ASAP7_75t_L g334 ( .A(n_114), .Y(n_334) );
INVx1_ASAP7_75t_L g602 ( .A(n_115), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_116), .Y(n_1028) );
INVx2_ASAP7_75t_L g345 ( .A(n_117), .Y(n_345) );
INVx1_ASAP7_75t_L g444 ( .A(n_117), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_118), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_119), .A2(n_247), .B1(n_403), .B2(n_405), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_119), .A2(n_184), .B1(n_425), .B2(n_426), .Y(n_438) );
INVx1_ASAP7_75t_L g947 ( .A(n_120), .Y(n_947) );
INVx1_ASAP7_75t_L g654 ( .A(n_121), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_122), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_124), .A2(n_235), .B1(n_336), .B2(n_339), .Y(n_732) );
OAI22xp33_ASAP7_75t_SL g780 ( .A1(n_125), .A2(n_127), .B1(n_633), .B2(n_636), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_125), .A2(n_134), .B1(n_738), .B2(n_739), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g1326 ( .A1(n_126), .A2(n_1327), .B1(n_1384), .B2(n_1386), .C1(n_1389), .C2(n_1391), .Y(n_1326) );
XNOR2xp5_ASAP7_75t_L g1329 ( .A(n_126), .B(n_1330), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_128), .A2(n_238), .B1(n_1128), .B2(n_1129), .Y(n_1152) );
INVx1_ASAP7_75t_L g1097 ( .A(n_129), .Y(n_1097) );
AOI22xp5_ASAP7_75t_L g1133 ( .A1(n_131), .A2(n_132), .B1(n_1123), .B2(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g670 ( .A(n_133), .Y(n_670) );
INVx1_ASAP7_75t_L g779 ( .A(n_134), .Y(n_779) );
INVx1_ASAP7_75t_L g945 ( .A(n_135), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_137), .A2(n_140), .B1(n_1128), .B2(n_1129), .Y(n_1141) );
CKINVDCx5p33_ASAP7_75t_R g1041 ( .A(n_138), .Y(n_1041) );
INVx1_ASAP7_75t_L g545 ( .A(n_139), .Y(n_545) );
INVx1_ASAP7_75t_L g801 ( .A(n_142), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_142), .A2(n_216), .B1(n_336), .B2(n_339), .Y(n_828) );
INVx1_ASAP7_75t_L g893 ( .A(n_143), .Y(n_893) );
INVx1_ASAP7_75t_L g962 ( .A(n_144), .Y(n_962) );
OAI211xp5_ASAP7_75t_L g966 ( .A1(n_144), .A2(n_474), .B(n_627), .C(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g794 ( .A(n_145), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_146), .Y(n_813) );
INVx1_ASAP7_75t_L g1356 ( .A(n_147), .Y(n_1356) );
BUFx3_ASAP7_75t_L g303 ( .A(n_149), .Y(n_303) );
OAI211xp5_ASAP7_75t_SL g776 ( .A1(n_150), .A2(n_613), .B(n_627), .C(n_777), .Y(n_776) );
OAI211xp5_ASAP7_75t_SL g784 ( .A1(n_150), .A2(n_507), .B(n_588), .C(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g939 ( .A(n_151), .Y(n_939) );
INVx1_ASAP7_75t_L g462 ( .A(n_152), .Y(n_462) );
INVx1_ASAP7_75t_L g942 ( .A(n_153), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_154), .Y(n_990) );
INVx1_ASAP7_75t_L g1081 ( .A(n_155), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_156), .A2(n_241), .B1(n_282), .B2(n_562), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_156), .A2(n_241), .B1(n_581), .B2(n_582), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_157), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_158), .A2(n_159), .B1(n_1128), .B2(n_1129), .Y(n_1156) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_160), .Y(n_961) );
XNOR2x1_ASAP7_75t_L g933 ( .A(n_161), .B(n_934), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_162), .A2(n_219), .B1(n_1123), .B2(n_1134), .Y(n_1160) );
OAI22xp33_ASAP7_75t_L g1050 ( .A1(n_163), .A2(n_261), .B1(n_336), .B2(n_339), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_164), .Y(n_1029) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_165), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_166), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_167), .Y(n_807) );
INVx1_ASAP7_75t_L g554 ( .A(n_168), .Y(n_554) );
INVx1_ASAP7_75t_L g874 ( .A(n_169), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_170), .Y(n_1021) );
INVx1_ASAP7_75t_L g1359 ( .A(n_172), .Y(n_1359) );
INVx1_ASAP7_75t_L g573 ( .A(n_173), .Y(n_573) );
OAI211xp5_ASAP7_75t_L g583 ( .A1(n_173), .A2(n_584), .B(n_588), .C(n_589), .Y(n_583) );
INVx1_ASAP7_75t_L g1086 ( .A(n_174), .Y(n_1086) );
INVx1_ASAP7_75t_L g1062 ( .A(n_176), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_177), .Y(n_707) );
INVx1_ASAP7_75t_L g486 ( .A(n_178), .Y(n_486) );
INVx1_ASAP7_75t_L g862 ( .A(n_179), .Y(n_862) );
INVx1_ASAP7_75t_L g1346 ( .A(n_181), .Y(n_1346) );
INVx1_ASAP7_75t_L g806 ( .A(n_182), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_182), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g308 ( .A(n_183), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_184), .A2(n_191), .B1(n_397), .B2(n_400), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_186), .B(n_325), .Y(n_873) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_186), .Y(n_881) );
OAI211xp5_ASAP7_75t_SL g1058 ( .A1(n_187), .A2(n_588), .B(n_1059), .C(n_1060), .Y(n_1058) );
INVx1_ASAP7_75t_L g1073 ( .A(n_187), .Y(n_1073) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_188), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_189), .Y(n_1025) );
OAI211xp5_ASAP7_75t_L g723 ( .A1(n_190), .A2(n_613), .B(n_627), .C(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g740 ( .A(n_190), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_191), .A2(n_247), .B1(n_425), .B2(n_426), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_192), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g1064 ( .A1(n_193), .A2(n_254), .B1(n_1065), .B2(n_1066), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_193), .A2(n_254), .B1(n_575), .B2(n_1075), .Y(n_1074) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_194), .Y(n_286) );
INVx1_ASAP7_75t_L g1042 ( .A(n_197), .Y(n_1042) );
OAI211xp5_ASAP7_75t_L g1047 ( .A1(n_197), .A2(n_641), .B(n_1010), .C(n_1048), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_198), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_199), .Y(n_978) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_200), .A2(n_250), .B1(n_432), .B2(n_433), .C(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g857 ( .A(n_201), .Y(n_857) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_204), .A2(n_564), .B(n_568), .C(n_570), .Y(n_563) );
INVx1_ASAP7_75t_L g594 ( .A(n_204), .Y(n_594) );
INVx1_ASAP7_75t_L g665 ( .A(n_205), .Y(n_665) );
INVx1_ASAP7_75t_L g944 ( .A(n_206), .Y(n_944) );
INVxp67_ASAP7_75t_SL g883 ( .A(n_207), .Y(n_883) );
INVx1_ASAP7_75t_L g1339 ( .A(n_208), .Y(n_1339) );
OAI211xp5_ASAP7_75t_L g1380 ( .A1(n_208), .A2(n_588), .B(n_1059), .C(n_1381), .Y(n_1380) );
XNOR2xp5_ASAP7_75t_L g1387 ( .A(n_209), .B(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g895 ( .A(n_210), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_211), .Y(n_1003) );
INVx1_ASAP7_75t_L g660 ( .A(n_213), .Y(n_660) );
XOR2xp5_ASAP7_75t_L g744 ( .A(n_214), .B(n_745), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_215), .Y(n_763) );
INVx1_ASAP7_75t_L g803 ( .A(n_216), .Y(n_803) );
BUFx3_ASAP7_75t_L g290 ( .A(n_217), .Y(n_290) );
INVx1_ASAP7_75t_L g358 ( .A(n_217), .Y(n_358) );
XOR2x2_ASAP7_75t_L g1053 ( .A(n_220), .B(n_1054), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_221), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_223), .Y(n_754) );
INVx1_ASAP7_75t_L g851 ( .A(n_224), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_225), .A2(n_250), .B1(n_913), .B2(n_914), .Y(n_912) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_226), .A2(n_627), .B(n_1001), .C(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1049 ( .A(n_226), .Y(n_1049) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_227), .Y(n_473) );
INVx1_ASAP7_75t_L g652 ( .A(n_228), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_229), .Y(n_986) );
INVx1_ASAP7_75t_L g1094 ( .A(n_230), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_231), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_232), .A2(n_626), .B(n_627), .C(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g644 ( .A(n_232), .Y(n_644) );
INVx1_ASAP7_75t_L g350 ( .A(n_233), .Y(n_350) );
INVx2_ASAP7_75t_L g412 ( .A(n_233), .Y(n_412) );
INVx1_ASAP7_75t_L g443 ( .A(n_233), .Y(n_443) );
INVx1_ASAP7_75t_L g458 ( .A(n_234), .Y(n_458) );
INVx1_ASAP7_75t_L g948 ( .A(n_237), .Y(n_948) );
XNOR2x1_ASAP7_75t_L g537 ( .A(n_239), .B(n_538), .Y(n_537) );
XNOR2xp5_ASAP7_75t_L g889 ( .A(n_240), .B(n_890), .Y(n_889) );
XNOR2xp5_ASAP7_75t_L g451 ( .A(n_242), .B(n_452), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_243), .Y(n_712) );
INVx1_ASAP7_75t_L g1353 ( .A(n_244), .Y(n_1353) );
INVx1_ASAP7_75t_L g861 ( .A(n_245), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_246), .Y(n_899) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_248), .Y(n_612) );
INVx1_ASAP7_75t_L g337 ( .A(n_249), .Y(n_337) );
INVx1_ASAP7_75t_L g546 ( .A(n_251), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g815 ( .A1(n_252), .A2(n_416), .B(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g834 ( .A(n_252), .Y(n_834) );
INVx1_ASAP7_75t_L g1096 ( .A(n_255), .Y(n_1096) );
XNOR2xp5_ASAP7_75t_L g1016 ( .A(n_256), .B(n_1017), .Y(n_1016) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_257), .A2(n_261), .B1(n_354), .B2(n_485), .Y(n_1043) );
INVx1_ASAP7_75t_L g1063 ( .A(n_258), .Y(n_1063) );
OAI211xp5_ASAP7_75t_L g1070 ( .A1(n_258), .A2(n_564), .B(n_568), .C(n_1071), .Y(n_1070) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_259), .Y(n_991) );
OAI211xp5_ASAP7_75t_L g1333 ( .A1(n_262), .A2(n_1334), .B(n_1335), .C(n_1336), .Y(n_1333) );
INVx1_ASAP7_75t_L g1382 ( .A(n_262), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_264), .Y(n_799) );
OAI211xp5_ASAP7_75t_L g958 ( .A1(n_265), .A2(n_641), .B(n_959), .C(n_960), .Y(n_958) );
INVx1_ASAP7_75t_L g968 ( .A(n_265), .Y(n_968) );
INVx1_ASAP7_75t_L g1354 ( .A(n_266), .Y(n_1354) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_291), .B(n_1109), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_276), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g1385 ( .A(n_270), .B(n_279), .Y(n_1385) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g1390 ( .A(n_272), .B(n_275), .Y(n_1390) );
INVx1_ASAP7_75t_L g1392 ( .A(n_272), .Y(n_1392) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g1395 ( .A(n_275), .B(n_1392), .Y(n_1395) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g391 ( .A(n_279), .B(n_392), .Y(n_391) );
AOI21xp5_ASAP7_75t_SL g790 ( .A1(n_279), .A2(n_791), .B(n_804), .Y(n_790) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g419 ( .A(n_280), .B(n_290), .Y(n_419) );
AND2x4_ASAP7_75t_L g817 ( .A(n_280), .B(n_289), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_281), .A2(n_356), .B1(n_499), .B2(n_500), .Y(n_498) );
AND2x4_ASAP7_75t_SL g1384 ( .A(n_281), .B(n_1385), .Y(n_1384) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x6_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
OR2x6_ASAP7_75t_L g576 ( .A(n_283), .B(n_357), .Y(n_576) );
BUFx4f_ASAP7_75t_L g601 ( .A(n_283), .Y(n_601) );
OR2x2_ASAP7_75t_L g633 ( .A(n_283), .B(n_357), .Y(n_633) );
INVx1_ASAP7_75t_L g690 ( .A(n_283), .Y(n_690) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g355 ( .A(n_284), .Y(n_355) );
BUFx4f_ASAP7_75t_L g678 ( .A(n_284), .Y(n_678) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g359 ( .A(n_286), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g365 ( .A(n_286), .B(n_287), .Y(n_365) );
INVx1_ASAP7_75t_L g375 ( .A(n_286), .Y(n_375) );
INVx2_ASAP7_75t_L g383 ( .A(n_286), .Y(n_383) );
INVx2_ASAP7_75t_L g389 ( .A(n_286), .Y(n_389) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_286), .B(n_287), .Y(n_461) );
INVx2_ASAP7_75t_L g360 ( .A(n_287), .Y(n_360) );
BUFx2_ASAP7_75t_L g371 ( .A(n_287), .Y(n_371) );
INVx1_ASAP7_75t_L g384 ( .A(n_287), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_287), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g406 ( .A(n_287), .B(n_389), .Y(n_406) );
OR2x2_ASAP7_75t_L g457 ( .A(n_287), .B(n_383), .Y(n_457) );
OR2x6_ASAP7_75t_L g354 ( .A(n_288), .B(n_355), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_288), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_798) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g377 ( .A(n_289), .Y(n_377) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g370 ( .A(n_290), .Y(n_370) );
AND2x4_ASAP7_75t_L g373 ( .A(n_290), .B(n_374), .Y(n_373) );
XNOR2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_694), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_621), .B1(n_692), .B2(n_693), .Y(n_292) );
INVx1_ASAP7_75t_L g693 ( .A(n_293), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B1(n_449), .B2(n_620), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_342), .B1(n_351), .B2(n_390), .C(n_394), .Y(n_296) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_315), .C(n_333), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_308), .B2(n_309), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_299), .A2(n_308), .B1(n_353), .B2(n_356), .Y(n_352) );
INVx2_ASAP7_75t_SL g581 ( .A(n_300), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_300), .A2(n_743), .B1(n_893), .B2(n_895), .Y(n_905) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_SL g509 ( .A(n_301), .Y(n_509) );
INVx1_ASAP7_75t_L g830 ( .A(n_301), .Y(n_830) );
OR2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_306), .Y(n_301) );
OR2x4_ASAP7_75t_L g336 ( .A(n_302), .B(n_310), .Y(n_336) );
BUFx4f_ASAP7_75t_L g653 ( .A(n_302), .Y(n_653) );
INVx2_ASAP7_75t_L g989 ( .A(n_302), .Y(n_989) );
BUFx3_ASAP7_75t_L g1082 ( .A(n_302), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1349 ( .A(n_302), .Y(n_1349) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g314 ( .A(n_303), .Y(n_314) );
AND2x4_ASAP7_75t_L g318 ( .A(n_303), .B(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_303), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_303), .B(n_320), .Y(n_341) );
INVx1_ASAP7_75t_L g436 ( .A(n_304), .Y(n_436) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_L g313 ( .A(n_305), .Y(n_313) );
INVx1_ASAP7_75t_L g310 ( .A(n_306), .Y(n_310) );
AND2x4_ASAP7_75t_L g332 ( .A(n_306), .B(n_318), .Y(n_332) );
OR2x6_ASAP7_75t_L g339 ( .A(n_306), .B(n_340), .Y(n_339) );
NAND3x1_ASAP7_75t_L g441 ( .A(n_306), .B(n_442), .C(n_444), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_306), .B(n_444), .Y(n_674) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g325 ( .A(n_307), .Y(n_325) );
NAND2xp33_ASAP7_75t_SL g526 ( .A(n_307), .B(n_345), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_309), .A2(n_499), .B1(n_500), .B2(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g582 ( .A(n_309), .Y(n_582) );
INVx1_ASAP7_75t_L g639 ( .A(n_309), .Y(n_639) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g743 ( .A(n_310), .B(n_311), .Y(n_743) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_311), .Y(n_425) );
INVx2_ASAP7_75t_L g518 ( .A(n_311), .Y(n_518) );
INVx2_ASAP7_75t_L g528 ( .A(n_311), .Y(n_528) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g544 ( .A(n_312), .Y(n_544) );
BUFx8_ASAP7_75t_L g659 ( .A(n_312), .Y(n_659) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_312), .Y(n_711) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x4_ASAP7_75t_L g435 ( .A(n_314), .B(n_436), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_321), .C(n_332), .Y(n_315) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g432 ( .A(n_318), .Y(n_432) );
INVx2_ASAP7_75t_L g505 ( .A(n_318), .Y(n_505) );
BUFx2_ASAP7_75t_L g523 ( .A(n_318), .Y(n_523) );
BUFx2_ASAP7_75t_L g557 ( .A(n_318), .Y(n_557) );
BUFx2_ASAP7_75t_L g837 ( .A(n_318), .Y(n_837) );
INVx1_ASAP7_75t_L g428 ( .A(n_319), .Y(n_428) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_323), .A2(n_736), .B1(n_778), .B2(n_786), .Y(n_785) );
AOI222xp33_ASAP7_75t_L g872 ( .A1(n_323), .A2(n_329), .B1(n_523), .B2(n_873), .C1(n_874), .C2(n_875), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_323), .B(n_899), .Y(n_908) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_323), .A2(n_329), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_323), .A2(n_329), .B1(n_1003), .B2(n_1014), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_323), .A2(n_329), .B1(n_1041), .B2(n_1049), .Y(n_1048) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
AND2x2_ASAP7_75t_L g329 ( .A(n_324), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g591 ( .A(n_324), .B(n_326), .Y(n_591) );
AND2x4_ASAP7_75t_L g593 ( .A(n_324), .B(n_330), .Y(n_593) );
AND2x4_ASAP7_75t_L g643 ( .A(n_324), .B(n_326), .Y(n_643) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND3x4_ASAP7_75t_L g429 ( .A(n_325), .B(n_345), .C(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g736 ( .A(n_325), .B(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g427 ( .A(n_327), .B(n_428), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_327), .B(n_331), .Y(n_587) );
INVx2_ASAP7_75t_L g739 ( .A(n_327), .Y(n_739) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_L g507 ( .A(n_329), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_329), .A2(n_629), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI32xp33_ASAP7_75t_L g735 ( .A1(n_329), .A2(n_726), .A3(n_736), .B1(n_738), .B2(n_740), .Y(n_735) );
INVxp67_ASAP7_75t_L g827 ( .A(n_329), .Y(n_827) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI211xp5_ASAP7_75t_L g503 ( .A1(n_332), .A2(n_491), .B(n_504), .C(n_506), .Y(n_503) );
CKINVDCx8_ASAP7_75t_R g588 ( .A(n_332), .Y(n_588) );
CKINVDCx8_ASAP7_75t_R g641 ( .A(n_332), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g824 ( .A(n_332), .B(n_825), .C(n_828), .Y(n_824) );
NOR3xp33_ASAP7_75t_L g906 ( .A(n_332), .B(n_907), .C(n_909), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_337), .B2(n_338), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_334), .A2(n_337), .B1(n_380), .B2(n_385), .Y(n_379) );
INVx2_ASAP7_75t_L g597 ( .A(n_335), .Y(n_597) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g512 ( .A(n_336), .Y(n_512) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_336), .Y(n_1065) );
INVx1_ASAP7_75t_L g596 ( .A(n_338), .Y(n_596) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g513 ( .A(n_339), .Y(n_513) );
INVx1_ASAP7_75t_L g1067 ( .A(n_339), .Y(n_1067) );
BUFx3_ASAP7_75t_L g519 ( .A(n_340), .Y(n_519) );
INVx1_ASAP7_75t_L g662 ( .A(n_340), .Y(n_662) );
BUFx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g531 ( .A(n_341), .Y(n_531) );
OAI31xp33_ASAP7_75t_L g579 ( .A1(n_342), .A2(n_580), .A3(n_583), .B(n_595), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_342), .A2(n_823), .B(n_832), .Y(n_822) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_342), .Y(n_1068) );
OAI31xp33_ASAP7_75t_L g1378 ( .A1(n_342), .A2(n_1379), .A3(n_1380), .B(n_1383), .Y(n_1378) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_343), .B(n_346), .Y(n_342) );
AND2x2_ASAP7_75t_L g515 ( .A(n_343), .B(n_346), .Y(n_515) );
AND2x2_ASAP7_75t_L g648 ( .A(n_343), .B(n_346), .Y(n_648) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g421 ( .A(n_348), .Y(n_421) );
OR2x2_ASAP7_75t_L g525 ( .A(n_348), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_348), .B(n_419), .Y(n_687) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_361), .C(n_379), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g894 ( .A(n_354), .Y(n_894) );
BUFx3_ASAP7_75t_L g616 ( .A(n_355), .Y(n_616) );
BUFx3_ASAP7_75t_L g766 ( .A(n_355), .Y(n_766) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_355), .Y(n_869) );
CKINVDCx16_ASAP7_75t_R g562 ( .A(n_356), .Y(n_562) );
INVx4_ASAP7_75t_L g636 ( .A(n_356), .Y(n_636) );
INVx3_ASAP7_75t_SL g792 ( .A(n_356), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_356), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_892) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g399 ( .A(n_359), .Y(n_399) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_359), .Y(n_417) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B(n_367), .C(n_376), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_362), .B(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g918 ( .A(n_363), .Y(n_918) );
INVx1_ASAP7_75t_L g920 ( .A(n_363), .Y(n_920) );
BUFx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g378 ( .A(n_364), .Y(n_378) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_369), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_369), .A2(n_631), .B1(n_778), .B2(n_779), .Y(n_777) );
BUFx3_ASAP7_75t_L g1337 ( .A(n_369), .Y(n_1337) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g380 ( .A(n_370), .B(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g386 ( .A(n_370), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g572 ( .A(n_370), .B(n_371), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g793 ( .A1(n_370), .A2(n_794), .B(n_795), .C(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g800 ( .A(n_370), .Y(n_800) );
AND2x2_ASAP7_75t_L g490 ( .A(n_371), .B(n_377), .Y(n_490) );
INVx2_ASAP7_75t_L g1072 ( .A(n_372), .Y(n_1072) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g493 ( .A(n_373), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_373), .A2(n_571), .B1(n_572), .B2(n_573), .Y(n_570) );
BUFx3_ASAP7_75t_L g631 ( .A(n_373), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_373), .A2(n_490), .B1(n_899), .B2(n_900), .Y(n_898) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g497 ( .A(n_376), .Y(n_497) );
INVx2_ASAP7_75t_L g627 ( .A(n_376), .Y(n_627) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g569 ( .A(n_377), .B(n_401), .Y(n_569) );
OR2x2_ASAP7_75t_L g634 ( .A(n_377), .B(n_387), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_380), .A2(n_483), .B1(n_484), .B2(n_486), .C(n_487), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_380), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g404 ( .A(n_382), .Y(n_404) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g577 ( .A(n_385), .Y(n_577) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g485 ( .A(n_386), .Y(n_485) );
INVx1_ASAP7_75t_L g729 ( .A(n_386), .Y(n_729) );
INVx8_ASAP7_75t_L g605 ( .A(n_387), .Y(n_605) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI31xp33_ASAP7_75t_SL g624 ( .A1(n_390), .A2(n_625), .A3(n_632), .B(n_635), .Y(n_624) );
BUFx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g501 ( .A(n_391), .Y(n_501) );
BUFx2_ASAP7_75t_L g578 ( .A(n_391), .Y(n_578) );
OAI31xp33_ASAP7_75t_L g774 ( .A1(n_391), .A2(n_775), .A3(n_776), .B(n_780), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g878 ( .A1(n_391), .A2(n_879), .B(n_886), .Y(n_878) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_391), .Y(n_1077) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_414), .C(n_423), .D(n_437), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_402), .C(n_407), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_401), .Y(n_496) );
BUFx3_ASAP7_75t_L g795 ( .A(n_401), .Y(n_795) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
INVx2_ASAP7_75t_L g819 ( .A(n_404), .Y(n_819) );
INVx2_ASAP7_75t_SL g913 ( .A(n_404), .Y(n_913) );
INVx1_ASAP7_75t_L g922 ( .A(n_404), .Y(n_922) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g466 ( .A(n_406), .Y(n_466) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_406), .Y(n_479) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g911 ( .A(n_409), .Y(n_911) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g468 ( .A(n_410), .Y(n_468) );
INVx2_ASAP7_75t_L g680 ( .A(n_410), .Y(n_680) );
INVx2_ASAP7_75t_L g1099 ( .A(n_410), .Y(n_1099) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
OR2x2_ASAP7_75t_L g673 ( .A(n_411), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g821 ( .A(n_411), .Y(n_821) );
OR2x6_ASAP7_75t_L g863 ( .A(n_411), .B(n_674), .Y(n_863) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g430 ( .A(n_412), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .C(n_422), .Y(n_414) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g917 ( .A(n_417), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_418), .Y(n_618) );
INVx2_ASAP7_75t_L g1377 ( .A(n_418), .Y(n_1377) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_419), .B(n_420), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g808 ( .A1(n_419), .A2(n_609), .B1(n_809), .B2(n_810), .C(n_811), .Y(n_808) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_429), .C(n_431), .Y(n_423) );
INVx2_ASAP7_75t_SL g552 ( .A(n_425), .Y(n_552) );
BUFx12f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g839 ( .A(n_427), .Y(n_839) );
INVx1_ASAP7_75t_L g737 ( .A(n_428), .Y(n_737) );
INVx1_ASAP7_75t_L g932 ( .A(n_429), .Y(n_932) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_432), .Y(n_646) );
BUFx2_ASAP7_75t_L g556 ( .A(n_433), .Y(n_556) );
INVx8_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g522 ( .A(n_434), .Y(n_522) );
INVx2_ASAP7_75t_L g845 ( .A(n_434), .Y(n_845) );
INVx8_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g448 ( .A(n_435), .Y(n_448) );
BUFx3_ASAP7_75t_L g836 ( .A(n_435), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .C(n_445), .Y(n_437) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g535 ( .A(n_440), .Y(n_535) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g559 ( .A(n_441), .Y(n_559) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
INVx1_ASAP7_75t_L g620 ( .A(n_449), .Y(n_620) );
OA22x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_536), .B1(n_537), .B2(n_619), .Y(n_449) );
INVx1_ASAP7_75t_L g619 ( .A(n_450), .Y(n_619) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_481), .C(n_502), .D(n_516), .Y(n_452) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_467), .B1(n_469), .B2(n_480), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B1(n_459), .B2(n_462), .C(n_463), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_455), .A2(n_474), .B1(n_852), .B2(n_862), .Y(n_867) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g682 ( .A(n_456), .Y(n_682) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g472 ( .A(n_457), .Y(n_472) );
INVx2_ASAP7_75t_L g611 ( .A(n_457), .Y(n_611) );
BUFx3_ASAP7_75t_L g771 ( .A(n_457), .Y(n_771) );
BUFx2_ASAP7_75t_L g953 ( .A(n_457), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_458), .A2(n_518), .B1(n_519), .B2(n_520), .C(n_521), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_459), .A2(n_682), .B1(n_754), .B2(n_758), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_459), .A2(n_938), .B1(n_947), .B2(n_953), .Y(n_952) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_460), .Y(n_474) );
BUFx4f_ASAP7_75t_L g613 ( .A(n_460), .Y(n_613) );
INVx4_ASAP7_75t_L g684 ( .A(n_460), .Y(n_684) );
BUFx4f_ASAP7_75t_L g814 ( .A(n_460), .Y(n_814) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g567 ( .A(n_461), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_462), .A2(n_528), .B1(n_529), .B2(n_532), .C(n_533), .Y(n_527) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g914 ( .A(n_466), .Y(n_914) );
OA33x2_ASAP7_75t_L g598 ( .A1(n_467), .A2(n_599), .A3(n_606), .B1(n_608), .B2(n_615), .B3(n_618), .Y(n_598) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI33xp33_ASAP7_75t_L g764 ( .A1(n_468), .A2(n_686), .A3(n_765), .B1(n_769), .B2(n_770), .B3(n_773), .Y(n_764) );
OAI33xp33_ASAP7_75t_L g1019 ( .A1(n_468), .A2(n_998), .A3(n_1020), .B1(n_1024), .B2(n_1027), .B3(n_1030), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g1364 ( .A1(n_468), .A2(n_1365), .A3(n_1366), .B1(n_1369), .B2(n_1373), .B3(n_1377), .Y(n_1364) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .B1(n_474), .B2(n_475), .C(n_476), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_470), .A2(n_545), .B1(n_553), .B2(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_470), .A2(n_1353), .B1(n_1356), .B2(n_1367), .Y(n_1366) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_474), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_474), .A2(n_995), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_498), .B(n_501), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_483), .A2(n_486), .B1(n_511), .B2(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g1075 ( .A(n_484), .Y(n_1075) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g1342 ( .A(n_485), .Y(n_1342) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .C(n_497), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_488) );
INVx1_ASAP7_75t_L g797 ( .A(n_490), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g1002 ( .A1(n_490), .A2(n_492), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_490), .A2(n_631), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_492), .A2(n_572), .B1(n_725), .B2(n_726), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_492), .A2(n_572), .B1(n_961), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_492), .A2(n_1337), .B1(n_1338), .B2(n_1339), .Y(n_1336) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_497), .B(n_898), .C(n_901), .Y(n_897) );
AO21x1_ASAP7_75t_L g891 ( .A1(n_501), .A2(n_892), .B(n_896), .Y(n_891) );
AOI31xp33_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_508), .A3(n_510), .B(n_514), .Y(n_502) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g928 ( .A(n_505), .Y(n_928) );
INVx2_ASAP7_75t_L g1057 ( .A(n_509), .Y(n_1057) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g877 ( .A(n_513), .Y(n_877) );
AO21x1_ASAP7_75t_L g904 ( .A1(n_514), .A2(n_905), .B(n_906), .Y(n_904) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_524), .B1(n_527), .B2(n_534), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_519), .A2(n_542), .B1(n_545), .B2(n_546), .C(n_547), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_519), .A2(n_552), .B1(n_553), .B2(n_554), .C(n_555), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_519), .A2(n_1091), .B1(n_1093), .B2(n_1094), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_519), .A2(n_528), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
OAI22xp5_ASAP7_75t_L g1355 ( .A1(n_519), .A2(n_1356), .B1(n_1357), .B2(n_1359), .Y(n_1355) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_524), .A2(n_833), .B1(n_840), .B2(n_841), .Y(n_832) );
OAI33xp33_ASAP7_75t_L g849 ( .A1(n_524), .A2(n_850), .A3(n_853), .B1(n_856), .B2(n_860), .B3(n_863), .Y(n_849) );
OAI33xp33_ASAP7_75t_L g1079 ( .A1(n_524), .A2(n_840), .A3(n_1080), .B1(n_1085), .B2(n_1090), .B3(n_1095), .Y(n_1079) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx4f_ASAP7_75t_L g550 ( .A(n_525), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_528), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_528), .A2(n_756), .B1(n_981), .B2(n_982), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_528), .A2(n_756), .B1(n_1025), .B2(n_1031), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_529), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_529), .A2(n_710), .B1(n_938), .B2(n_939), .Y(n_937) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g756 ( .A(n_530), .Y(n_756) );
CKINVDCx8_ASAP7_75t_R g843 ( .A(n_530), .Y(n_843) );
INVx3_ASAP7_75t_L g858 ( .A(n_530), .Y(n_858) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g667 ( .A(n_531), .Y(n_667) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND4xp75_ASAP7_75t_L g538 ( .A(n_539), .B(n_560), .C(n_579), .D(n_598), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_549), .B1(n_551), .B2(n_558), .Y(n_540) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g985 ( .A(n_543), .Y(n_985) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g842 ( .A(n_544), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_546), .A2(n_554), .B1(n_616), .B2(n_617), .Y(n_615) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI33xp33_ASAP7_75t_L g650 ( .A1(n_550), .A2(n_651), .A3(n_656), .B1(n_663), .B2(n_669), .B3(n_673), .Y(n_650) );
OAI33xp33_ASAP7_75t_L g702 ( .A1(n_550), .A2(n_673), .A3(n_703), .B1(n_706), .B2(n_709), .B3(n_714), .Y(n_702) );
OAI33xp33_ASAP7_75t_L g747 ( .A1(n_550), .A2(n_673), .A3(n_748), .B1(n_753), .B2(n_757), .B3(n_761), .Y(n_747) );
OAI33xp33_ASAP7_75t_L g936 ( .A1(n_550), .A2(n_673), .A3(n_937), .B1(n_940), .B2(n_943), .B3(n_946), .Y(n_936) );
OAI33xp33_ASAP7_75t_L g976 ( .A1(n_550), .A2(n_673), .A3(n_977), .B1(n_980), .B2(n_983), .B3(n_987), .Y(n_976) );
OAI33xp33_ASAP7_75t_L g1033 ( .A1(n_550), .A2(n_673), .A3(n_1034), .B1(n_1035), .B2(n_1036), .B3(n_1037), .Y(n_1033) );
OAI33xp33_ASAP7_75t_L g1344 ( .A1(n_550), .A2(n_1345), .A3(n_1352), .B1(n_1355), .B2(n_1360), .B3(n_1361), .Y(n_1344) );
OAI211xp5_ASAP7_75t_L g833 ( .A1(n_552), .A2(n_834), .B(n_835), .C(n_838), .Y(n_833) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_559), .Y(n_840) );
INVx2_ASAP7_75t_L g1360 ( .A(n_559), .Y(n_1360) );
OAI31xp33_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .A3(n_574), .B(n_578), .Y(n_560) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g1334 ( .A(n_566), .Y(n_1334) );
BUFx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_SL g607 ( .A(n_567), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_567), .A2(n_654), .B1(n_672), .B2(n_682), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_567), .A2(n_953), .B1(n_979), .B2(n_991), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_567), .A2(n_995), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1368 ( .A(n_567), .Y(n_1368) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g1335 ( .A(n_569), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_571), .A2(n_590), .B1(n_592), .B2(n_594), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g880 ( .A1(n_572), .A2(n_631), .B1(n_795), .B2(n_874), .C1(n_875), .C2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_572), .A2(n_1062), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g1341 ( .A(n_576), .Y(n_1341) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_578), .A2(n_723), .A3(n_727), .B(n_730), .Y(n_722) );
OAI31xp33_ASAP7_75t_SL g964 ( .A1(n_578), .A2(n_965), .A3(n_966), .B(n_969), .Y(n_964) );
OAI31xp33_ASAP7_75t_L g999 ( .A1(n_578), .A2(n_1000), .A3(n_1005), .B(n_1006), .Y(n_999) );
OAI31xp33_ASAP7_75t_L g1038 ( .A1(n_578), .A2(n_1039), .A3(n_1043), .B(n_1044), .Y(n_1038) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g826 ( .A(n_585), .Y(n_826) );
INVx2_ASAP7_75t_L g1059 ( .A(n_585), .Y(n_1059) );
INVx1_ASAP7_75t_L g1351 ( .A(n_585), .Y(n_1351) );
INVx4_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_586), .Y(n_655) );
INVx3_ASAP7_75t_L g751 ( .A(n_586), .Y(n_751) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx3_ASAP7_75t_L g671 ( .A(n_587), .Y(n_671) );
BUFx2_ASAP7_75t_L g1012 ( .A(n_587), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_590), .A2(n_592), .B1(n_1338), .B2(n_1382), .Y(n_1381) );
BUFx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_591), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_592), .A2(n_1061), .B1(n_1062), .B2(n_1063), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B1(n_602), .B2(n_603), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_601), .A2(n_603), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx5_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx6_ASAP7_75t_L g617 ( .A(n_604), .Y(n_617) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g679 ( .A(n_605), .Y(n_679) );
INVx4_ASAP7_75t_L g691 ( .A(n_605), .Y(n_691) );
INVx2_ASAP7_75t_L g768 ( .A(n_605), .Y(n_768) );
INVx1_ASAP7_75t_L g951 ( .A(n_605), .Y(n_951) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_605), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_609), .A2(n_1086), .B1(n_1093), .B2(n_1105), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_609), .A2(n_1001), .B1(n_1083), .B2(n_1097), .Y(n_1106) );
INVx4_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g995 ( .A(n_611), .Y(n_995) );
INVx2_ASAP7_75t_L g1372 ( .A(n_611), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_613), .A2(n_771), .B1(n_854), .B2(n_857), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_617), .A2(n_1081), .B1(n_1096), .B2(n_1101), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_617), .A2(n_1089), .B1(n_1094), .B2(n_1101), .Y(n_1107) );
OAI33xp33_ASAP7_75t_L g1098 ( .A1(n_618), .A2(n_1099), .A3(n_1100), .B1(n_1104), .B2(n_1106), .B3(n_1107), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g692 ( .A(n_622), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_637), .C(n_649), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g879 ( .A(n_627), .B(n_880), .C(n_882), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_630), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g885 ( .A(n_634), .Y(n_885) );
OAI31xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .A3(n_647), .B(n_648), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .C(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g734 ( .A(n_643), .Y(n_734) );
OAI31xp33_ASAP7_75t_SL g731 ( .A1(n_648), .A2(n_732), .A3(n_733), .B(n_741), .Y(n_731) );
OAI31xp33_ASAP7_75t_SL g781 ( .A1(n_648), .A2(n_782), .A3(n_783), .B(n_784), .Y(n_781) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_648), .A2(n_871), .B(n_876), .Y(n_870) );
OAI31xp33_ASAP7_75t_L g956 ( .A1(n_648), .A2(n_957), .A3(n_958), .B(n_963), .Y(n_956) );
OAI31xp33_ASAP7_75t_SL g1007 ( .A1(n_648), .A2(n_1008), .A3(n_1009), .B(n_1015), .Y(n_1007) );
OAI31xp33_ASAP7_75t_SL g1045 ( .A1(n_648), .A2(n_1046), .A3(n_1047), .B(n_1050), .Y(n_1045) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_675), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_652), .A2(n_670), .B1(n_677), .B2(n_679), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_653), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_653), .A2(n_655), .B1(n_704), .B2(n_705), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_653), .A2(n_671), .B1(n_715), .B2(n_716), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_653), .A2(n_749), .B1(n_750), .B2(n_752), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_653), .A2(n_671), .B1(n_762), .B2(n_763), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_653), .A2(n_826), .B1(n_851), .B2(n_852), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g860 ( .A1(n_653), .A2(n_655), .B1(n_861), .B2(n_862), .Y(n_860) );
OAI22xp5_ASAP7_75t_SL g940 ( .A1(n_653), .A2(n_750), .B1(n_941), .B2(n_942), .Y(n_940) );
OAI22xp33_ASAP7_75t_L g943 ( .A1(n_653), .A2(n_671), .B1(n_944), .B2(n_945), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_653), .A2(n_750), .B1(n_978), .B2(n_979), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_655), .A2(n_988), .B1(n_1021), .B2(n_1028), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_657), .A2(n_665), .B1(n_682), .B2(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_658), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_SL g664 ( .A(n_659), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_660), .A2(n_668), .B1(n_689), .B2(n_691), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_661), .A2(n_664), .B1(n_707), .B2(n_708), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_661), .A2(n_759), .B1(n_947), .B2(n_948), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_661), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_666), .B2(n_668), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_666), .A2(n_710), .B1(n_712), .B2(n_713), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_666), .A2(n_842), .B1(n_854), .B2(n_855), .Y(n_853) );
BUFx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx6f_ASAP7_75t_L g959 ( .A(n_671), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_671), .A2(n_988), .B1(n_990), .B2(n_991), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_671), .A2(n_988), .B1(n_1023), .B2(n_1029), .Y(n_1037) );
OAI33xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_680), .A3(n_681), .B1(n_685), .B2(n_686), .B3(n_688), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_677), .A2(n_691), .B1(n_704), .B2(n_715), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g950 ( .A1(n_677), .A2(n_941), .B1(n_944), .B2(n_951), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_677), .A2(n_691), .B1(n_939), .B2(n_948), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_677), .A2(n_767), .B1(n_978), .B2(n_990), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_677), .A2(n_691), .B1(n_982), .B2(n_986), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_677), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_677), .A2(n_767), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
INVx4_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g1103 ( .A(n_678), .Y(n_1103) );
BUFx6f_ASAP7_75t_L g1375 ( .A(n_678), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_679), .A2(n_1101), .B1(n_1346), .B2(n_1362), .Y(n_1365) );
OAI33xp33_ASAP7_75t_L g717 ( .A1(n_680), .A2(n_686), .A3(n_718), .B1(n_719), .B2(n_720), .B3(n_721), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g864 ( .A1(n_680), .A2(n_686), .A3(n_865), .B1(n_866), .B2(n_867), .B3(n_868), .Y(n_864) );
OAI33xp33_ASAP7_75t_L g949 ( .A1(n_680), .A2(n_686), .A3(n_950), .B1(n_952), .B2(n_954), .B3(n_955), .Y(n_949) );
OAI33xp33_ASAP7_75t_L g992 ( .A1(n_680), .A2(n_993), .A3(n_994), .B1(n_996), .B2(n_997), .B3(n_998), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_682), .A2(n_683), .B1(n_707), .B2(n_712), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_682), .A2(n_683), .B1(n_705), .B2(n_716), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_682), .A2(n_683), .B1(n_942), .B2(n_945), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_683), .A2(n_981), .B1(n_984), .B2(n_995), .Y(n_994) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g772 ( .A(n_684), .Y(n_772) );
INVx1_ASAP7_75t_L g809 ( .A(n_684), .Y(n_809) );
INVx1_ASAP7_75t_L g1001 ( .A(n_684), .Y(n_1001) );
INVx2_ASAP7_75t_L g1105 ( .A(n_684), .Y(n_1105) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI33xp33_ASAP7_75t_L g910 ( .A1(n_687), .A2(n_911), .A3(n_912), .B1(n_915), .B2(n_919), .B3(n_921), .Y(n_910) );
INVx2_ASAP7_75t_L g998 ( .A(n_687), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_689), .A2(n_691), .B1(n_708), .B2(n_713), .Y(n_721) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_691), .A2(n_755), .B1(n_760), .B2(n_766), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_691), .A2(n_766), .B1(n_851), .B2(n_861), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_1052), .B2(n_1108), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_887), .Y(n_696) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_787), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_744), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_722), .C(n_731), .Y(n_700) );
NOR2xp33_ASAP7_75t_SL g701 ( .A(n_702), .B(n_717), .Y(n_701) );
INVx2_ASAP7_75t_L g1092 ( .A(n_710), .Y(n_1092) );
INVx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g759 ( .A(n_711), .Y(n_759) );
INVx2_ASAP7_75t_SL g926 ( .A(n_711), .Y(n_926) );
INVx5_ASAP7_75t_L g1088 ( .A(n_711), .Y(n_1088) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g802 ( .A(n_729), .B(n_803), .Y(n_802) );
INVx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_743), .A2(n_799), .B1(n_830), .B2(n_831), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_774), .C(n_781), .Y(n_745) );
NOR2xp33_ASAP7_75t_SL g746 ( .A(n_747), .B(n_764), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_749), .A2(n_762), .B1(n_766), .B2(n_767), .Y(n_765) );
INVx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g1084 ( .A(n_751), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_752), .A2(n_763), .B1(n_771), .B2(n_772), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_759), .A2(n_858), .B1(n_1026), .B2(n_1032), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_767), .A2(n_855), .B1(n_859), .B2(n_869), .Y(n_868) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
XOR2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_846), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_820), .B(n_822), .Y(n_789) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_808), .B(n_812), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g841 ( .A1(n_807), .A2(n_813), .B1(n_842), .B2(n_843), .C(n_844), .Y(n_841) );
OAI211xp5_ASAP7_75t_SL g812 ( .A1(n_813), .A2(n_814), .B(n_815), .C(n_818), .Y(n_812) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
BUFx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g823 ( .A(n_824), .B(n_829), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_843), .A2(n_1086), .B1(n_1087), .B2(n_1089), .Y(n_1085) );
NAND3xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_870), .C(n_878), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_864), .Y(n_848) );
INVx1_ASAP7_75t_L g929 ( .A(n_863), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_970), .B1(n_971), .B2(n_1051), .Y(n_887) );
INVx1_ASAP7_75t_L g1051 ( .A(n_888), .Y(n_1051) );
XNOR2x1_ASAP7_75t_SL g888 ( .A(n_889), .B(n_933), .Y(n_888) );
NAND4xp75_ASAP7_75t_L g890 ( .A(n_891), .B(n_904), .C(n_910), .D(n_923), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_903), .Y(n_896) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
AOI32xp33_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_927), .A3(n_929), .B1(n_930), .B2(n_931), .Y(n_923) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AND3x1_ASAP7_75t_L g934 ( .A(n_935), .B(n_956), .C(n_964), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_936), .B(n_949), .Y(n_935) );
BUFx3_ASAP7_75t_L g1376 ( .A(n_951), .Y(n_1376) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_959), .A2(n_1082), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
XNOR2x1_ASAP7_75t_L g971 ( .A(n_972), .B(n_1016), .Y(n_971) );
XNOR2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_974), .Y(n_972) );
AND3x1_ASAP7_75t_L g974 ( .A(n_975), .B(n_999), .C(n_1007), .Y(n_974) );
NOR2xp33_ASAP7_75t_SL g975 ( .A(n_976), .B(n_992), .Y(n_975) );
INVx2_ASAP7_75t_SL g988 ( .A(n_989), .Y(n_988) );
OAI22xp33_ASAP7_75t_L g1095 ( .A1(n_1010), .A2(n_1082), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
AND3x1_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1038), .C(n_1045), .Y(n_1017) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1033), .Y(n_1018) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1053), .Y(n_1108) );
NAND3xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1069), .C(n_1078), .Y(n_1054) );
OAI31xp33_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1058), .A3(n_1064), .B(n_1068), .Y(n_1055) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
OAI31xp33_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1074), .A3(n_1076), .B(n_1077), .Y(n_1069) );
OAI31xp33_ASAP7_75t_L g1331 ( .A1(n_1077), .A2(n_1332), .A3(n_1333), .B(n_1340), .Y(n_1331) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1098), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1080) );
BUFx3_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx8_ASAP7_75t_L g1358 ( .A(n_1088), .Y(n_1358) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_1103), .Y(n_1102) );
OAI21xp33_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1117), .B(n_1326), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g1110 ( .A(n_1111), .Y(n_1110) );
CKINVDCx5p33_ASAP7_75t_R g1111 ( .A(n_1112), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
AND2x6_ASAP7_75t_L g1123 ( .A(n_1113), .B(n_1124), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1113), .B(n_1126), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_1113), .B(n_1114), .Y(n_1128) );
AND2x6_ASAP7_75t_L g1129 ( .A(n_1113), .B(n_1130), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1113), .B(n_1126), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1113), .B(n_1126), .Y(n_1155) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_1114), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1116), .Y(n_1114) );
AND3x1_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1263), .C(n_1300), .Y(n_1117) );
AOI211xp5_ASAP7_75t_SL g1118 ( .A1(n_1119), .A2(n_1136), .B(n_1190), .C(n_1239), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1131), .Y(n_1120) );
INVx3_ASAP7_75t_L g1211 ( .A(n_1121), .Y(n_1211) );
A2O1A1Ixp33_ASAP7_75t_L g1229 ( .A1(n_1121), .A2(n_1230), .B(n_1231), .C(n_1232), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1121), .B(n_1189), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1127), .Y(n_1121) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1131), .Y(n_1202) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1131), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1131), .B(n_1171), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1131), .B(n_1238), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1131), .B(n_1153), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1277 ( .A(n_1131), .B(n_1247), .C(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1132), .B(n_1189), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1132), .B(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1132), .Y(n_1208) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1132), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1132), .B(n_1153), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1135), .Y(n_1132) );
OAI211xp5_ASAP7_75t_SL g1136 ( .A1(n_1137), .A2(n_1147), .B(n_1161), .C(n_1178), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1143), .Y(n_1138) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1139), .B(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1140), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1140), .B(n_1166), .Y(n_1175) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1140), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1140), .B(n_1165), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1140), .B(n_1144), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1140), .B(n_1143), .Y(n_1216) );
NAND2x1_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1143), .B(n_1174), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1143), .B(n_1183), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1143), .B(n_1186), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1143), .B(n_1175), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1143), .B(n_1205), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1143), .B(n_1223), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1143), .B(n_1164), .Y(n_1284) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1144), .B(n_1158), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1144), .B(n_1177), .Y(n_1176) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_1144), .A2(n_1179), .B1(n_1181), .B2(n_1185), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1144), .B(n_1169), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1245 ( .A(n_1144), .B(n_1246), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1144), .B(n_1165), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1144), .B(n_1205), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1144), .B(n_1166), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1144), .B(n_1166), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1146), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1157), .Y(n_1147) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1148), .Y(n_1238) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1148), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1153), .Y(n_1148) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1149), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1149), .B(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1150), .B(n_1153), .Y(n_1180) );
INVx2_ASAP7_75t_SL g1188 ( .A(n_1150), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1150), .B(n_1186), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1150), .B(n_1189), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1150), .B(n_1192), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1152), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_1153), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_1153), .A2(n_1164), .B1(n_1192), .B2(n_1195), .C(n_1199), .Y(n_1191) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1153), .A2(n_1166), .B1(n_1213), .B2(n_1217), .C(n_1220), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1153), .B(n_1158), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1153), .B(n_1320), .Y(n_1319) );
AND2x4_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1156), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1157), .B(n_1164), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1157), .B(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1157), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1157), .B(n_1257), .Y(n_1256) );
OAI211xp5_ASAP7_75t_L g1265 ( .A1(n_1157), .A2(n_1266), .B(n_1268), .C(n_1270), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1157), .B(n_1299), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1157), .B(n_1216), .Y(n_1318) );
CKINVDCx5p33_ASAP7_75t_R g1157 ( .A(n_1158), .Y(n_1157) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1158), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1158), .B(n_1202), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1158), .B(n_1197), .Y(n_1322) );
AND2x4_ASAP7_75t_SL g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g1161 ( .A1(n_1162), .A2(n_1171), .B1(n_1172), .B2(n_1176), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1171), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1170), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1164), .B(n_1234), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1169), .Y(n_1164) );
OAI322xp33_ASAP7_75t_L g1199 ( .A1(n_1165), .A2(n_1171), .A3(n_1200), .B1(n_1203), .B2(n_1205), .C1(n_1206), .C2(n_1209), .Y(n_1199) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1166), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1168), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1170), .B(n_1223), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1170), .B(n_1175), .Y(n_1286) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1171), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1171), .B(n_1269), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1171), .B(n_1286), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1171), .B(n_1181), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1171), .B(n_1202), .Y(n_1325) );
O2A1O1Ixp33_ASAP7_75t_L g1309 ( .A1(n_1172), .A2(n_1310), .B(n_1312), .C(n_1313), .Y(n_1309) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1174), .B(n_1194), .Y(n_1193) );
OAI22xp5_ASAP7_75t_SL g1301 ( .A1(n_1174), .A2(n_1206), .B1(n_1302), .B2(n_1303), .Y(n_1301) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1179), .B(n_1207), .Y(n_1206) );
AOI322xp5_ASAP7_75t_L g1227 ( .A1(n_1179), .A2(n_1201), .A3(n_1228), .B1(n_1229), .B2(n_1233), .C1(n_1235), .C2(n_1236), .Y(n_1227) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1181), .B(n_1186), .Y(n_1324) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1183), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1183), .B(n_1252), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1186), .B(n_1219), .Y(n_1218) );
CKINVDCx14_ASAP7_75t_R g1250 ( .A(n_1186), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1186), .B(n_1197), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1186), .B(n_1188), .Y(n_1278) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1187), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1189), .Y(n_1187) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1188), .Y(n_1197) );
A2O1A1Ixp33_ASAP7_75t_L g1282 ( .A1(n_1188), .A2(n_1283), .B(n_1285), .C(n_1287), .Y(n_1282) );
A2O1A1Ixp33_ASAP7_75t_L g1314 ( .A1(n_1188), .A2(n_1255), .B(n_1315), .C(n_1317), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1189), .B(n_1211), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1189), .B(n_1249), .Y(n_1248) );
OAI221xp5_ASAP7_75t_SL g1190 ( .A1(n_1191), .A2(n_1210), .B1(n_1212), .B2(n_1224), .C(n_1227), .Y(n_1190) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1194), .Y(n_1234) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1198), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_1197), .B(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1198), .Y(n_1232) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1204), .Y(n_1260) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1205), .Y(n_1247) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
CKINVDCx14_ASAP7_75t_R g1264 ( .A(n_1210), .Y(n_1264) );
OAI221xp5_ASAP7_75t_L g1288 ( .A1(n_1210), .A2(n_1289), .B1(n_1292), .B2(n_1293), .C(n_1294), .Y(n_1288) );
OAI31xp33_ASAP7_75t_SL g1300 ( .A1(n_1210), .A2(n_1301), .A3(n_1304), .B(n_1307), .Y(n_1300) );
CKINVDCx14_ASAP7_75t_R g1210 ( .A(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1211), .B(n_1226), .Y(n_1225) );
AOI322xp5_ASAP7_75t_L g1244 ( .A1(n_1213), .A2(n_1245), .A3(n_1248), .B1(n_1250), .B2(n_1251), .C1(n_1254), .C2(n_1256), .Y(n_1244) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1219), .B(n_1222), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1219), .B(n_1290), .Y(n_1293) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1246 ( .A(n_1223), .B(n_1247), .Y(n_1246) );
CKINVDCx14_ASAP7_75t_R g1224 ( .A(n_1225), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1226), .B(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1228), .Y(n_1321) );
OAI211xp5_ASAP7_75t_SL g1307 ( .A1(n_1232), .A2(n_1308), .B(n_1309), .C(n_1323), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1234), .B(n_1247), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1303 ( .A(n_1235), .B(n_1275), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1235), .B(n_1242), .Y(n_1306) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
OAI211xp5_ASAP7_75t_SL g1239 ( .A1(n_1240), .A2(n_1241), .B(n_1244), .C(n_1258), .Y(n_1239) );
INVxp67_ASAP7_75t_SL g1287 ( .A(n_1240), .Y(n_1287) );
INVxp67_ASAP7_75t_L g1269 ( .A(n_1241), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1243), .Y(n_1241) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1243), .Y(n_1275) );
AOI221xp5_ASAP7_75t_SL g1270 ( .A1(n_1248), .A2(n_1271), .B1(n_1272), .B2(n_1275), .C(n_1276), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1249), .B(n_1259), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1250), .B(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1253), .Y(n_1299) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1255), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1261), .Y(n_1259) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
AOI211xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B(n_1279), .C(n_1288), .Y(n_1263) );
INVxp67_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
OAI21xp5_ASAP7_75t_L g1294 ( .A1(n_1275), .A2(n_1295), .B(n_1297), .Y(n_1294) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
OAI21xp5_ASAP7_75t_L g1279 ( .A1(n_1280), .A2(n_1281), .B(n_1282), .Y(n_1279) );
OAI21xp33_ASAP7_75t_L g1323 ( .A1(n_1283), .A2(n_1324), .B(n_1325), .Y(n_1323) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NAND2xp5_ASAP7_75t_SL g1313 ( .A(n_1314), .B(n_1319), .Y(n_1313) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
HB1xp67_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1330), .Y(n_1388) );
AND3x1_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1343), .C(n_1378), .Y(n_1330) );
NOR2xp33_ASAP7_75t_SL g1343 ( .A(n_1344), .B(n_1364), .Y(n_1343) );
OAI22xp33_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1347), .B1(n_1350), .B2(n_1351), .Y(n_1345) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVxp67_ASAP7_75t_SL g1348 ( .A(n_1349), .Y(n_1348) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_1350), .A2(n_1363), .B1(n_1367), .B2(n_1370), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_1354), .A2(n_1359), .B1(n_1374), .B2(n_1376), .Y(n_1373) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx5_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx2_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVxp67_ASAP7_75t_SL g1386 ( .A(n_1387), .Y(n_1386) );
HB1xp67_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
OAI21xp5_ASAP7_75t_L g1391 ( .A1(n_1392), .A2(n_1393), .B(n_1394), .Y(n_1391) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
endmodule