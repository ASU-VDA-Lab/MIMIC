module real_jpeg_23198_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_49;
wire n_52;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_27;
wire n_48;
wire n_19;
wire n_20;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_0),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_7),
.B(n_16),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_9),
.C(n_22),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_6),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_16),
.B(n_22),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_7),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_15),
.B1(n_25),
.B2(n_26),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_10),
.A2(n_21),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

OAI31xp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_30),
.A3(n_33),
.B(n_37),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_27),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_25),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_21),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_47),
.C(n_51),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

AOI31xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.A3(n_44),
.B(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);


endmodule