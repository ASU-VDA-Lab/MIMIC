module fake_jpeg_26592_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_23),
.B1(n_31),
.B2(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_43),
.A2(n_44),
.B1(n_51),
.B2(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_52),
.B1(n_55),
.B2(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_30),
.B1(n_23),
.B2(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_18),
.B1(n_17),
.B2(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_0),
.Y(n_90)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_76),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_68),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_72),
.B1(n_27),
.B2(n_1),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_16),
.B1(n_20),
.B2(n_33),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_41),
.A3(n_38),
.B1(n_33),
.B2(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_78),
.B1(n_46),
.B2(n_66),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_38),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_89),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_38),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_45),
.B1(n_66),
.B2(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_56),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_87),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_59),
.C(n_58),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_100),
.B1(n_107),
.B2(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_99),
.B(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_65),
.B1(n_64),
.B2(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_106),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_0),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_80),
.B1(n_79),
.B2(n_74),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_9),
.C(n_14),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_9),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_84),
.B1(n_83),
.B2(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_129),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_82),
.B1(n_73),
.B2(n_68),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_77),
.B1(n_75),
.B2(n_81),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_101),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_130),
.B(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_125),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_108),
.B1(n_93),
.B2(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_88),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_103),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_79),
.B1(n_69),
.B2(n_87),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_110),
.B1(n_106),
.B2(n_94),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_4),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_126),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_153),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_99),
.B(n_108),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_145),
.B(n_142),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_103),
.B(n_94),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_126),
.A3(n_129),
.B1(n_118),
.B2(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_158),
.B1(n_131),
.B2(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_161),
.B1(n_10),
.B2(n_11),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_111),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_93),
.B1(n_95),
.B2(n_114),
.Y(n_158)
);

AOI22x1_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_114),
.B1(n_105),
.B2(n_6),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_11),
.B(n_13),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_105),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_119),
.Y(n_172)
);

OAI22x1_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_5),
.C(n_7),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_134),
.C(n_141),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_10),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_167),
.B(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_176),
.B(n_182),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_178),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_157),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_137),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_161),
.B1(n_168),
.B2(n_169),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_191),
.B1(n_169),
.B2(n_144),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_155),
.A2(n_133),
.B1(n_137),
.B2(n_12),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_156),
.B1(n_152),
.B2(n_148),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_11),
.B(n_12),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_195),
.B(n_163),
.C(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_204),
.B1(n_190),
.B2(n_175),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_219),
.B(n_195),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_160),
.C(n_143),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_203),
.C(n_209),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_153),
.C(n_145),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_150),
.C(n_162),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

FAx1_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_146),
.CI(n_151),
.CON(n_211),
.SN(n_211)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_174),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_216),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_148),
.C(n_14),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_194),
.C(n_191),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_13),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_177),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_230),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_189),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_206),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_179),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_187),
.C(n_197),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_236),
.C(n_208),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_180),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_193),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_180),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_219),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_199),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_192),
.C(n_185),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_192),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_208),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_250),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_239),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_220),
.B1(n_204),
.B2(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_252),
.B(n_219),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_212),
.Y(n_250)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_228),
.C(n_229),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_227),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_221),
.B1(n_233),
.B2(n_200),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_223),
.B(n_200),
.Y(n_260)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_222),
.C(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_264),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_186),
.B1(n_211),
.B2(n_225),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_273),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_241),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_266),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_268),
.B(n_271),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_277),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_265),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_262),
.C(n_261),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_275),
.B1(n_254),
.B2(n_222),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.C(n_259),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_258),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_289),
.B(n_286),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_282),
.B(n_290),
.Y(n_292)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_276),
.B1(n_243),
.B2(n_211),
.C(n_206),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_199),
.B(n_15),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_199),
.B(n_15),
.Y(n_295)
);


endmodule