module real_jpeg_26042_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_24),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_70),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_62),
.B1(n_64),
.B2(n_70),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_204)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_5),
.A2(n_15),
.B(n_304),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_5),
.B(n_305),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_21),
.B1(n_25),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_41),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_41),
.B1(n_62),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_8),
.A2(n_41),
.B1(n_83),
.B2(n_84),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_20),
.B1(n_31),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_20),
.B1(n_62),
.B2(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_20),
.B1(n_83),
.B2(n_84),
.Y(n_99)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_11),
.B1(n_25),
.B2(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_11),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_52),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_11),
.A2(n_52),
.B1(n_83),
.B2(n_84),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_11),
.B(n_30),
.C(n_33),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_11),
.B(n_29),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_11),
.B(n_59),
.C(n_62),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_11),
.B(n_80),
.C(n_83),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_11),
.B(n_13),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_11),
.B(n_113),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_11),
.B(n_73),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_13),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_13),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_44),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_42),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_27),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_19),
.A2(n_29),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_24),
.B1(n_30),
.B2(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_26),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_28),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_29),
.A2(n_35),
.B1(n_51),
.B2(n_67),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_33),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_38),
.B(n_46),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_49),
.B(n_50),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_86),
.B(n_303),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_47),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_47),
.B(n_301),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.CI(n_65),
.CON(n_47),
.SN(n_47)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_49),
.A2(n_50),
.B(n_68),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_56),
.A2(n_61),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_73),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_57),
.B(n_118),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_61),
.A2(n_117),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_64),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_62),
.B(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.C(n_74),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_66),
.B(n_136),
.C(n_144),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_66),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_66),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_66),
.A2(n_144),
.B1(n_145),
.B2(n_158),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_66),
.A2(n_115),
.B1(n_158),
.B2(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_66),
.B(n_115),
.C(n_197),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_71),
.A2(n_74),
.B1(n_125),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_71),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_74),
.A2(n_125),
.B1(n_126),
.B2(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_74),
.B(n_121),
.C(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_85),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_76),
.B(n_104),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_104),
.B1(n_113),
.B2(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_82),
.A2(n_103),
.B(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_83),
.B(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_300),
.B(n_302),
.Y(n_86)
);

OAI211xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_146),
.B(n_160),
.C(n_299),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_130),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_130),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_108),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_110),
.C(n_119),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_105),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_91),
.A2(n_105),
.B1(n_106),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_91),
.A2(n_101),
.B1(n_133),
.B2(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_93),
.B(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_99),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_94),
.Y(n_203)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_101),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_119),
.B2(n_120),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_111),
.B(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_115),
.B(n_217),
.C(n_219),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_115),
.A2(n_207),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_122),
.B1(n_154),
.B2(n_159),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_121),
.B(n_144),
.C(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_121),
.A2(n_122),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_121),
.A2(n_122),
.B1(n_179),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_170),
.C(n_179),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_122),
.B(n_150),
.C(n_154),
.Y(n_301)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_135),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_134),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_137),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_141),
.A2(n_142),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_141),
.A2(n_142),
.B1(n_230),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_142),
.B(n_224),
.C(n_230),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_142),
.B(n_202),
.C(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_144),
.A2(n_145),
.B1(n_193),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_144),
.A2(n_145),
.B1(n_177),
.B2(n_190),
.Y(n_267)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_145),
.B(n_177),
.C(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_161),
.C(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_148),
.B(n_149),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_183),
.B(n_298),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_181),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_164),
.B(n_181),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_165),
.B(n_167),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_169),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_170),
.A2(n_171),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_177),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_204),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_177),
.A2(n_190),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_177),
.B(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_179),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_293),
.B(n_297),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_220),
.B(n_279),
.C(n_292),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_209),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_186),
.B(n_209),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_196),
.B2(n_208),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_189),
.B(n_195),
.C(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_206),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_201),
.A2(n_202),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_253),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.C(n_216),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_211),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_216),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_278),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_239),
.B(n_277),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_223),
.B(n_236),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_225),
.B1(n_273),
.B2(n_275),
.Y(n_272)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_229),
.B(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_270),
.B(n_276),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_264),
.B(n_269),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_256),
.B(n_263),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_248),
.B(n_255),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_252),
.B(n_254),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_258),
.Y(n_263)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_291),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_289),
.C(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);


endmodule