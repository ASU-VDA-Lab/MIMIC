module fake_jpeg_5889_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_6),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_17),
.B1(n_32),
.B2(n_21),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_56),
.B1(n_33),
.B2(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_17),
.B1(n_32),
.B2(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_32),
.B1(n_17),
.B2(n_45),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_64),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_17),
.B1(n_32),
.B2(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_18),
.B1(n_29),
.B2(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_69),
.B(n_81),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_72),
.A2(n_52),
.B1(n_97),
.B2(n_94),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_77),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_23),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_83),
.C(n_96),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_39),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_28),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_30),
.B1(n_35),
.B2(n_26),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_28),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_28),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_42),
.B1(n_35),
.B2(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_54),
.B1(n_31),
.B2(n_29),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_27),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_27),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_48),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_19),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_50),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_51),
.B1(n_52),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_111),
.B1(n_117),
.B2(n_123),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_56),
.C(n_39),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_106),
.C(n_127),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_39),
.C(n_55),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_51),
.B1(n_52),
.B2(n_36),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_51),
.B1(n_52),
.B2(n_37),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_130),
.B1(n_78),
.B2(n_82),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_54),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_40),
.B1(n_37),
.B2(n_31),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_75),
.C(n_100),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_70),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_136),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_138),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_140),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_148),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_144),
.Y(n_195)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_72),
.B1(n_87),
.B2(n_76),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_153),
.B1(n_161),
.B2(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_155),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_72),
.B(n_83),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_80),
.B(n_83),
.C(n_84),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_85),
.C(n_80),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_156),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_106),
.B(n_124),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_154),
.B(n_31),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_82),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_109),
.B(n_78),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_115),
.B(n_88),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_39),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_162),
.B(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_121),
.B1(n_126),
.B2(n_109),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_178),
.B1(n_180),
.B2(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_181),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_104),
.B1(n_115),
.B2(n_93),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_171),
.B1(n_183),
.B2(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_150),
.B1(n_156),
.B2(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_174),
.B(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_182),
.C(n_20),
.Y(n_197)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_131),
.B1(n_146),
.B2(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_104),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_93),
.B1(n_112),
.B2(n_110),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_122),
.B1(n_107),
.B2(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_107),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_122),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_113),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_129),
.B1(n_98),
.B2(n_95),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_20),
.CI(n_19),
.CON(n_206),
.SN(n_206)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_201),
.C(n_208),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_90),
.B1(n_40),
.B2(n_34),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_215),
.B1(n_175),
.B2(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_209),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_172),
.C(n_182),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_19),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_164),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_222),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_68),
.B1(n_34),
.B2(n_24),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_175),
.B1(n_194),
.B2(n_192),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_20),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_213),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_20),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_218),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_34),
.B1(n_24),
.B2(n_19),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_19),
.C(n_20),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_225),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_19),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_219),
.C(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_68),
.C(n_73),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_162),
.B(n_163),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_34),
.C(n_24),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_0),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_170),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_230),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_184),
.B(n_196),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_1),
.B(n_4),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_187),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_244),
.C(n_247),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_249),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_166),
.B(n_183),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_241),
.B1(n_223),
.B2(n_214),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_209),
.B1(n_225),
.B2(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_217),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_193),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_203),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_169),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_181),
.B1(n_24),
.B2(n_3),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_199),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_207),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_219),
.C(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_269),
.C(n_235),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_231),
.A2(n_205),
.B1(n_218),
.B2(n_206),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_267),
.B(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_226),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_264),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_212),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_243),
.B(n_220),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_206),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_246),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_4),
.B(n_5),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_1),
.C(n_4),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_1),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_11),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_247),
.C(n_232),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_282),
.Y(n_302)
);

BUFx12_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_277),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_258),
.B(n_237),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_231),
.Y(n_280)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_287),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_254),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_230),
.Y(n_301)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_257),
.B1(n_261),
.B2(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_256),
.C(n_253),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_293),
.C(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_285),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_254),
.C(n_235),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_267),
.B1(n_260),
.B2(n_264),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_281),
.B1(n_289),
.B2(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_295),
.A2(n_285),
.B1(n_276),
.B2(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_229),
.C(n_269),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_297),
.A2(n_290),
.B(n_293),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_270),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_273),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_303),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_276),
.B(n_236),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_276),
.B(n_273),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_305),
.A2(n_291),
.B(n_302),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_306),
.B(n_314),
.CI(n_5),
.CON(n_324),
.SN(n_324)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_288),
.B1(n_284),
.B2(n_242),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_309),
.B(n_312),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_287),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_11),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_297),
.C(n_302),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_300),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_312),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_323),
.B(n_325),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.C(n_311),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_12),
.B(n_7),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_316),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_7),
.B(n_10),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_326),
.B(n_328),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_311),
.Y(n_329)
);

AO21x2_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_331),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_318),
.B(n_11),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_324),
.B(n_13),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_332),
.A2(n_333),
.B(n_327),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_13),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_12),
.B(n_15),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_15),
.Y(n_339)
);


endmodule