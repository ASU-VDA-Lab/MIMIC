module fake_ibex_1542_n_964 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_964);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_964;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_167;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_506;
wire n_444;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_927;
wire n_684;
wire n_775;
wire n_934;
wire n_784;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_39),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_60),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_54),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_75),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_92),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_1),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_69),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_58),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_82),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_72),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_38),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_5),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_44),
.B(n_32),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_17),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_119),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_41),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_56),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_103),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g212 ( 
.A(n_81),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_32),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_26),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_16),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_107),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_145),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_12),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_33),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_39),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_110),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_57),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g230 ( 
.A(n_115),
.B(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_123),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_114),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_51),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_59),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_33),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_87),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_134),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_146),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_67),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_117),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_106),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_99),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_147),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_138),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_50),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_113),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_61),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_3),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_80),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_101),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_86),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_85),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_91),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_116),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_139),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_52),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g272 ( 
.A(n_131),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_149),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_93),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_27),
.B(n_104),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_122),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_46),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_6),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_148),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_25),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_160),
.B(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_185),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_181),
.B(n_4),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_194),
.B(n_4),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_254),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_161),
.B(n_8),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_216),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_250),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_254),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_202),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_216),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_194),
.B(n_11),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_165),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_216),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_163),
.B(n_13),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_179),
.Y(n_310)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_249),
.B(n_45),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_13),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_167),
.B(n_15),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_182),
.B(n_189),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_168),
.B(n_15),
.Y(n_315)
);

CKINVDCx8_ASAP7_75t_R g316 ( 
.A(n_164),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_169),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_170),
.B(n_16),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_171),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_193),
.B(n_17),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_172),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_222),
.B(n_18),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_174),
.A2(n_66),
.B(n_155),
.Y(n_323)
);

OAI22x1_ASAP7_75t_L g324 ( 
.A1(n_256),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_198),
.B(n_21),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_176),
.A2(n_70),
.B(n_154),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_204),
.B(n_22),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_202),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_209),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_177),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_178),
.B(n_180),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_213),
.B(n_23),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_215),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_223),
.B(n_240),
.Y(n_335)
);

AND2x4_ASAP7_75t_SL g336 ( 
.A(n_165),
.B(n_79),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_164),
.B(n_76),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_183),
.A2(n_88),
.B(n_153),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_186),
.B(n_27),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_271),
.B(n_68),
.Y(n_341)
);

OR2x6_ASAP7_75t_L g342 ( 
.A(n_196),
.B(n_28),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_187),
.B(n_29),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g345 ( 
.A(n_173),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_191),
.B(n_29),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_195),
.B(n_30),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_199),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_201),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_214),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_206),
.B(n_90),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_207),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_208),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_217),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_279),
.B(n_30),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_216),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_218),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_225),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_219),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_212),
.A2(n_272),
.B1(n_197),
.B2(n_211),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_221),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_224),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_226),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

CKINVDCx11_ASAP7_75t_R g366 ( 
.A(n_281),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_245),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_227),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_173),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_283),
.B(n_286),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_175),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_298),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_228),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_229),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_285),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_320),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_287),
.B(n_233),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_235),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

INVx6_ASAP7_75t_L g383 ( 
.A(n_294),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_184),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_314),
.B(n_237),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_354),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_239),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_R g388 ( 
.A(n_297),
.B(n_184),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_284),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_289),
.B(n_241),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_289),
.B(n_243),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_244),
.Y(n_397)
);

INVx4_ASAP7_75t_SL g398 ( 
.A(n_311),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_316),
.B(n_166),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_190),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_342),
.B(n_245),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_246),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_314),
.B(n_248),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_288),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_294),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_296),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_257),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_352),
.B(n_259),
.Y(n_408)
);

BUFx8_ASAP7_75t_SL g409 ( 
.A(n_307),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_297),
.Y(n_410)
);

XNOR2x2_ASAP7_75t_SL g411 ( 
.A(n_293),
.B(n_281),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_352),
.B(n_317),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_327),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_332),
.A2(n_260),
.B1(n_263),
.B2(n_276),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_342),
.B(n_230),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_317),
.B(n_261),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_299),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_319),
.B(n_262),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_290),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_290),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_292),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_342),
.A2(n_316),
.B1(n_361),
.B2(n_327),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_292),
.Y(n_428)
);

AND3x2_ASAP7_75t_L g429 ( 
.A(n_367),
.B(n_252),
.C(n_265),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_319),
.B(n_264),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_321),
.B(n_274),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_300),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_321),
.B(n_274),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_330),
.B(n_274),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_300),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_301),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_366),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_301),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_331),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_305),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_330),
.B(n_274),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_303),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_349),
.B(n_234),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_310),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_349),
.B(n_234),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_350),
.B(n_200),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_331),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_296),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_295),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_333),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_329),
.Y(n_453)
);

AO21x2_ASAP7_75t_L g454 ( 
.A1(n_338),
.A2(n_275),
.B(n_277),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_295),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_341),
.B(n_203),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_306),
.B(n_242),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_331),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_363),
.B(n_280),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_364),
.A2(n_334),
.B1(n_340),
.B2(n_343),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_296),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_306),
.B(n_280),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_356),
.B(n_277),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_SL g465 ( 
.A(n_291),
.B(n_273),
.C(n_270),
.Y(n_465)
);

NAND2x1p5_ASAP7_75t_L g466 ( 
.A(n_322),
.B(n_267),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_304),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_346),
.B(n_282),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_304),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_322),
.B(n_166),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_309),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_336),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_313),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_304),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_311),
.A2(n_273),
.B1(n_270),
.B2(n_258),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_339),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_307),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_356),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_312),
.B(n_255),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_338),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_423),
.B(n_337),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_405),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_383),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_383),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

AO22x1_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_231),
.B1(n_232),
.B2(n_238),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_369),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_439),
.B(n_232),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_439),
.B(n_253),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_383),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_366),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_448),
.B(n_238),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_401),
.B(n_324),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_412),
.A2(n_318),
.B1(n_315),
.B2(n_348),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_448),
.B(n_458),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_458),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_443),
.B(n_451),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_374),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_253),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_455),
.B(n_220),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_318),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_412),
.A2(n_348),
.B1(n_324),
.B2(n_302),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_468),
.B(n_326),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_384),
.B(n_326),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_326),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_427),
.A2(n_328),
.B1(n_323),
.B2(n_365),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_437),
.A2(n_323),
.B1(n_34),
.B2(n_35),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_371),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_463),
.B(n_385),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_480),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_401),
.B(n_365),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_416),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_385),
.B(n_365),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_409),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_466),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_94),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_478),
.B(n_31),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_450),
.B(n_34),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_408),
.A2(n_357),
.B1(n_308),
.B2(n_37),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_386),
.A2(n_357),
.B(n_308),
.C(n_38),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_389),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_409),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_401),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_386),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_417),
.B(n_43),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_387),
.B(n_44),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_L g539 ( 
.A(n_472),
.B(n_47),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_370),
.A2(n_49),
.B1(n_53),
.B2(n_55),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_389),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_471),
.B(n_65),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_473),
.B(n_89),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_403),
.B(n_447),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_476),
.B(n_95),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_393),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_380),
.B(n_373),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_466),
.B(n_127),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_437),
.B(n_130),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_136),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_395),
.A2(n_396),
.B1(n_374),
.B2(n_390),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_428),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_374),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_445),
.B(n_453),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_461),
.B(n_460),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_461),
.B(n_410),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_475),
.B(n_376),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_374),
.B(n_396),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_378),
.B(n_391),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_396),
.A2(n_374),
.B1(n_465),
.B2(n_457),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_388),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_430),
.B(n_420),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_546),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_520),
.B(n_429),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_501),
.B(n_457),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_561),
.A2(n_422),
.B(n_407),
.C(n_402),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_519),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_547),
.B(n_457),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_524),
.B(n_470),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_518),
.Y(n_574)
);

BUFx12f_ASAP7_75t_L g575 ( 
.A(n_524),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_SL g576 ( 
.A(n_565),
.B(n_415),
.C(n_397),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_SL g577 ( 
.A(n_565),
.B(n_407),
.C(n_381),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_533),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_502),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_484),
.B(n_421),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_504),
.Y(n_582)
);

INVx8_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_507),
.B(n_430),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_506),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_R g588 ( 
.A(n_534),
.B(n_470),
.Y(n_588)
);

O2A1O1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_512),
.A2(n_381),
.B(n_397),
.C(n_459),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_488),
.B(n_442),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_537),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_559),
.A2(n_470),
.B1(n_456),
.B2(n_454),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_516),
.B(n_429),
.Y(n_593)
);

BUFx4f_ASAP7_75t_L g594 ( 
.A(n_519),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_544),
.B(n_456),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_494),
.B(n_426),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_552),
.A2(n_440),
.B1(n_446),
.B2(n_444),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_456),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_496),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_496),
.B(n_440),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_517),
.B(n_454),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_564),
.A2(n_558),
.B1(n_496),
.B2(n_537),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_505),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_500),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_537),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_SL g607 ( 
.A(n_535),
.B(n_411),
.C(n_441),
.Y(n_607)
);

BUFx8_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_496),
.A2(n_433),
.B1(n_434),
.B2(n_431),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_527),
.B(n_411),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_500),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_555),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_487),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_562),
.A2(n_398),
.B1(n_474),
.B2(n_467),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_R g615 ( 
.A(n_562),
.B(n_372),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_503),
.B(n_372),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_563),
.A2(n_377),
.B1(n_379),
.B2(n_382),
.Y(n_617)
);

OA22x2_ASAP7_75t_L g618 ( 
.A1(n_499),
.A2(n_377),
.B1(n_379),
.B2(n_382),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_514),
.B(n_379),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_542),
.A2(n_406),
.B(n_449),
.C(n_462),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_497),
.A2(n_462),
.B1(n_469),
.B2(n_508),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_549),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_550),
.Y(n_623)
);

O2A1O1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_536),
.A2(n_538),
.B(n_532),
.C(n_531),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_529),
.B(n_566),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_550),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_553),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_551),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_553),
.B(n_560),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_566),
.A2(n_489),
.B1(n_483),
.B2(n_493),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_SL g634 ( 
.A(n_532),
.B(n_543),
.C(n_545),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_491),
.A2(n_495),
.B(n_492),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_486),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_554),
.B(n_485),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_522),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_491),
.A2(n_498),
.B(n_481),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_526),
.B(n_481),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_571),
.B(n_490),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_567),
.A2(n_594),
.B1(n_586),
.B2(n_619),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_638),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_590),
.B(n_521),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_610),
.B(n_587),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_582),
.B(n_515),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_571),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_602),
.A2(n_540),
.B1(n_522),
.B2(n_528),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_578),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_626),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_580),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_585),
.B(n_528),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_606),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_622),
.B(n_530),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_608),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_603),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_579),
.Y(n_658)
);

AO32x2_ASAP7_75t_L g659 ( 
.A1(n_617),
.A2(n_609),
.A3(n_597),
.B1(n_634),
.B2(n_618),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_635),
.A2(n_625),
.B(n_629),
.C(n_639),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_636),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_571),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_595),
.A2(n_572),
.B(n_616),
.C(n_569),
.Y(n_663)
);

NOR2x1_ASAP7_75t_R g664 ( 
.A(n_575),
.B(n_613),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_577),
.A2(n_576),
.B(n_619),
.C(n_623),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_592),
.A2(n_627),
.B1(n_633),
.B2(n_591),
.Y(n_666)
);

NOR2x1_ASAP7_75t_SL g667 ( 
.A(n_628),
.B(n_631),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_607),
.A2(n_568),
.B(n_593),
.C(n_596),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_605),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_583),
.B(n_588),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_583),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_608),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_600),
.B(n_598),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_637),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_574),
.A2(n_614),
.B(n_630),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_628),
.A2(n_599),
.B1(n_584),
.B2(n_632),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_604),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_618),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_581),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_573),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_581),
.B(n_611),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_615),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_604),
.A2(n_611),
.B1(n_612),
.B2(n_579),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_586),
.B(n_414),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_586),
.B(n_414),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_602),
.A2(n_586),
.B1(n_629),
.B2(n_594),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_601),
.A2(n_427),
.B(n_512),
.C(n_520),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_601),
.A2(n_570),
.B(n_589),
.C(n_624),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_567),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_586),
.B(n_414),
.Y(n_691)
);

BUFx12f_ASAP7_75t_L g692 ( 
.A(n_575),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

BUFx12f_ASAP7_75t_L g694 ( 
.A(n_575),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_601),
.A2(n_427),
.B(n_512),
.C(n_520),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_638),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_619),
.A2(n_427),
.B1(n_602),
.B2(n_601),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_640),
.A2(n_509),
.B(n_510),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_601),
.A2(n_570),
.B(n_589),
.C(n_624),
.Y(n_700)
);

INVx6_ASAP7_75t_SL g701 ( 
.A(n_628),
.Y(n_701)
);

AO21x1_ASAP7_75t_L g702 ( 
.A1(n_621),
.A2(n_602),
.B(n_512),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_567),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_567),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_586),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_586),
.B(n_516),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_583),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_640),
.A2(n_509),
.B(n_510),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_567),
.B(n_367),
.Y(n_709)
);

OA21x2_ASAP7_75t_L g710 ( 
.A1(n_620),
.A2(n_511),
.B(n_510),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_586),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_586),
.B(n_582),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_601),
.A2(n_427),
.B(n_512),
.C(n_520),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_601),
.A2(n_570),
.B(n_589),
.C(n_624),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_601),
.A2(n_509),
.B(n_510),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_610),
.A2(n_427),
.B1(n_401),
.B2(n_470),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_568),
.B(n_520),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_601),
.A2(n_427),
.B(n_512),
.C(n_520),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_586),
.B(n_516),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_586),
.B(n_414),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_586),
.B(n_414),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_634),
.B(n_592),
.C(n_621),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_601),
.A2(n_570),
.B(n_589),
.C(n_624),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_638),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_586),
.B(n_414),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_638),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_567),
.B(n_367),
.Y(n_727)
);

AO31x2_ASAP7_75t_L g728 ( 
.A1(n_621),
.A2(n_601),
.A3(n_512),
.B(n_620),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_414),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_586),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_567),
.B(n_367),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_601),
.A2(n_570),
.B(n_589),
.C(n_624),
.Y(n_732)
);

AO31x2_ASAP7_75t_L g733 ( 
.A1(n_621),
.A2(n_601),
.A3(n_512),
.B(n_620),
.Y(n_733)
);

AO21x1_ASAP7_75t_L g734 ( 
.A1(n_621),
.A2(n_602),
.B(n_512),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_586),
.Y(n_735)
);

CKINVDCx6p67_ASAP7_75t_R g736 ( 
.A(n_575),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_567),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_602),
.A2(n_586),
.B1(n_629),
.B2(n_594),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_602),
.A2(n_586),
.B1(n_629),
.B2(n_594),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_640),
.A2(n_509),
.B(n_510),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_586),
.B(n_582),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_SL g742 ( 
.A1(n_716),
.A2(n_676),
.B(n_698),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_702),
.A2(n_734),
.B(n_722),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_707),
.B(n_656),
.Y(n_744)
);

OA21x2_ASAP7_75t_L g745 ( 
.A1(n_722),
.A2(n_700),
.B(n_689),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_706),
.B(n_719),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_711),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_684),
.B(n_685),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_641),
.Y(n_749)
);

CKINVDCx14_ASAP7_75t_R g750 ( 
.A(n_736),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_730),
.Y(n_751)
);

OA21x2_ASAP7_75t_L g752 ( 
.A1(n_714),
.A2(n_723),
.B(n_732),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_735),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_704),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_715),
.A2(n_708),
.B(n_740),
.Y(n_755)
);

OAI21x1_ASAP7_75t_SL g756 ( 
.A1(n_686),
.A2(n_739),
.B(n_738),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_698),
.A2(n_686),
.B1(n_738),
.B2(n_739),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_649),
.A2(n_660),
.A3(n_663),
.B(n_699),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_646),
.A2(n_674),
.B1(n_701),
.B2(n_712),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_712),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_691),
.B(n_720),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_671),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_704),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_688),
.A2(n_713),
.B(n_696),
.C(n_718),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_690),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_690),
.B(n_741),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_721),
.B(n_725),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_671),
.B(n_692),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_741),
.B(n_729),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_661),
.Y(n_770)
);

OAI211xp5_ASAP7_75t_L g771 ( 
.A1(n_668),
.A2(n_717),
.B(n_665),
.C(n_676),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_678),
.A2(n_642),
.B1(n_653),
.B2(n_645),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_671),
.B(n_695),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_667),
.A2(n_678),
.B1(n_672),
.B2(n_707),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_655),
.B(n_654),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_643),
.B(n_697),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_650),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_709),
.B(n_731),
.Y(n_778)
);

OAI211xp5_ASAP7_75t_L g779 ( 
.A1(n_687),
.A2(n_703),
.B(n_693),
.C(n_727),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_666),
.A2(n_675),
.B(n_647),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_724),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_675),
.A2(n_657),
.B(n_669),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_701),
.A2(n_652),
.B1(n_726),
.B2(n_673),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_737),
.B(n_679),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_644),
.B(n_648),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_662),
.A2(n_682),
.B1(n_681),
.B2(n_670),
.Y(n_786)
);

OA21x2_ASAP7_75t_L g787 ( 
.A1(n_728),
.A2(n_733),
.B(n_659),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_658),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_683),
.A2(n_710),
.B(n_651),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_680),
.B(n_677),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_658),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_694),
.B(n_658),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_659),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_664),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_705),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_709),
.B(n_590),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_671),
.B(n_586),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_698),
.A2(n_738),
.B1(n_739),
.B2(n_686),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_705),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_705),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_706),
.B(n_719),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_690),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_705),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_704),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_705),
.Y(n_805)
);

OAI221xp5_ASAP7_75t_L g806 ( 
.A1(n_716),
.A2(n_607),
.B1(n_427),
.B2(n_520),
.C(n_496),
.Y(n_806)
);

OAI211xp5_ASAP7_75t_SL g807 ( 
.A1(n_716),
.A2(n_607),
.B(n_668),
.C(n_520),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_695),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_706),
.B(n_719),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_706),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_706),
.B(n_719),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_706),
.B(n_719),
.Y(n_812)
);

AOI221xp5_ASAP7_75t_L g813 ( 
.A1(n_688),
.A2(n_427),
.B1(n_520),
.B2(n_713),
.C(n_696),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_686),
.Y(n_814)
);

OA21x2_ASAP7_75t_L g815 ( 
.A1(n_702),
.A2(n_734),
.B(n_722),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_705),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_706),
.B(n_719),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_705),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_742),
.A2(n_807),
.B1(n_806),
.B2(n_813),
.Y(n_819)
);

AOI221x1_ASAP7_75t_SL g820 ( 
.A1(n_777),
.A2(n_818),
.B1(n_800),
.B2(n_803),
.C(n_805),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_752),
.B(n_745),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_SL g822 ( 
.A1(n_757),
.A2(n_798),
.B(n_772),
.Y(n_822)
);

OAI211xp5_ASAP7_75t_L g823 ( 
.A1(n_779),
.A2(n_759),
.B(n_771),
.C(n_807),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_760),
.B(n_745),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_752),
.B(n_766),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_802),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_789),
.B(n_814),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_756),
.A2(n_769),
.B1(n_759),
.B2(n_814),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_764),
.A2(n_780),
.B(n_755),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_SL g830 ( 
.A1(n_762),
.A2(n_797),
.B(n_786),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_810),
.A2(n_809),
.B1(n_811),
.B2(n_812),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_793),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_787),
.B(n_782),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_787),
.B(n_743),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_743),
.B(n_815),
.Y(n_835)
);

INVx3_ASAP7_75t_SL g836 ( 
.A(n_744),
.Y(n_836)
);

OAI211xp5_ASAP7_75t_L g837 ( 
.A1(n_779),
.A2(n_771),
.B(n_774),
.C(n_783),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_802),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_788),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_749),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_770),
.B(n_758),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_SL g842 ( 
.A(n_774),
.B(n_783),
.C(n_765),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_781),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_SL g844 ( 
.A1(n_762),
.A2(n_797),
.B(n_786),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_810),
.A2(n_817),
.B1(n_801),
.B2(n_746),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_781),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_751),
.Y(n_847)
);

OA21x2_ASAP7_75t_L g848 ( 
.A1(n_791),
.A2(n_795),
.B(n_747),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_753),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_799),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_778),
.B(n_796),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_748),
.A2(n_761),
.B(n_767),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_841),
.B(n_816),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_848),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_841),
.B(n_785),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_832),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_841),
.B(n_776),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_827),
.B(n_744),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_824),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_839),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_821),
.B(n_825),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_821),
.B(n_775),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_824),
.B(n_744),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_847),
.B(n_775),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_830),
.B(n_773),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_833),
.B(n_808),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_833),
.B(n_804),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_833),
.B(n_754),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_819),
.A2(n_794),
.B1(n_792),
.B2(n_763),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_840),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_847),
.B(n_790),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_825),
.B(n_792),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_840),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_856),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_861),
.B(n_846),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_861),
.B(n_834),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_861),
.B(n_834),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_861),
.B(n_846),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_854),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_860),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_853),
.B(n_834),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_865),
.B(n_836),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_859),
.B(n_835),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_856),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_857),
.B(n_843),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_858),
.B(n_827),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_860),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_855),
.B(n_825),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_876),
.B(n_867),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_874),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_820),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_887),
.B(n_858),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_876),
.B(n_867),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_884),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_884),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_883),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_888),
.B(n_820),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_883),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_879),
.B(n_837),
.C(n_823),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_887),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_886),
.B(n_858),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_891),
.B(n_876),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_897),
.B(n_877),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_889),
.B(n_877),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_896),
.B(n_877),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_900),
.B(n_879),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_896),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_900),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_899),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_889),
.B(n_881),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_893),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_898),
.B(n_883),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_898),
.B(n_875),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_893),
.B(n_890),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_913),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_907),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_913),
.Y(n_917)
);

OAI21xp33_ASAP7_75t_L g918 ( 
.A1(n_909),
.A2(n_892),
.B(n_901),
.Y(n_918)
);

OAI21xp33_ASAP7_75t_L g919 ( 
.A1(n_902),
.A2(n_892),
.B(n_901),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_903),
.A2(n_837),
.B1(n_823),
.B2(n_901),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_914),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_906),
.A2(n_865),
.B(n_844),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_904),
.B(n_881),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_912),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_908),
.A2(n_882),
.B(n_865),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_904),
.B(n_890),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_911),
.A2(n_873),
.B(n_870),
.Y(n_927)
);

NOR2x1_ASAP7_75t_SL g928 ( 
.A(n_923),
.B(n_910),
.Y(n_928)
);

OAI211xp5_ASAP7_75t_SL g929 ( 
.A1(n_920),
.A2(n_869),
.B(n_750),
.C(n_819),
.Y(n_929)
);

OAI322xp33_ASAP7_75t_L g930 ( 
.A1(n_915),
.A2(n_905),
.A3(n_875),
.B1(n_878),
.B2(n_885),
.C1(n_822),
.C2(n_863),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_919),
.A2(n_858),
.B1(n_910),
.B2(n_872),
.Y(n_931)
);

AOI321xp33_ASAP7_75t_L g932 ( 
.A1(n_918),
.A2(n_869),
.A3(n_872),
.B1(n_828),
.B2(n_866),
.C(n_868),
.Y(n_932)
);

AOI211xp5_ASAP7_75t_L g933 ( 
.A1(n_922),
.A2(n_794),
.B(n_836),
.C(n_768),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_917),
.A2(n_886),
.B(n_878),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_927),
.B(n_880),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_921),
.A2(n_858),
.B1(n_872),
.B2(n_886),
.Y(n_936)
);

OAI221xp5_ASAP7_75t_L g937 ( 
.A1(n_932),
.A2(n_925),
.B1(n_924),
.B2(n_926),
.C(n_916),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_SL g938 ( 
.A1(n_933),
.A2(n_852),
.B(n_916),
.C(n_829),
.Y(n_938)
);

AOI222xp33_ASAP7_75t_L g939 ( 
.A1(n_928),
.A2(n_935),
.B1(n_934),
.B2(n_929),
.C1(n_923),
.C2(n_842),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_931),
.A2(n_936),
.B1(n_858),
.B2(n_872),
.Y(n_940)
);

XNOR2xp5_ASAP7_75t_L g941 ( 
.A(n_930),
.B(n_867),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_SL g942 ( 
.A1(n_928),
.A2(n_866),
.B1(n_868),
.B2(n_862),
.Y(n_942)
);

AOI21xp33_ASAP7_75t_SL g943 ( 
.A1(n_935),
.A2(n_836),
.B(n_792),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_938),
.A2(n_939),
.B(n_943),
.C(n_937),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_942),
.B(n_842),
.C(n_852),
.Y(n_945)
);

NAND4xp25_ASAP7_75t_L g946 ( 
.A(n_940),
.B(n_828),
.C(n_831),
.D(n_845),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_941),
.Y(n_947)
);

NOR3xp33_ASAP7_75t_L g948 ( 
.A(n_938),
.B(n_784),
.C(n_851),
.Y(n_948)
);

OR5x1_ASAP7_75t_L g949 ( 
.A(n_944),
.B(n_836),
.C(n_794),
.D(n_851),
.E(n_863),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_948),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_SL g951 ( 
.A(n_947),
.B(n_829),
.C(n_851),
.Y(n_951)
);

XNOR2x1_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_794),
.Y(n_952)
);

NAND4xp25_ASAP7_75t_L g953 ( 
.A(n_945),
.B(n_845),
.C(n_831),
.D(n_863),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_944),
.B(n_871),
.C(n_864),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_950),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_954),
.B(n_868),
.Y(n_956)
);

NOR4xp25_ASAP7_75t_L g957 ( 
.A(n_951),
.B(n_847),
.C(n_864),
.D(n_850),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_955),
.A2(n_952),
.B1(n_949),
.B2(n_953),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_956),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_957),
.B(n_956),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_959),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_961),
.A2(n_838),
.B1(n_826),
.B2(n_866),
.Y(n_962)
);

AO221x1_ASAP7_75t_L g963 ( 
.A1(n_962),
.A2(n_850),
.B1(n_849),
.B2(n_895),
.C(n_894),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_963),
.A2(n_838),
.B1(n_826),
.B2(n_843),
.Y(n_964)
);


endmodule