module fake_jpeg_4410_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_31),
.B1(n_19),
.B2(n_22),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_66),
.B(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_60),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_69),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_31),
.B1(n_19),
.B2(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_26),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_23),
.B(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_27),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_73),
.A2(n_78),
.B1(n_81),
.B2(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_25),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_31),
.B1(n_19),
.B2(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_31),
.B1(n_19),
.B2(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_91),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_97),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_66),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_67),
.B1(n_61),
.B2(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_118),
.B1(n_28),
.B2(n_17),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_110),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_62),
.B1(n_56),
.B2(n_54),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_50),
.B1(n_48),
.B2(n_52),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_72),
.B1(n_76),
.B2(n_82),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_115),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_56),
.B1(n_54),
.B2(n_59),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_120),
.B1(n_82),
.B2(n_27),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_47),
.B1(n_27),
.B2(n_32),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_42),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_64),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_135),
.B1(n_97),
.B2(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_129),
.A2(n_18),
.B1(n_20),
.B2(n_33),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_29),
.B(n_17),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_16),
.B(n_28),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_137),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_89),
.B1(n_29),
.B2(n_28),
.Y(n_168)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_41),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_116),
.B1(n_111),
.B2(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_169),
.B(n_173),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_105),
.B1(n_118),
.B2(n_95),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_157),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_161),
.C(n_127),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_116),
.B(n_113),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_156),
.B(n_163),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_108),
.B(n_32),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_102),
.C(n_42),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_132),
.B1(n_130),
.B2(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_51),
.B1(n_24),
.B2(n_30),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_138),
.B1(n_136),
.B2(n_142),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_176),
.B1(n_18),
.B2(n_138),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_124),
.A2(n_30),
.A3(n_33),
.B1(n_23),
.B2(n_42),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_122),
.B1(n_141),
.B2(n_135),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_198),
.C(n_93),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_181),
.B(n_183),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_143),
.B(n_127),
.C(n_125),
.D(n_139),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_165),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_140),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_185),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_140),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_195),
.B(n_197),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_162),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_138),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_196),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_176),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_42),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_58),
.C(n_64),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_40),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_202),
.B1(n_151),
.B2(n_157),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_224),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_177),
.A2(n_170),
.B1(n_149),
.B2(n_163),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_225),
.B1(n_223),
.B2(n_208),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_30),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_179),
.B1(n_181),
.B2(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_223),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_175),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_172),
.B1(n_153),
.B2(n_136),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_200),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_198),
.C(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_136),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_212),
.C(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_189),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_221),
.C(n_213),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_189),
.B(n_203),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_240),
.B(n_245),
.Y(n_260)
);

BUFx12_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_246),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_203),
.B(n_199),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_205),
.B(n_186),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_199),
.B(n_142),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_206),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_142),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_238),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_261),
.B(n_235),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_255),
.C(n_262),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_211),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_267),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_221),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_265),
.B(n_266),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_233),
.C(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_12),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_237),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_93),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

NOR4xp25_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_243),
.C(n_247),
.D(n_230),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_271),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_279),
.C(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_3),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_280),
.B1(n_268),
.B2(n_33),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_242),
.B1(n_240),
.B2(n_234),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_267),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_258),
.A2(n_244),
.B1(n_234),
.B2(n_249),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_239),
.B(n_114),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_13),
.C(n_15),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_255),
.C(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_290),
.C(n_292),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_254),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_294),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_103),
.B1(n_93),
.B2(n_90),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_289),
.B1(n_294),
.B2(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_90),
.C(n_84),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_90),
.B1(n_33),
.B2(n_30),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_273),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_1),
.C(n_2),
.Y(n_294)
);

NOR2x1_ASAP7_75t_SL g298 ( 
.A(n_296),
.B(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_300),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_5),
.C(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_275),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_305),
.B1(n_7),
.B2(n_8),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_269),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_5),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_6),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_282),
.B1(n_6),
.B2(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_311),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_313),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_299),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_10),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_302),
.C(n_307),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_320),
.A3(n_316),
.B1(n_306),
.B2(n_318),
.C1(n_305),
.C2(n_314),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_310),
.B(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_10),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_10),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_11),
.C(n_13),
.Y(n_325)
);

OAI221xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_143),
.Y(n_326)
);


endmodule