module fake_jpeg_4063_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_34),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_54),
.B(n_20),
.C(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_18),
.B1(n_19),
.B2(n_16),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_24),
.B(n_20),
.C(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_16),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_16),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_72),
.B1(n_19),
.B2(n_16),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_67),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_75),
.Y(n_100)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_87),
.B1(n_74),
.B2(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_20),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_44),
.B1(n_49),
.B2(n_42),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_64),
.C(n_61),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_42),
.B1(n_63),
.B2(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_77),
.B1(n_67),
.B2(n_70),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_92),
.C(n_114),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_15),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_58),
.B1(n_59),
.B2(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_58),
.B1(n_51),
.B2(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

AOI22x1_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_63),
.B1(n_39),
.B2(n_40),
.Y(n_102)
);

NAND5xp2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_68),
.C(n_51),
.D(n_55),
.E(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_63),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_63),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_114),
.B(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_26),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_83),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_123),
.B(n_108),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_23),
.B(n_27),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_126),
.B(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_78),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_90),
.B1(n_111),
.B2(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_120),
.B(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_76),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_68),
.C(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

OAI31xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_48),
.A3(n_55),
.B(n_27),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_102),
.B(n_109),
.C(n_110),
.D(n_95),
.Y(n_142)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_69),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_30),
.B(n_19),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_97),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_51),
.C(n_62),
.Y(n_141)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_136),
.Y(n_183)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_148),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_155),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_89),
.B1(n_100),
.B2(n_93),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_139),
.B1(n_115),
.B2(n_121),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_105),
.B1(n_99),
.B2(n_108),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_162),
.B1(n_163),
.B2(n_167),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_30),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_128),
.B(n_117),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_134),
.B(n_141),
.Y(n_175)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_105),
.B1(n_103),
.B2(n_30),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_55),
.B1(n_17),
.B2(n_82),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_145),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_171),
.C(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_116),
.C(n_122),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_190),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_129),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_191),
.B(n_165),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_167),
.B(n_148),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_119),
.B1(n_115),
.B2(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_153),
.A2(n_142),
.B1(n_164),
.B2(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_116),
.B1(n_123),
.B2(n_140),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_137),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_136),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_136),
.B1(n_118),
.B2(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_159),
.B1(n_158),
.B2(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_189),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_17),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_26),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_26),
.B(n_23),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_163),
.B1(n_143),
.B2(n_162),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_167),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_143),
.C(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_196),
.B(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_166),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_204),
.B(n_184),
.Y(n_223)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_219),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_217),
.Y(n_234)
);

XOR2x2_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_148),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_187),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_26),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_147),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_183),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_175),
.C(n_182),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_226),
.C(n_229),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_206),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_181),
.B1(n_185),
.B2(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_233),
.B1(n_238),
.B2(n_205),
.Y(n_244)
);

NOR3xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_197),
.C(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_180),
.C(n_179),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_172),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_212),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_177),
.B1(n_186),
.B2(n_192),
.Y(n_233)
);

XOR2x2_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_191),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_198),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_190),
.C(n_188),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_237),
.C(n_240),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_148),
.B1(n_147),
.B2(n_97),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_106),
.C(n_26),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_256),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_255),
.B(n_28),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_257),
.B1(n_13),
.B2(n_11),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_198),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_212),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_254),
.B1(n_10),
.B2(n_11),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_211),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_230),
.A2(n_211),
.B1(n_201),
.B2(n_214),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_236),
.B1(n_228),
.B2(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_201),
.C(n_106),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_106),
.C(n_28),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_240),
.B1(n_227),
.B2(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

OAI321xp33_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_229),
.A3(n_224),
.B1(n_28),
.B2(n_27),
.C(n_23),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_241),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_259),
.B1(n_252),
.B2(n_255),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_270),
.B1(n_10),
.B2(n_1),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_245),
.C(n_28),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_269),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_23),
.B(n_27),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_267),
.B1(n_28),
.B2(n_27),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_26),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_241),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_265),
.A3(n_269),
.B1(n_272),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_278),
.C(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_273),
.B(n_245),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_26),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_266),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_2),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_274),
.B(n_13),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_288),
.C(n_0),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_82),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_286),
.B(n_3),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_0),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_264),
.C(n_275),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_293),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_292),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_280),
.A3(n_282),
.B1(n_281),
.B2(n_288),
.C1(n_277),
.C2(n_287),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_0),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_298),
.Y(n_300)
);

OAI221xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_4),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_1),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_4),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_5),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_9),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_5),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_296),
.B(n_293),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_307),
.A2(n_297),
.B(n_7),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_309),
.B(n_310),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_289),
.C(n_8),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_314),
.B1(n_312),
.B2(n_307),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_6),
.Y(n_317)
);


endmodule