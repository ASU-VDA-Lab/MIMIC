module fake_jpeg_29776_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_38),
.B(n_15),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_43),
.C(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_69),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_46),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_54),
.B1(n_50),
.B2(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_52),
.B1(n_17),
.B2(n_18),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_82),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_50),
.B1(n_41),
.B2(n_52),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_36),
.B1(n_11),
.B2(n_12),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_14),
.B1(n_20),
.B2(n_21),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_86),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_46),
.C(n_16),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_9),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_5),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_5),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_8),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_6),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_29),
.C(n_30),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_10),
.B(n_13),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_23),
.C(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_107),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_27),
.B(n_28),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_109),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_115),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_92),
.C(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_114),
.C(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_93),
.B1(n_95),
.B2(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_112),
.B1(n_104),
.B2(n_102),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_116),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_113),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_31),
.B(n_32),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_33),
.Y(n_123)
);


endmodule