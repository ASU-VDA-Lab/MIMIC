module real_jpeg_11128_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_1),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_6),
.B(n_65),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_56),
.B1(n_60),
.B2(n_68),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_6),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_71),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_38),
.B(n_42),
.C(n_127),
.D(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_6),
.B(n_38),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_6),
.B(n_80),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_24),
.B(n_142),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_64),
.B(n_76),
.C(n_94),
.D(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_6),
.B(n_64),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g78 ( 
.A(n_9),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_13),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_60),
.B1(n_68),
.B2(n_82),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_82),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_82),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_14),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_85),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_85),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_104),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_24),
.A2(n_31),
.B1(n_33),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_24),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_25),
.A2(n_30),
.B1(n_103),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_25),
.A2(n_30),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_25),
.B(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_26),
.B(n_43),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_26),
.B(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_27),
.A2(n_45),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_30),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_33),
.A2(n_148),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_33),
.B(n_67),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_33),
.A2(n_156),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_49),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_38),
.A2(n_39),
.B1(n_77),
.B2(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_38),
.B(n_77),
.Y(n_178)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_39),
.A2(n_79),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_41),
.A2(n_49),
.B1(n_139),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_41),
.A2(n_170),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_55),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_49),
.A2(n_53),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_49),
.B(n_67),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.C(n_73),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_51),
.A2(n_52),
.B1(n_73),
.B2(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_66),
.B(n_69),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_61),
.B(n_67),
.C(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_77),
.B(n_79),
.C(n_80),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_77),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_84),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_83),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_96),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_101),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_109),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_105),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_116),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_111),
.A2(n_112),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_115),
.B(n_116),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_117),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_196),
.B(n_201),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_183),
.B(n_195),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_164),
.B(n_182),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_144),
.B(n_163),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_125),
.B(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_127),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_141),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_152),
.B(n_162),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_150),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_157),
.B(n_161),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_166),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_175),
.B2(n_181),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_174),
.C(n_181),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_179),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_185),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_191),
.C(n_193),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_190),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);


endmodule