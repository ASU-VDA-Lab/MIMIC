module fake_jpeg_26955_n_254 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_36),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_26),
.B1(n_31),
.B2(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_64),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_18),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_20),
.B1(n_30),
.B2(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_85),
.B1(n_38),
.B2(n_44),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_69),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_51),
.B1(n_47),
.B2(n_21),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_77),
.B1(n_82),
.B2(n_89),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_75),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_35),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_79),
.B(n_92),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_18),
.B1(n_30),
.B2(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_36),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_86),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_38),
.B1(n_44),
.B2(n_34),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_40),
.B(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_25),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_36),
.C(n_43),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_36),
.C(n_43),
.Y(n_104)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_68),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_43),
.B1(n_59),
.B2(n_40),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_121),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_115),
.C(n_1),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_28),
.B1(n_17),
.B2(n_25),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_28),
.B1(n_17),
.B2(n_32),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_29),
.A3(n_32),
.B1(n_19),
.B2(n_24),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_32),
.A3(n_29),
.B1(n_73),
.B2(n_90),
.C(n_24),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_36),
.C(n_32),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_29),
.B(n_19),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_97),
.B(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_28),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_88),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_32),
.B1(n_19),
.B2(n_36),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_86),
.B1(n_70),
.B2(n_66),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_145),
.B1(n_146),
.B2(n_131),
.Y(n_162)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_70),
.B1(n_76),
.B2(n_82),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_133),
.B1(n_117),
.B2(n_123),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_84),
.B1(n_81),
.B2(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_124),
.B1(n_101),
.B2(n_109),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_134),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_93),
.B1(n_91),
.B2(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_91),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_147),
.B(n_115),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_124),
.B1(n_109),
.B2(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_29),
.B1(n_24),
.B2(n_2),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_29),
.B1(n_24),
.B2(n_2),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_118),
.B(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_105),
.B(n_0),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_2),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_167),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_104),
.C(n_121),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_164),
.C(n_170),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_130),
.A3(n_148),
.B1(n_134),
.B2(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_126),
.B1(n_141),
.B2(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_101),
.C(n_114),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_145),
.B1(n_125),
.B2(n_129),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_126),
.B1(n_138),
.B2(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_168),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_3),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_6),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_3),
.C(n_4),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_3),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_186),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_185),
.B1(n_163),
.B2(n_12),
.Y(n_206)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_209)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_190)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_8),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_167),
.B(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_9),
.B(n_10),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_153),
.C(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_207),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_191),
.B(n_188),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_165),
.B1(n_172),
.B2(n_157),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_192),
.B1(n_181),
.B2(n_189),
.Y(n_220)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_171),
.A3(n_169),
.B1(n_156),
.B2(n_154),
.C1(n_170),
.C2(n_152),
.Y(n_203)
);

OA21x2_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_191),
.B(n_193),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_164),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_208),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_211),
.B1(n_179),
.B2(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_11),
.C(n_12),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_13),
.C(n_14),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_13),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_208),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_223),
.Y(n_224)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_218),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_180),
.B(n_188),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_183),
.B(n_205),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_209),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_220),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_206),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_219),
.B(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_233),
.Y(n_240)
);

OAI221xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_222),
.B1(n_207),
.B2(n_213),
.C(n_221),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_225),
.B(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_227),
.B1(n_224),
.B2(n_231),
.Y(n_242)
);

AOI31xp33_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_217),
.A3(n_221),
.B(n_213),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_198),
.C(n_177),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_245),
.B(n_196),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_238),
.B1(n_237),
.B2(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_249),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_196),
.B(n_15),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_250),
.B(n_246),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_16),
.Y(n_254)
);


endmodule