module fake_jpeg_3552_n_127 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_42),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_32),
.B1(n_41),
.B2(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_34),
.C(n_35),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_41),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_51),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_71),
.C(n_68),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_43),
.C(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_58),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_3),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_40),
.B1(n_5),
.B2(n_6),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_4),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_40),
.C(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_5),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_14),
.C(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_6),
.B(n_7),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_20),
.B(n_30),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_13),
.B(n_29),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_106),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_107)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_8),
.C(n_9),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_99),
.C(n_101),
.Y(n_117)
);

OAI322xp33_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_100),
.A3(n_8),
.B1(n_10),
.B2(n_12),
.C1(n_22),
.C2(n_24),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_120),
.B(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_115),
.B1(n_114),
.B2(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_11),
.Y(n_122)
);

OAI321xp33_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_115),
.A3(n_98),
.B1(n_116),
.B2(n_109),
.C(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_117),
.Y(n_127)
);


endmodule