module fake_jpeg_28132_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_16),
.B1(n_17),
.B2(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_20),
.B1(n_17),
.B2(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_16),
.B1(n_23),
.B2(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_38),
.B1(n_10),
.B2(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_20),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_23),
.B(n_2),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_10),
.B(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_34),
.B1(n_11),
.B2(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_35),
.B(n_38),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_32),
.C(n_21),
.Y(n_52)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_5),
.B(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_34),
.B1(n_18),
.B2(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_42),
.B1(n_2),
.B2(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_48),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_32),
.C(n_14),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_56),
.C(n_46),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_32),
.C(n_4),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.C(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_4),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_55),
.C(n_50),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_61),
.C(n_7),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_64),
.C(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_7),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);


endmodule