module fake_jpeg_16884_n_61 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_59;
wire n_20;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_24;
wire n_26;
wire n_36;
wire n_56;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_4),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.C(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_5),
.B1(n_16),
.B2(n_22),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_38),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_51),
.B2(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_39),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_25),
.B(n_37),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_19),
.B(n_20),
.C(n_31),
.D(n_32),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_34),
.B(n_35),
.C(n_26),
.Y(n_61)
);


endmodule