module fake_netlist_6_4862_n_837 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_837);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_837;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_817;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_45),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_12),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_36),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_82),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_85),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_27),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_10),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_77),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_22),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_23),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_10),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_98),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_34),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_19),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_90),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_88),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_105),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_153),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_75),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_144),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_132),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_24),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_128),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_53),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_100),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_41),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_121),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_26),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_7),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_101),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_44),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_67),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_69),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_143),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_109),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_83),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_107),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_12),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_17),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_174),
.B(n_220),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_180),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

CKINVDCx6p67_ASAP7_75t_R g247 ( 
.A(n_170),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_176),
.A2(n_240),
.B1(n_229),
.B2(n_199),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_201),
.Y(n_250)
);

CKINVDCx11_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g254 ( 
.A(n_171),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_169),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_174),
.B(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_172),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_171),
.Y(n_264)
);

BUFx8_ASAP7_75t_SL g265 ( 
.A(n_214),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_179),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

BUFx8_ASAP7_75t_SL g269 ( 
.A(n_219),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_181),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_228),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_177),
.B(n_1),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_177),
.B(n_1),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_185),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_182),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_196),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_196),
.B(n_18),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_183),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_187),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_2),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_192),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_232),
.B(n_3),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_195),
.A2(n_86),
.B(n_165),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_225),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_256),
.B(n_207),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_SL g302 ( 
.A(n_243),
.B(n_226),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_184),
.Y(n_307)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_256),
.B(n_186),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_276),
.B(n_243),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_276),
.B(n_189),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_270),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_193),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_245),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_265),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_259),
.B(n_203),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_260),
.A2(n_262),
.B1(n_248),
.B2(n_258),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_255),
.B(n_194),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g330 ( 
.A(n_260),
.B(n_204),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_253),
.B(n_197),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_272),
.B(n_205),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_257),
.B(n_198),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_245),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_267),
.B(n_263),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_321),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_282),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_285),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_282),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_294),
.B(n_248),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_271),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_254),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_330),
.B(n_268),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_317),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_254),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_SL g363 ( 
.A(n_297),
.B(n_275),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_317),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_247),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_261),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_279),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_302),
.A2(n_231),
.B1(n_244),
.B2(n_292),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_295),
.A2(n_329),
.B(n_327),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_302),
.A2(n_324),
.B1(n_307),
.B2(n_309),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_344),
.B(n_274),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_311),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_320),
.B(n_274),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_320),
.B(n_290),
.Y(n_381)
);

NAND3xp33_ASAP7_75t_L g382 ( 
.A(n_307),
.B(n_287),
.C(n_275),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_292),
.C(n_287),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_297),
.B(n_290),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_286),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_337),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_300),
.B(n_202),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_312),
.B(n_288),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_312),
.B(n_251),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_312),
.B(n_291),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_300),
.B(n_208),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_339),
.B(n_209),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_339),
.B(n_210),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_339),
.B(n_212),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_251),
.Y(n_401)
);

AO221x1_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_236),
.B1(n_215),
.B2(n_218),
.C(n_223),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_L g403 ( 
.A(n_303),
.B(n_283),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_303),
.B(n_213),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_304),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_304),
.B(n_216),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_305),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_305),
.B(n_250),
.Y(n_408)
);

AO32x1_ASAP7_75t_L g409 ( 
.A1(n_405),
.A2(n_344),
.A3(n_343),
.B1(n_338),
.B2(n_335),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_360),
.B(n_217),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_357),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_246),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_378),
.A2(n_343),
.B(n_338),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_378),
.A2(n_335),
.B(n_333),
.Y(n_415)
);

O2A1O1Ixp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_363),
.B(n_382),
.C(n_353),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_358),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_369),
.A2(n_333),
.B(n_328),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_211),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_382),
.A2(n_383),
.B(n_371),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_398),
.A2(n_328),
.B(n_325),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_399),
.A2(n_325),
.B(n_318),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_351),
.B(n_313),
.Y(n_427)
);

BUFx8_ASAP7_75t_SL g428 ( 
.A(n_362),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_400),
.A2(n_318),
.B(n_316),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_345),
.B(n_313),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_367),
.A2(n_293),
.B(n_224),
.C(n_230),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_349),
.B(n_314),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_364),
.Y(n_433)
);

AO21x1_ASAP7_75t_L g434 ( 
.A1(n_403),
.A2(n_233),
.B(n_238),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_379),
.A2(n_222),
.B1(n_234),
.B2(n_237),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_368),
.B(n_314),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_373),
.A2(n_242),
.B1(n_283),
.B2(n_315),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_392),
.A2(n_249),
.B(n_315),
.C(n_316),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_374),
.B(n_388),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_380),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_359),
.A2(n_283),
.B1(n_250),
.B2(n_269),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_348),
.A2(n_393),
.B(n_387),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_283),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_20),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_375),
.B(n_3),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_355),
.B(n_21),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_25),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_396),
.A2(n_91),
.B(n_164),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_346),
.A2(n_87),
.B1(n_163),
.B2(n_162),
.Y(n_453)
);

AND3x1_ASAP7_75t_SL g454 ( 
.A(n_402),
.B(n_4),
.C(n_5),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_397),
.A2(n_81),
.B(n_161),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_385),
.B(n_29),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_408),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_394),
.B(n_4),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_366),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_6),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_30),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_390),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_404),
.A2(n_93),
.B(n_159),
.Y(n_465)
);

BUFx4f_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_31),
.Y(n_467)
);

NAND2x1p5_ASAP7_75t_L g468 ( 
.A(n_350),
.B(n_33),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_352),
.B(n_8),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_376),
.B(n_8),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_382),
.A2(n_9),
.B(n_11),
.C(n_13),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_378),
.A2(n_94),
.B(n_158),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_354),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_347),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_351),
.B(n_9),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_351),
.B(n_38),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_452),
.A2(n_459),
.B(n_432),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_420),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_412),
.B(n_11),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_419),
.B(n_473),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_166),
.B(n_97),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_411),
.B(n_39),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_424),
.A2(n_99),
.B(n_156),
.Y(n_485)
);

AND2x6_ASAP7_75t_SL g486 ( 
.A(n_462),
.B(n_13),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_14),
.Y(n_487)
);

AO31x2_ASAP7_75t_L g488 ( 
.A1(n_431),
.A2(n_15),
.A3(n_16),
.B(n_40),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

OAI22x1_ASAP7_75t_L g490 ( 
.A1(n_448),
.A2(n_15),
.B1(n_16),
.B2(n_42),
.Y(n_490)
);

NOR2x1_ASAP7_75t_SL g491 ( 
.A(n_476),
.B(n_43),
.Y(n_491)
);

BUFx8_ASAP7_75t_SL g492 ( 
.A(n_428),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_442),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_416),
.A2(n_46),
.B(n_47),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_427),
.B(n_48),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_433),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_430),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_418),
.A2(n_49),
.B(n_50),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_457),
.B(n_51),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_464),
.A2(n_52),
.B(n_54),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_443),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_56),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_421),
.B(n_57),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_466),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_458),
.B(n_62),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_420),
.B(n_63),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_421),
.B(n_65),
.Y(n_511)
);

AO32x2_ASAP7_75t_L g512 ( 
.A1(n_453),
.A2(n_68),
.A3(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_439),
.B(n_78),
.Y(n_513)
);

AO31x2_ASAP7_75t_L g514 ( 
.A1(n_434),
.A2(n_79),
.A3(n_80),
.B(n_84),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_425),
.A2(n_92),
.B(n_102),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_417),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_111),
.Y(n_517)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_456),
.A2(n_112),
.B(n_113),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_429),
.A2(n_116),
.B(n_117),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_422),
.B(n_120),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_122),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_461),
.B(n_470),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_435),
.B(n_123),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_414),
.A2(n_415),
.B(n_467),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_463),
.A2(n_124),
.B(n_125),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_437),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_410),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_446),
.A2(n_129),
.B(n_133),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_471),
.B(n_134),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_449),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_444),
.B(n_139),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_525),
.A2(n_450),
.B(n_447),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_482),
.A2(n_440),
.B(n_472),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_502),
.A2(n_460),
.B1(n_438),
.B2(n_468),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_477),
.A2(n_465),
.B(n_455),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_487),
.A2(n_451),
.B1(n_454),
.B2(n_409),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_495),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_498),
.B(n_522),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_509),
.B(n_449),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

OA21x2_ASAP7_75t_L g545 ( 
.A1(n_494),
.A2(n_145),
.B(n_146),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_495),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_499),
.A2(n_147),
.B(n_148),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_520),
.A2(n_155),
.B(n_157),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_493),
.B(n_507),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_513),
.A2(n_496),
.B(n_515),
.Y(n_550)
);

AO21x2_ASAP7_75t_L g551 ( 
.A1(n_523),
.A2(n_517),
.B(n_530),
.Y(n_551)
);

A2O1A1Ixp33_ASAP7_75t_L g552 ( 
.A1(n_533),
.A2(n_484),
.B(n_479),
.C(n_531),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_503),
.B(n_500),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_L g554 ( 
.A(n_480),
.B(n_511),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_490),
.A2(n_509),
.B1(n_528),
.B2(n_533),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_478),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_483),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_519),
.A2(n_521),
.B(n_529),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_492),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_483),
.B(n_504),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_532),
.Y(n_563)
);

AO31x2_ASAP7_75t_L g564 ( 
.A1(n_518),
.A2(n_491),
.A3(n_506),
.B(n_516),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_481),
.B(n_505),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_524),
.B(n_510),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_501),
.A2(n_526),
.B(n_485),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_481),
.B(n_512),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_512),
.B(n_488),
.Y(n_569)
);

OA21x2_ASAP7_75t_L g570 ( 
.A1(n_485),
.A2(n_488),
.B(n_512),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_508),
.B(n_486),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_514),
.A2(n_488),
.B(n_508),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_514),
.A2(n_477),
.B(n_496),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

AND2x2_ASAP7_75t_SL g575 ( 
.A(n_487),
.B(n_475),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_489),
.Y(n_576)
);

AOI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_490),
.A2(n_367),
.B(n_359),
.Y(n_577)
);

AO21x2_ASAP7_75t_L g578 ( 
.A1(n_494),
.A2(n_499),
.B(n_423),
.Y(n_578)
);

OA21x2_ASAP7_75t_L g579 ( 
.A1(n_494),
.A2(n_525),
.B(n_431),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_493),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_498),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_497),
.Y(n_582)
);

CKINVDCx6p67_ASAP7_75t_R g583 ( 
.A(n_489),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_581),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_557),
.B(n_562),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_581),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_543),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_582),
.Y(n_589)
);

OA21x2_ASAP7_75t_L g590 ( 
.A1(n_572),
.A2(n_574),
.B(n_573),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_580),
.B(n_549),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_575),
.B(n_540),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_560),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_561),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_561),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_575),
.B(n_553),
.Y(n_596)
);

AO31x2_ASAP7_75t_L g597 ( 
.A1(n_538),
.A2(n_573),
.A3(n_536),
.B(n_552),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_545),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_535),
.A2(n_537),
.B(n_558),
.Y(n_599)
);

AOI21x1_ASAP7_75t_L g600 ( 
.A1(n_579),
.A2(n_538),
.B(n_567),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_545),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

CKINVDCx11_ASAP7_75t_R g605 ( 
.A(n_583),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_546),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_534),
.A2(n_550),
.B(n_548),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_579),
.A2(n_536),
.B(n_570),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_566),
.A2(n_549),
.B1(n_568),
.B2(n_565),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_557),
.B(n_555),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_569),
.A2(n_554),
.B(n_551),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_552),
.A2(n_566),
.B(n_577),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_539),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_541),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_547),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_544),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_547),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_578),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_580),
.B(n_542),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_544),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_578),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_559),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_592),
.B(n_542),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_587),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_587),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_585),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_627),
.Y(n_632)
);

NOR2x1_ASAP7_75t_L g633 ( 
.A(n_584),
.B(n_542),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_611),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_586),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_592),
.B(n_564),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_585),
.B(n_564),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_594),
.B(n_564),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_593),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_597),
.B(n_555),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_627),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_594),
.B(n_563),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_611),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_595),
.B(n_564),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_588),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_595),
.B(n_563),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_588),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_593),
.B(n_563),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_622),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_622),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_589),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_614),
.A2(n_571),
.B1(n_576),
.B2(n_559),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_610),
.B(n_576),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_589),
.B(n_571),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_591),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_596),
.B(n_617),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_623),
.B(n_571),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_623),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_612),
.B(n_586),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_625),
.B(n_597),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_602),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_597),
.B(n_615),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_603),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_606),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_597),
.B(n_624),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_615),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_624),
.B(n_616),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_597),
.B(n_613),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_608),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_618),
.B(n_620),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_598),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_673),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_656),
.B(n_621),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_639),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_655),
.B(n_626),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_658),
.B(n_621),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_659),
.B(n_626),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_634),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_658),
.B(n_619),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_661),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_646),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_634),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_629),
.B(n_619),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_631),
.Y(n_686)
);

NOR2x1_ASAP7_75t_L g687 ( 
.A(n_633),
.B(n_632),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_643),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_643),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_652),
.B(n_601),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_646),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_632),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_649),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_636),
.B(n_609),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_649),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_650),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_653),
.B(n_598),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_653),
.B(n_601),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_630),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_636),
.B(n_590),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_663),
.B(n_590),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_630),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_664),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_640),
.A2(n_600),
.B1(n_605),
.B2(n_607),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_663),
.B(n_600),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_665),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_635),
.B(n_607),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_628),
.B(n_599),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_648),
.B(n_605),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_695),
.B(n_666),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_680),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_695),
.B(n_666),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_702),
.B(n_710),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_684),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_688),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_693),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_689),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_686),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_703),
.B(n_660),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_705),
.B(n_640),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_686),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_694),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_676),
.Y(n_725)
);

NOR2x1p5_ASAP7_75t_L g726 ( 
.A(n_711),
.B(n_657),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_674),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_683),
.B(n_628),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_674),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_692),
.B(n_644),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_708),
.B(n_660),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_675),
.B(n_638),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_709),
.B(n_669),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_696),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_679),
.B(n_638),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_698),
.B(n_644),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_697),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_707),
.B(n_700),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_678),
.B(n_637),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_699),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_681),
.B(n_648),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_682),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_725),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_712),
.B(n_707),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_713),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_713),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_712),
.B(n_714),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_718),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_733),
.B(n_727),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_715),
.B(n_670),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_735),
.B(n_690),
.Y(n_752)
);

AND3x1_ASAP7_75t_L g753 ( 
.A(n_729),
.B(n_677),
.C(n_657),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_717),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_714),
.B(n_670),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_738),
.B(n_685),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_717),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_743),
.B(n_693),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_716),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_722),
.A2(n_691),
.B(n_687),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_742),
.B(n_691),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_739),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_728),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_746),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_751),
.B(n_738),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_760),
.A2(n_753),
.B(n_761),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_748),
.B(n_745),
.Y(n_767)
);

NOR2x1_ASAP7_75t_L g768 ( 
.A(n_758),
.B(n_718),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_747),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_761),
.A2(n_706),
.B(n_662),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_746),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_763),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_750),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_762),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_752),
.A2(n_654),
.B(n_642),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_R g776 ( 
.A(n_772),
.B(n_654),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_766),
.B(n_756),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_766),
.B(n_745),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_769),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_767),
.B(n_773),
.Y(n_780)
);

INVxp67_ASAP7_75t_SL g781 ( 
.A(n_774),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_764),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_771),
.Y(n_783)
);

AOI21xp33_ASAP7_75t_SL g784 ( 
.A1(n_777),
.A2(n_770),
.B(n_775),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_778),
.A2(n_770),
.B(n_775),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_781),
.A2(n_768),
.B(n_744),
.Y(n_786)
);

AOI221xp5_ASAP7_75t_L g787 ( 
.A1(n_781),
.A2(n_759),
.B1(n_757),
.B2(n_750),
.C(n_773),
.Y(n_787)
);

AOI211xp5_ASAP7_75t_SL g788 ( 
.A1(n_779),
.A2(n_730),
.B(n_731),
.C(n_739),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_L g789 ( 
.A(n_782),
.B(n_749),
.C(n_632),
.Y(n_789)
);

AOI221xp5_ASAP7_75t_L g790 ( 
.A1(n_776),
.A2(n_750),
.B1(n_719),
.B2(n_754),
.C(n_734),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_789),
.Y(n_791)
);

NOR2x1_ASAP7_75t_L g792 ( 
.A(n_786),
.B(n_783),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_784),
.B(n_785),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_787),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_790),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_793),
.B(n_780),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_792),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_795),
.B(n_788),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_794),
.B(n_765),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_797),
.B(n_791),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_799),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_798),
.B(n_726),
.Y(n_802)
);

NOR4xp75_ASAP7_75t_L g803 ( 
.A(n_796),
.B(n_641),
.C(n_748),
.D(n_732),
.Y(n_803)
);

NOR2x1_ASAP7_75t_L g804 ( 
.A(n_800),
.B(n_749),
.Y(n_804)
);

XNOR2x1_ASAP7_75t_L g805 ( 
.A(n_802),
.B(n_642),
.Y(n_805)
);

XOR2x1_ASAP7_75t_L g806 ( 
.A(n_801),
.B(n_668),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_803),
.B(n_749),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_800),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_801),
.B(n_755),
.Y(n_809)
);

XNOR2x1_ASAP7_75t_L g810 ( 
.A(n_808),
.B(n_642),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_809),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_804),
.B(n_641),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_807),
.B(n_755),
.Y(n_813)
);

AOI221xp5_ASAP7_75t_L g814 ( 
.A1(n_806),
.A2(n_671),
.B1(n_668),
.B2(n_737),
.C(n_754),
.Y(n_814)
);

OAI211xp5_ASAP7_75t_SL g815 ( 
.A1(n_805),
.A2(n_667),
.B(n_736),
.C(n_740),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_808),
.A2(n_672),
.B(n_668),
.C(n_724),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_808),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_817),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_811),
.B(n_672),
.C(n_718),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_813),
.B(n_721),
.Y(n_820)
);

AO22x2_ASAP7_75t_L g821 ( 
.A1(n_810),
.A2(n_693),
.B1(n_741),
.B2(n_724),
.Y(n_821)
);

OAI21x1_ASAP7_75t_SL g822 ( 
.A1(n_816),
.A2(n_814),
.B(n_812),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_815),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_818),
.Y(n_824)
);

AOI21xp33_ASAP7_75t_SL g825 ( 
.A1(n_823),
.A2(n_819),
.B(n_822),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_820),
.A2(n_741),
.B1(n_723),
.B2(n_720),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_821),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_823),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_824),
.A2(n_651),
.B(n_645),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_828),
.A2(n_720),
.B1(n_723),
.B2(n_733),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_827),
.A2(n_645),
.B(n_647),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_826),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_832),
.A2(n_825),
.B(n_651),
.Y(n_833)
);

AO221x1_ASAP7_75t_L g834 ( 
.A1(n_830),
.A2(n_635),
.B1(n_704),
.B2(n_701),
.C(n_647),
.Y(n_834)
);

OA21x2_ASAP7_75t_L g835 ( 
.A1(n_833),
.A2(n_831),
.B(n_829),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_835),
.B(n_834),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_836),
.A2(n_635),
.B1(n_733),
.B2(n_709),
.Y(n_837)
);


endmodule