module fake_netlist_5_1051_n_1030 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1030);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1030;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_615;
wire n_469;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1024;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_918;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_952;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_870;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_57),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_0),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_142),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_147),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_155),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_175),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_162),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_53),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_112),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_52),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_111),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_64),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_102),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_167),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_80),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_40),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_51),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_165),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_127),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_88),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_28),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_31),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_93),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_198),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_105),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_22),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_4),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_22),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_194),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_73),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_179),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_76),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_86),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_23),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_140),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_89),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_72),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_59),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_45),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_92),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_125),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_61),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_91),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_209),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_74),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_193),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_183),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_191),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_163),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_187),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_7),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_65),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_121),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_186),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_132),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_58),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_204),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_158),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_48),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_56),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_150),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_106),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_138),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_78),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_27),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_55),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_54),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_20),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_265),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_265),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_311),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_221),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_229),
.B(n_1),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_222),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_224),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_227),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_228),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_284),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_230),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_245),
.B(n_1),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_241),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_238),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_248),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_2),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_3),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_241),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_239),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_220),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_226),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_240),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_242),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_223),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_301),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_244),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_225),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_255),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_267),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_267),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_246),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_232),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_277),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_3),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_277),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_234),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_236),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_313),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_226),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_343),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_343),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_371),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_365),
.Y(n_383)
);

AND3x2_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_309),
.C(n_307),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_309),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_319),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_369),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_322),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_323),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_324),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_220),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_278),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_320),
.A2(n_312),
.B(n_243),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_329),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_359),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_350),
.Y(n_402)
);

CKINVDCx8_ASAP7_75t_R g403 ( 
.A(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_328),
.A2(n_276),
.B1(n_272),
.B2(n_294),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_335),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_344),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_231),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_347),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_356),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_361),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_332),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_318),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_359),
.B(n_250),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_360),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_355),
.B(n_312),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_363),
.B(n_251),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_341),
.B(n_237),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_342),
.B(n_249),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_348),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_254),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_220),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_374),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_235),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_310),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_258),
.Y(n_444)
);

NAND3x1_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_262),
.C(n_259),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_253),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_268),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_270),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_411),
.B(n_273),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_386),
.A2(n_308),
.B1(n_304),
.B2(n_303),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_279),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_387),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_386),
.B(n_220),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_427),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_395),
.B(n_269),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_402),
.B(n_331),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_419),
.B(n_256),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

BUFx4f_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_418),
.B(n_269),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_421),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_414),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_282),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_405),
.B(n_364),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_257),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_412),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_372),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_424),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_373),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_378),
.B(n_260),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_394),
.B(n_261),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_406),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_394),
.B(n_266),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_390),
.B(n_363),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_388),
.B(n_269),
.Y(n_493)
);

INVx4_ASAP7_75t_SL g494 ( 
.A(n_394),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_394),
.B(n_271),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_394),
.B(n_396),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_403),
.B(n_269),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_391),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_388),
.B(n_305),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_415),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_436),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_446),
.B(n_417),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_285),
.Y(n_509)
);

A2O1A1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_441),
.A2(n_274),
.B(n_275),
.C(n_280),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_479),
.B(n_281),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_283),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

NAND2x1_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_435),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_430),
.Y(n_515)
);

NAND2x1_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_435),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_480),
.A2(n_366),
.B1(n_368),
.B2(n_370),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_286),
.Y(n_518)
);

O2A1O1Ixp33_ASAP7_75t_L g519 ( 
.A1(n_459),
.A2(n_392),
.B(n_423),
.C(n_385),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_431),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_287),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_481),
.B(n_289),
.Y(n_522)
);

NOR3xp33_ASAP7_75t_L g523 ( 
.A(n_452),
.B(n_292),
.C(n_290),
.Y(n_523)
);

NOR3x1_ASAP7_75t_L g524 ( 
.A(n_458),
.B(n_317),
.C(n_316),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_466),
.A2(n_293),
.B1(n_306),
.B2(n_300),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_438),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_443),
.B(n_442),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_472),
.B(n_305),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_506),
.A2(n_370),
.B1(n_366),
.B2(n_368),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_299),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_490),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_472),
.B(n_305),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_476),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_463),
.B(n_305),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_474),
.B(n_36),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_489),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_459),
.B(n_37),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_485),
.B(n_424),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_506),
.A2(n_316),
.B1(n_317),
.B2(n_420),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_467),
.B(n_39),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_497),
.A2(n_422),
.B1(n_398),
.B2(n_377),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_382),
.Y(n_546)
);

A2O1A1Ixp33_ASAP7_75t_L g547 ( 
.A1(n_496),
.A2(n_382),
.B(n_398),
.C(n_377),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_41),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_437),
.A2(n_376),
.B1(n_6),
.B2(n_7),
.Y(n_549)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_472),
.B(n_42),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_486),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_486),
.B(n_433),
.Y(n_552)
);

AND2x6_ASAP7_75t_SL g553 ( 
.A(n_492),
.B(n_376),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_493),
.B(n_503),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_503),
.B(n_5),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_482),
.B(n_5),
.Y(n_558)
);

AND3x1_ASAP7_75t_L g559 ( 
.A(n_499),
.B(n_6),
.C(n_8),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_482),
.B(n_43),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_462),
.B(n_8),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_462),
.B(n_9),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_477),
.B(n_44),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_487),
.A2(n_118),
.B(n_217),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_477),
.B(n_47),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_437),
.B(n_49),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_434),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_437),
.B(n_50),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_437),
.B(n_60),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_499),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_473),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_501),
.B(n_9),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_501),
.B(n_10),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_444),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_468),
.Y(n_576)
);

INVx8_ASAP7_75t_L g577 ( 
.A(n_498),
.Y(n_577)
);

NAND2x1p5_ASAP7_75t_L g578 ( 
.A(n_472),
.B(n_62),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_444),
.B(n_63),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_444),
.B(n_66),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_470),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_500),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_447),
.B(n_67),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_470),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_457),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_448),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_433),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_457),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_SL g589 ( 
.A(n_505),
.B(n_10),
.C(n_11),
.Y(n_589)
);

AOI221xp5_ASAP7_75t_L g590 ( 
.A1(n_448),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_502),
.B(n_12),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_556),
.B(n_433),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_527),
.B(n_498),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_572),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_542),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_556),
.B(n_498),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_455),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_553),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_SL g600 ( 
.A(n_517),
.B(n_504),
.C(n_491),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_587),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_498),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_509),
.B(n_512),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_520),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_SL g606 ( 
.A(n_517),
.B(n_495),
.C(n_488),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_512),
.B(n_498),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_573),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_568),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_584),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_513),
.B(n_447),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_555),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_577),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_585),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_534),
.Y(n_616)
);

CKINVDCx11_ASAP7_75t_R g617 ( 
.A(n_529),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_557),
.A2(n_448),
.B(n_456),
.C(n_450),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_SL g620 ( 
.A(n_529),
.B(n_445),
.C(n_450),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

CKINVDCx8_ASAP7_75t_R g622 ( 
.A(n_582),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_546),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_450),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_SL g625 ( 
.A(n_543),
.B(n_445),
.C(n_456),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_552),
.B(n_455),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_576),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_540),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_549),
.B(n_456),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_581),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_591),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_544),
.B(n_548),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_588),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_507),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_531),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_586),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_554),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_567),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_538),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_550),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_550),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_558),
.B(n_447),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_475),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_514),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_551),
.B(n_460),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_521),
.B(n_475),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_521),
.B(n_475),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_557),
.B(n_571),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_516),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_578),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_545),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_579),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_580),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_547),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_583),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_604),
.B(n_621),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_615),
.A2(n_537),
.B(n_563),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_650),
.B(n_560),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_648),
.A2(n_575),
.B(n_469),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_615),
.A2(n_565),
.B(n_536),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_650),
.B(n_530),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_649),
.A2(n_469),
.B(n_541),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_597),
.A2(n_510),
.B(n_511),
.Y(n_666)
);

AO21x1_ASAP7_75t_L g667 ( 
.A1(n_633),
.A2(n_564),
.B(n_523),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_593),
.A2(n_522),
.B(n_518),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_633),
.A2(n_439),
.B(n_566),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_612),
.A2(n_439),
.B(n_569),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_630),
.A2(n_549),
.B(n_590),
.C(n_574),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_627),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_609),
.B(n_523),
.Y(n_673)
);

NAND2x1p5_ASAP7_75t_L g674 ( 
.A(n_614),
.B(n_460),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_608),
.A2(n_449),
.B(n_440),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_638),
.Y(n_676)
);

AO21x1_ASAP7_75t_L g677 ( 
.A1(n_630),
.A2(n_570),
.B(n_519),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_593),
.B(n_525),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_615),
.A2(n_440),
.B(n_449),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_652),
.A2(n_451),
.B(n_528),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_614),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_636),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_618),
.A2(n_528),
.B(n_533),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_637),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_644),
.A2(n_545),
.B1(n_526),
.B2(n_543),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_632),
.B(n_561),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_653),
.B(n_595),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_645),
.B(n_464),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_641),
.B(n_464),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_596),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_641),
.B(n_465),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_623),
.Y(n_692)
);

OAI21x1_ASAP7_75t_SL g693 ( 
.A1(n_643),
.A2(n_451),
.B(n_559),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_603),
.A2(n_533),
.B(n_562),
.C(n_589),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_607),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_601),
.B(n_465),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_618),
.A2(n_465),
.B(n_589),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_654),
.B(n_478),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_656),
.B(n_465),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_627),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_628),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_594),
.A2(n_655),
.B(n_652),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_655),
.A2(n_634),
.B(n_631),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_602),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_607),
.A2(n_457),
.B(n_478),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_631),
.A2(n_465),
.B(n_471),
.Y(n_706)
);

AOI21x1_ASAP7_75t_L g707 ( 
.A1(n_610),
.A2(n_457),
.B(n_478),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_635),
.A2(n_494),
.B(n_478),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_653),
.A2(n_524),
.B1(n_14),
.B2(n_15),
.Y(n_709)
);

AO21x1_ASAP7_75t_L g710 ( 
.A1(n_643),
.A2(n_13),
.B(n_15),
.Y(n_710)
);

AOI31xp33_ASAP7_75t_L g711 ( 
.A1(n_599),
.A2(n_16),
.A3(n_17),
.B(n_18),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_623),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_607),
.A2(n_494),
.B(n_471),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_659),
.B(n_657),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_672),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_679),
.A2(n_635),
.B(n_640),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_672),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_665),
.A2(n_643),
.B(n_624),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_692),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_690),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_700),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_700),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_675),
.A2(n_635),
.B(n_640),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_600),
.B(n_606),
.C(n_625),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_682),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_681),
.B(n_598),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_684),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_695),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_663),
.A2(n_640),
.B(n_639),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_704),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_690),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_685),
.B(n_620),
.C(n_617),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_676),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_664),
.B(n_634),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_701),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_687),
.B(n_622),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_680),
.A2(n_660),
.B(n_707),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_680),
.A2(n_639),
.B(n_611),
.Y(n_738)
);

AO21x2_ASAP7_75t_L g739 ( 
.A1(n_666),
.A2(n_629),
.B(n_592),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_669),
.A2(n_592),
.B(n_613),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_661),
.B(n_598),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_702),
.A2(n_613),
.B(n_651),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_708),
.A2(n_651),
.B(n_646),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_667),
.A2(n_646),
.A3(n_642),
.B(n_624),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_671),
.A2(n_616),
.B1(n_626),
.B2(n_598),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_695),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_681),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_708),
.A2(n_642),
.B(n_624),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_668),
.A2(n_624),
.B(n_642),
.Y(n_749)
);

NOR4xp25_ASAP7_75t_L g750 ( 
.A(n_709),
.B(n_617),
.C(n_622),
.D(n_605),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_689),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_712),
.Y(n_752)
);

OA21x2_ASAP7_75t_L g753 ( 
.A1(n_697),
.A2(n_647),
.B(n_626),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_686),
.A2(n_626),
.B1(n_647),
.B2(n_599),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_670),
.A2(n_642),
.B(n_619),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_687),
.B(n_678),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_676),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_703),
.A2(n_619),
.B(n_614),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_683),
.A2(n_619),
.B(n_614),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_694),
.A2(n_647),
.B(n_619),
.C(n_18),
.Y(n_760)
);

OA21x2_ASAP7_75t_L g761 ( 
.A1(n_662),
.A2(n_471),
.B(n_494),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_705),
.A2(n_471),
.B(n_131),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_698),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_691),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_718),
.A2(n_677),
.B(n_698),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_719),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_747),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_727),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_750),
.A2(n_709),
.B1(n_711),
.B2(n_673),
.C(n_694),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_756),
.B(n_681),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_719),
.Y(n_771)
);

OAI221xp5_ASAP7_75t_L g772 ( 
.A1(n_724),
.A2(n_688),
.B1(n_699),
.B2(n_696),
.C(n_706),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_714),
.A2(n_681),
.B1(n_674),
.B2(n_710),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_735),
.A2(n_674),
.B1(n_713),
.B2(n_693),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_749),
.A2(n_471),
.B(n_133),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_727),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_714),
.B(n_16),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_741),
.B(n_17),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_726),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_733),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_726),
.B(n_68),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_757),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_741),
.B(n_734),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_725),
.Y(n_784)
);

OAI222xp33_ASAP7_75t_L g785 ( 
.A1(n_735),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.C1(n_23),
.C2(n_24),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_734),
.B(n_21),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_R g787 ( 
.A(n_736),
.B(n_69),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_732),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_715),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_SL g790 ( 
.A1(n_745),
.A2(n_752),
.B1(n_753),
.B2(n_733),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_754),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_720),
.A2(n_731),
.B1(n_752),
.B2(n_753),
.Y(n_792)
);

AND2x6_ASAP7_75t_L g793 ( 
.A(n_747),
.B(n_70),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_720),
.B(n_71),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_725),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_731),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_760),
.B(n_75),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_730),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_753),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_726),
.B(n_747),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_SL g801 ( 
.A1(n_753),
.A2(n_751),
.B1(n_747),
.B2(n_763),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_747),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_751),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_715),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_746),
.B(n_77),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_737),
.A2(n_149),
.B(n_216),
.Y(n_806)
);

AO21x2_ASAP7_75t_L g807 ( 
.A1(n_737),
.A2(n_729),
.B(n_739),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_717),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_717),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_721),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_728),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_729),
.A2(n_755),
.B(n_740),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_746),
.B(n_79),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_763),
.A2(n_35),
.B1(n_81),
.B2(n_82),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_721),
.Y(n_815)
);

OAI221xp5_ASAP7_75t_L g816 ( 
.A1(n_764),
.A2(n_83),
.B1(n_85),
.B2(n_87),
.C(n_90),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_728),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_722),
.B(n_95),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_722),
.B(n_218),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_764),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_755),
.A2(n_96),
.B(n_98),
.Y(n_821)
);

NAND3xp33_ASAP7_75t_SL g822 ( 
.A(n_739),
.B(n_101),
.C(n_103),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_769),
.A2(n_761),
.B1(n_744),
.B2(n_759),
.Y(n_823)
);

CKINVDCx11_ASAP7_75t_R g824 ( 
.A(n_771),
.Y(n_824)
);

OAI221xp5_ASAP7_75t_L g825 ( 
.A1(n_788),
.A2(n_761),
.B1(n_744),
.B2(n_739),
.C(n_759),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_767),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_783),
.B(n_744),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_800),
.B(n_748),
.Y(n_828)
);

AOI221xp5_ASAP7_75t_L g829 ( 
.A1(n_788),
.A2(n_744),
.B1(n_738),
.B2(n_740),
.C(n_742),
.Y(n_829)
);

AOI222xp33_ASAP7_75t_L g830 ( 
.A1(n_785),
.A2(n_742),
.B1(n_738),
.B2(n_762),
.C1(n_723),
.C2(n_758),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_796),
.A2(n_762),
.B1(n_723),
.B2(n_761),
.Y(n_831)
);

INVx3_ASAP7_75t_SL g832 ( 
.A(n_780),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_776),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_778),
.B(n_744),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_777),
.B(n_758),
.Y(n_835)
);

OAI22xp33_ASAP7_75t_L g836 ( 
.A1(n_787),
.A2(n_761),
.B1(n_748),
.B2(n_716),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_797),
.A2(n_716),
.B1(n_743),
.B2(n_108),
.Y(n_837)
);

AO22x1_ASAP7_75t_L g838 ( 
.A1(n_793),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_791),
.A2(n_743),
.B1(n_113),
.B2(n_114),
.Y(n_839)
);

OAI221xp5_ASAP7_75t_L g840 ( 
.A1(n_797),
.A2(n_110),
.B1(n_115),
.B2(n_116),
.C(n_117),
.Y(n_840)
);

AOI221xp5_ASAP7_75t_L g841 ( 
.A1(n_799),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.C(n_124),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_770),
.A2(n_126),
.B(n_129),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_797),
.A2(n_130),
.B1(n_135),
.B2(n_136),
.Y(n_843)
);

NOR2x1_ASAP7_75t_SL g844 ( 
.A(n_822),
.B(n_137),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_784),
.Y(n_845)
);

AOI21xp33_ASAP7_75t_L g846 ( 
.A1(n_773),
.A2(n_139),
.B(n_141),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_790),
.B(n_143),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_799),
.A2(n_215),
.B1(n_146),
.B2(n_148),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_775),
.A2(n_765),
.B(n_816),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_803),
.A2(n_144),
.B1(n_151),
.B2(n_152),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_786),
.B(n_153),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_803),
.A2(n_154),
.B1(n_156),
.B2(n_159),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_766),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_821),
.B(n_160),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_795),
.Y(n_855)
);

OAI211xp5_ASAP7_75t_L g856 ( 
.A1(n_809),
.A2(n_814),
.B(n_794),
.C(n_782),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_812),
.A2(n_161),
.B(n_164),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_780),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_767),
.Y(n_859)
);

AOI221xp5_ASAP7_75t_L g860 ( 
.A1(n_809),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.C(n_171),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_798),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_798),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_805),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_863)
);

AO21x2_ASAP7_75t_L g864 ( 
.A1(n_765),
.A2(n_177),
.B(n_178),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_779),
.B(n_180),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_767),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_L g867 ( 
.A1(n_792),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.C(n_188),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_805),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_847),
.A2(n_793),
.B1(n_813),
.B2(n_781),
.Y(n_869)
);

AO31x2_ASAP7_75t_L g870 ( 
.A1(n_823),
.A2(n_774),
.A3(n_815),
.B(n_820),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_827),
.B(n_801),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_834),
.B(n_807),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_845),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_861),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_855),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_862),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_835),
.B(n_807),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_828),
.B(n_820),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_833),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_828),
.B(n_768),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_825),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_858),
.B(n_808),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_853),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_832),
.B(n_810),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_864),
.B(n_779),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_864),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_857),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_836),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_832),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_866),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_836),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_854),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_854),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_866),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_831),
.B(n_804),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_830),
.B(n_789),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_866),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_854),
.B(n_800),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_831),
.B(n_819),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_844),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_866),
.Y(n_902)
);

AO21x2_ASAP7_75t_L g903 ( 
.A1(n_886),
.A2(n_849),
.B(n_846),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_873),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_890),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_R g906 ( 
.A(n_893),
.B(n_824),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_890),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_873),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_872),
.B(n_848),
.Y(n_909)
);

AOI211xp5_ASAP7_75t_L g910 ( 
.A1(n_887),
.A2(n_840),
.B(n_856),
.C(n_838),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_869),
.A2(n_843),
.B1(n_848),
.B2(n_850),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_883),
.B(n_851),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_872),
.B(n_837),
.Y(n_913)
);

OAI321xp33_ASAP7_75t_L g914 ( 
.A1(n_887),
.A2(n_843),
.A3(n_852),
.B1(n_841),
.B2(n_839),
.C(n_860),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_885),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_884),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_886),
.A2(n_806),
.B(n_842),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_893),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_881),
.A2(n_850),
.B(n_852),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_875),
.Y(n_920)
);

OAI221xp5_ASAP7_75t_L g921 ( 
.A1(n_881),
.A2(n_839),
.B1(n_868),
.B2(n_863),
.C(n_867),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_SL g922 ( 
.A1(n_894),
.A2(n_793),
.B1(n_859),
.B2(n_781),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_894),
.A2(n_774),
.B(n_772),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_875),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_916),
.B(n_871),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_924),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_904),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_918),
.B(n_871),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_904),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_918),
.B(n_877),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_924),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_908),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_907),
.B(n_901),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_908),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_915),
.B(n_877),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_915),
.B(n_892),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_905),
.B(n_889),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_906),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_939),
.A2(n_911),
.B1(n_919),
.B2(n_921),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_926),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_937),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_925),
.B(n_909),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_927),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_932),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_938),
.B(n_909),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_930),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_941),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_945),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_947),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_944),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_914),
.C(n_919),
.Y(n_952)
);

AOI31xp33_ASAP7_75t_L g953 ( 
.A1(n_940),
.A2(n_910),
.A3(n_922),
.B(n_934),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_944),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_943),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_955),
.B(n_942),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_948),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_953),
.B(n_934),
.Y(n_958)
);

AOI221xp5_ASAP7_75t_L g959 ( 
.A1(n_952),
.A2(n_940),
.B1(n_910),
.B2(n_914),
.C(n_923),
.Y(n_959)
);

NOR2x1p5_ASAP7_75t_L g960 ( 
.A(n_950),
.B(n_915),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_958),
.B(n_953),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_SL g962 ( 
.A1(n_959),
.A2(n_913),
.B(n_912),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_956),
.B(n_949),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_957),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_963),
.B(n_954),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_964),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_961),
.B(n_960),
.Y(n_967)
);

XNOR2xp5_ASAP7_75t_L g968 ( 
.A(n_962),
.B(n_922),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_963),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_969),
.B(n_951),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_966),
.B(n_929),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_936),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_968),
.B(n_937),
.Y(n_973)
);

AOI211xp5_ASAP7_75t_L g974 ( 
.A1(n_965),
.A2(n_901),
.B(n_913),
.C(n_889),
.Y(n_974)
);

AOI31xp33_ASAP7_75t_L g975 ( 
.A1(n_969),
.A2(n_884),
.A3(n_882),
.B(n_931),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_966),
.B(n_892),
.C(n_882),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_969),
.B(n_900),
.C(n_897),
.Y(n_977)
);

NAND4xp25_ASAP7_75t_SL g978 ( 
.A(n_974),
.B(n_936),
.C(n_900),
.D(n_897),
.Y(n_978)
);

NAND4xp25_ASAP7_75t_L g979 ( 
.A(n_970),
.B(n_899),
.C(n_876),
.D(n_826),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_977),
.A2(n_903),
.B(n_876),
.Y(n_980)
);

NAND4xp25_ASAP7_75t_L g981 ( 
.A(n_973),
.B(n_899),
.C(n_826),
.D(n_915),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_975),
.B(n_874),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_L g983 ( 
.A(n_971),
.B(n_865),
.C(n_818),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_976),
.A2(n_903),
.B(n_886),
.C(n_813),
.Y(n_984)
);

AOI221xp5_ASAP7_75t_L g985 ( 
.A1(n_972),
.A2(n_903),
.B1(n_874),
.B2(n_930),
.C(n_928),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_982),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_979),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_978),
.B(n_983),
.Y(n_989)
);

XNOR2xp5_ASAP7_75t_L g990 ( 
.A(n_980),
.B(n_899),
.Y(n_990)
);

NAND4xp75_ASAP7_75t_L g991 ( 
.A(n_985),
.B(n_793),
.C(n_818),
.D(n_819),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_984),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_980),
.A2(n_917),
.B(n_899),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_986),
.B(n_987),
.C(n_988),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_992),
.Y(n_995)
);

NOR2x1_ASAP7_75t_L g996 ( 
.A(n_989),
.B(n_802),
.Y(n_996)
);

AOI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_990),
.A2(n_195),
.B(n_196),
.Y(n_997)
);

OA22x2_ASAP7_75t_L g998 ( 
.A1(n_993),
.A2(n_991),
.B1(n_898),
.B2(n_895),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_993),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_986),
.A2(n_935),
.B1(n_933),
.B2(n_928),
.Y(n_1000)
);

NOR4xp75_ASAP7_75t_L g1001 ( 
.A(n_991),
.B(n_878),
.C(n_880),
.D(n_902),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_994),
.A2(n_888),
.B(n_879),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_999),
.B(n_802),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

NOR4xp25_ASAP7_75t_L g1005 ( 
.A(n_995),
.B(n_935),
.C(n_933),
.D(n_927),
.Y(n_1005)
);

NAND5xp2_ASAP7_75t_L g1006 ( 
.A(n_998),
.B(n_878),
.C(n_880),
.D(n_879),
.E(n_902),
.Y(n_1006)
);

NAND4xp25_ASAP7_75t_L g1007 ( 
.A(n_997),
.B(n_898),
.C(n_896),
.D(n_888),
.Y(n_1007)
);

OA22x2_ASAP7_75t_L g1008 ( 
.A1(n_1000),
.A2(n_891),
.B1(n_885),
.B2(n_920),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1001),
.Y(n_1009)
);

AND3x4_ASAP7_75t_L g1010 ( 
.A(n_1009),
.B(n_885),
.C(n_920),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1004),
.A2(n_920),
.B1(n_908),
.B2(n_896),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_1003),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1008),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1007),
.A2(n_1002),
.B1(n_1005),
.B2(n_1006),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_1004),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_1015),
.A2(n_917),
.B(n_885),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1013),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_1012),
.B(n_870),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1017),
.B(n_1014),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1018),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1019),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_1020),
.B(n_1010),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_1022),
.B(n_1016),
.C(n_1011),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1021),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1024),
.A2(n_802),
.B1(n_917),
.B2(n_811),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1023),
.A2(n_917),
.B(n_199),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_L g1027 ( 
.A(n_1026),
.B(n_197),
.C(n_200),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_SL g1028 ( 
.A(n_1025),
.B(n_201),
.C(n_202),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_1027),
.A2(n_203),
.B1(n_212),
.B2(n_213),
.C(n_214),
.Y(n_1029)
);

AOI211xp5_ASAP7_75t_L g1030 ( 
.A1(n_1029),
.A2(n_1028),
.B(n_811),
.C(n_817),
.Y(n_1030)
);


endmodule