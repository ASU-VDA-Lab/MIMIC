module fake_jpeg_7876_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_41),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_42),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_25),
.A2(n_8),
.B(n_15),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_27),
.B1(n_20),
.B2(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_28),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_25),
.B1(n_35),
.B2(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_69),
.B1(n_72),
.B2(n_36),
.Y(n_97)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_66),
.Y(n_93)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_25),
.B1(n_35),
.B2(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_35),
.B1(n_27),
.B2(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_27),
.B1(n_36),
.B2(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_86),
.B(n_90),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_82),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_99),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_119),
.B1(n_19),
.B2(n_21),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_21),
.B1(n_19),
.B2(n_23),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_78),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_120),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_33),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_115),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_31),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_31),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_65),
.B(n_17),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_34),
.B1(n_28),
.B2(n_29),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_21),
.B1(n_23),
.B2(n_9),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_32),
.B1(n_30),
.B2(n_17),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_58),
.B(n_32),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_22),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_55),
.B(n_24),
.Y(n_124)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_22),
.B(n_21),
.C(n_24),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_115),
.A3(n_108),
.B1(n_99),
.B2(n_111),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_123),
.B(n_93),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_115),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_146),
.B1(n_111),
.B2(n_117),
.Y(n_159)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_145),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_94),
.B1(n_88),
.B2(n_113),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_21),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_0),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_23),
.B1(n_9),
.B2(n_11),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_154),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_23),
.B1(n_9),
.B2(n_11),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_107),
.B1(n_100),
.B2(n_95),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_110),
.B(n_23),
.CI(n_1),
.CON(n_151),
.SN(n_151)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_151),
.B(n_13),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_102),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_136),
.B(n_151),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_163),
.B(n_165),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_186),
.B1(n_190),
.B2(n_176),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_160),
.A2(n_176),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_171),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_108),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_175),
.B1(n_133),
.B2(n_126),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_95),
.B(n_109),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_129),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_183),
.Y(n_204)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_89),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_170),
.B(n_174),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_178),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_121),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_109),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_181),
.B(n_184),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_113),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_179),
.B(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_152),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_138),
.B(n_135),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_186),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_132),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_94),
.B1(n_143),
.B2(n_126),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_189),
.B(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_159),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_203),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_184),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_195),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_153),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_156),
.C(n_155),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_199),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_156),
.C(n_155),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_202),
.B1(n_175),
.B2(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_206),
.B(n_212),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_210),
.A2(n_220),
.B(n_200),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_216),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_162),
.A2(n_127),
.A3(n_143),
.B1(n_15),
.B2(n_16),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_133),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_104),
.B(n_87),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_183),
.B1(n_168),
.B2(n_188),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_158),
.B1(n_165),
.B2(n_181),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_225),
.A2(n_246),
.B1(n_192),
.B2(n_218),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_158),
.B(n_163),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_244),
.B(n_199),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_232),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_235),
.B1(n_249),
.B2(n_205),
.Y(n_250)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_230),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_191),
.A3(n_222),
.B1(n_215),
.B2(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_160),
.B1(n_187),
.B2(n_163),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_180),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_195),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_8),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_215),
.B(n_214),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_167),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_201),
.C(n_197),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_91),
.B(n_106),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_265),
.B1(n_225),
.B2(n_239),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_261),
.C(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_260),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_266),
.B(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_240),
.C(n_241),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_241),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_211),
.C(n_198),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_269),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_203),
.B1(n_208),
.B2(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_219),
.B1(n_196),
.B2(n_193),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_243),
.B1(n_235),
.B2(n_242),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_270),
.B1(n_267),
.B2(n_266),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_252),
.B1(n_254),
.B2(n_268),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.C(n_263),
.Y(n_290)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_226),
.C(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_249),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_250),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_286),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_252),
.A2(n_230),
.B1(n_196),
.B2(n_8),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_287),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_259),
.B(n_230),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_255),
.B(n_6),
.Y(n_289)
);

AOI221xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_4),
.B1(n_6),
.B2(n_12),
.C(n_14),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_279),
.C(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_300),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_251),
.B(n_253),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_276),
.B(n_278),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_262),
.B1(n_2),
.B2(n_3),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_274),
.B(n_281),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_7),
.B1(n_13),
.B2(n_4),
.Y(n_300)
);

BUFx12_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_288),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_280),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_307),
.C(n_314),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_280),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_291),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_301),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_278),
.B(n_275),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_315),
.Y(n_325)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_273),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_315),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_302),
.B1(n_292),
.B2(n_295),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_318),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_296),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_324),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_302),
.B1(n_299),
.B2(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_285),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_296),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_322),
.B(n_325),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_307),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_314),
.C(n_305),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_327),
.C(n_326),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_338),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_316),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_333),
.B(n_304),
.Y(n_341)
);


endmodule