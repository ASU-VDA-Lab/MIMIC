module fake_ariane_2365_n_300 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_54, n_25, n_300);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_54;
input n_25;

output n_300;

wire n_295;
wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_289;
wire n_288;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_294;
wire n_110;
wire n_153;
wire n_221;
wire n_197;
wire n_86;
wire n_269;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_259;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_299;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_111;
wire n_242;
wire n_260;
wire n_274;
wire n_115;
wire n_272;
wire n_133;
wire n_66;
wire n_205;
wire n_236;
wire n_265;
wire n_71;
wire n_267;
wire n_109;
wire n_208;
wire n_245;
wire n_96;
wire n_156;
wire n_281;
wire n_209;
wire n_262;
wire n_291;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_283;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_235;
wire n_225;
wire n_200;
wire n_297;
wire n_166;
wire n_253;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_244;
wire n_246;
wire n_226;
wire n_271;
wire n_290;
wire n_220;
wire n_84;
wire n_261;
wire n_247;
wire n_199;
wire n_91;
wire n_189;
wire n_107;
wire n_159;
wire n_72;
wire n_128;
wire n_105;
wire n_217;
wire n_224;
wire n_240;
wire n_82;
wire n_178;
wire n_286;
wire n_57;
wire n_131;
wire n_263;
wire n_201;
wire n_229;
wire n_70;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_287;
wire n_85;
wire n_130;
wire n_144;
wire n_256;
wire n_214;
wire n_227;
wire n_94;
wire n_101;
wire n_243;
wire n_284;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_162;
wire n_112;
wire n_138;
wire n_278;
wire n_264;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_282;
wire n_122;
wire n_268;
wire n_257;
wire n_266;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_277;
wire n_157;
wire n_248;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_73;
wire n_77;
wire n_293;
wire n_171;
wire n_228;
wire n_121;
wire n_118;
wire n_93;
wire n_276;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_279;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_219;
wire n_140;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_270;
wire n_194;
wire n_97;
wire n_154;
wire n_280;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_285;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_298;
wire n_296;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_59;
wire n_63;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_273;

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_86),
.Y(n_115)
);

NAND2x1_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_102),
.Y(n_117)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_76),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_84),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_58),
.B1(n_63),
.B2(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_75),
.Y(n_123)
);

AO221x1_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_78),
.B1(n_74),
.B2(n_71),
.C(n_63),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_77),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_33),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_3),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_110),
.B1(n_109),
.B2(n_92),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_110),
.B1(n_106),
.B2(n_107),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_96),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_117),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_125),
.B1(n_130),
.B2(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_99),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_98),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_112),
.B1(n_118),
.B2(n_88),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_99),
.B(n_98),
.C(n_95),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_112),
.B1(n_92),
.B2(n_95),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_112),
.B1(n_88),
.B2(n_89),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_95),
.B(n_92),
.C(n_103),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_112),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_92),
.B1(n_95),
.B2(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_91),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_91),
.Y(n_167)
);

O2A1O1Ixp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_105),
.B(n_100),
.C(n_94),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_95),
.B1(n_92),
.B2(n_89),
.Y(n_176)
);

AOI222xp33_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_142),
.B1(n_137),
.B2(n_146),
.C1(n_148),
.C2(n_89),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_138),
.B1(n_142),
.B2(n_135),
.Y(n_181)
);

BUFx4f_ASAP7_75t_SL g182 ( 
.A(n_154),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_169),
.B1(n_155),
.B2(n_164),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_164),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_157),
.C(n_161),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_174),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_177),
.B1(n_181),
.B2(n_178),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_175),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_176),
.B(n_159),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_174),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_168),
.Y(n_212)
);

NAND4xp25_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_173),
.C(n_183),
.D(n_10),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_205),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_205),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_183),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_194),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_194),
.Y(n_224)
);

AOI33xp33_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_192),
.A3(n_10),
.B1(n_8),
.B2(n_158),
.B3(n_150),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_212),
.B1(n_203),
.B2(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_210),
.A3(n_211),
.B1(n_208),
.B2(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_220),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_214),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_207),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_226),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_220),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_226),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_219),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_219),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_196),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_208),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_R g254 ( 
.A(n_236),
.B(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_216),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_216),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_216),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_197),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_250),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_245),
.C(n_201),
.Y(n_269)
);

NOR3x1_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_251),
.C(n_253),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_261),
.C(n_260),
.Y(n_271)
);

AOI221xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_252),
.B1(n_240),
.B2(n_89),
.C(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_243),
.Y(n_273)
);

AOI222xp33_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_263),
.B1(n_89),
.B2(n_267),
.C1(n_264),
.C2(n_259),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_199),
.A3(n_257),
.B1(n_264),
.B2(n_254),
.C1(n_247),
.C2(n_151),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_254),
.B(n_247),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_209),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

NAND4xp25_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_273),
.C(n_268),
.D(n_150),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_276),
.B1(n_191),
.B2(n_209),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

AOI222xp33_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_191),
.B1(n_171),
.B2(n_149),
.C1(n_209),
.C2(n_20),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_14),
.Y(n_285)
);

NOR2x1p5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_171),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_15),
.C(n_17),
.Y(n_287)
);

AO22x2_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_29),
.C(n_30),
.Y(n_289)
);

NAND5xp2_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_31),
.C(n_32),
.D(n_35),
.E(n_36),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_40),
.C(n_41),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

OAI222xp33_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.C1(n_46),
.C2(n_48),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_49),
.B(n_50),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_171),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_295),
.B(n_292),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_282),
.B(n_293),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_298),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_297),
.B(n_296),
.Y(n_300)
);


endmodule