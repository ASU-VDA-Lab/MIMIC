module fake_ariane_1196_n_3095 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_3095);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_3095;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_3063;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_1491;
wire n_931;
wire n_2628;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3052;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_2853;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_3085;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2723;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_943;
wire n_2905;
wire n_2884;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_1321;
wire n_3050;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2700;
wire n_2606;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_1116;
wire n_3043;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_2974;
wire n_923;
wire n_1645;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_3091;
wire n_1024;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_898;
wire n_857;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_2967;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_3018;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2705;
wire n_2664;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_2917;
wire n_2544;
wire n_2085;
wire n_2432;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3094;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2678;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_815),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_753),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_803),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_666),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_835),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_295),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_218),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_584),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_144),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_475),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_777),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_671),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_771),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_414),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_579),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_821),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_339),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_665),
.Y(n_858)
);

BUFx8_ASAP7_75t_SL g859 ( 
.A(n_39),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_408),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_764),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_66),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_720),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_691),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_238),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_793),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_460),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_388),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_832),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_410),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_807),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_768),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_356),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_392),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_617),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_165),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_188),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_4),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_68),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_521),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_236),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_679),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_758),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_798),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_594),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_783),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_469),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_759),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_100),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_762),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_139),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_320),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_792),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_175),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_755),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_50),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_499),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_761),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_787),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_809),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_402),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_548),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_409),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_77),
.Y(n_904)
);

BUFx2_ASAP7_75t_SL g905 ( 
.A(n_383),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_659),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_483),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_488),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_672),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_215),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_667),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_436),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_389),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_752),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_351),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_784),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_300),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_167),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_642),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_168),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_543),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_403),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_630),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_749),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_37),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_362),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_786),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_57),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_765),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_702),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_781),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_553),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_466),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_270),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_61),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_673),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_561),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_804),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_649),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_205),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_828),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_234),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_801),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_154),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_611),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_776),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_819),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_284),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_355),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_827),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_710),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_567),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_18),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_120),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_839),
.Y(n_955)
);

CKINVDCx16_ASAP7_75t_R g956 ( 
.A(n_773),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_241),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_600),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_275),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_526),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_775),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_779),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_825),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_181),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_778),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_411),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_806),
.Y(n_967)
);

INVxp33_ASAP7_75t_SL g968 ( 
.A(n_132),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_441),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_121),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_785),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_255),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_791),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_829),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_15),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_357),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_450),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_474),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_13),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_287),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_831),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_162),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_49),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_103),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_747),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_644),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_619),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_46),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_665),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_109),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_183),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_474),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_730),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_627),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_706),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_780),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_20),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_249),
.Y(n_998)
);

CKINVDCx14_ASAP7_75t_R g999 ( 
.A(n_587),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_811),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_247),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_444),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_141),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_693),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_95),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_189),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_523),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_501),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_556),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_490),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_276),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_413),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_805),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_757),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_558),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_660),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_529),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_822),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_602),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_394),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_756),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_91),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_838),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_476),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_411),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_162),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_737),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_14),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_810),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_531),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_98),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_90),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_366),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_544),
.Y(n_1034)
);

BUFx5_ASAP7_75t_L g1035 ( 
.A(n_840),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_76),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_782),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_788),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_470),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_541),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_597),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_227),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_366),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_384),
.Y(n_1044)
);

CKINVDCx14_ASAP7_75t_R g1045 ( 
.A(n_52),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_772),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_237),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_790),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_774),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_607),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_797),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_90),
.Y(n_1052)
);

CKINVDCx14_ASAP7_75t_R g1053 ( 
.A(n_83),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_255),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_802),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_260),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_817),
.Y(n_1057)
);

CKINVDCx14_ASAP7_75t_R g1058 ( 
.A(n_28),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_456),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_113),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_823),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_11),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_554),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_607),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_374),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_672),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_269),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_48),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_359),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_662),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_670),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_403),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_11),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_431),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_418),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_40),
.Y(n_1076)
);

BUFx10_ASAP7_75t_L g1077 ( 
.A(n_769),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_598),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_268),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_242),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_559),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_92),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_267),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_697),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_483),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_669),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_208),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_824),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_305),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_201),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_86),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_107),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_818),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_124),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_541),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_31),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_3),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_808),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_285),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_796),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_813),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_751),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_71),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_84),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_767),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_445),
.Y(n_1106)
);

CKINVDCx14_ASAP7_75t_R g1107 ( 
.A(n_175),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_538),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_493),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_816),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_356),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_712),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_132),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_766),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_826),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_511),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_454),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_341),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_613),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_675),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_267),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_482),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_836),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_246),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_452),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_24),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_800),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_760),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_794),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_244),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_750),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_592),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_362),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_789),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_389),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_248),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_32),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_149),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_128),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_578),
.Y(n_1140)
);

BUFx5_ASAP7_75t_L g1141 ( 
.A(n_321),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_671),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_820),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_837),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_276),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_763),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_687),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_119),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_799),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_550),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_278),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_686),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_664),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_93),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_795),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_122),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_668),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_333),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_41),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_277),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_812),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_548),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_770),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_197),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_112),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_76),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_583),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_739),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_655),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_44),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_21),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_151),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_834),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_103),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_833),
.Y(n_1175)
);

BUFx10_ASAP7_75t_L g1176 ( 
.A(n_334),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_754),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_830),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_381),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_594),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_485),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_814),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_0),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_140),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_1042),
.Y(n_1185)
);

INVxp33_ASAP7_75t_SL g1186 ( 
.A(n_1092),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1042),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1141),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1141),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1141),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1141),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1141),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_844),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_850),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1007),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_873),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_874),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_859),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_898),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_999),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_892),
.Y(n_1201)
);

INVxp33_ASAP7_75t_SL g1202 ( 
.A(n_1017),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_896),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_901),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_930),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_902),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_950),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_909),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_963),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_848),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_910),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_912),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_913),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_848),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_919),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_1045),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_920),
.Y(n_1217)
);

INVxp33_ASAP7_75t_SL g1218 ( 
.A(n_1062),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_926),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_1053),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_928),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_933),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_944),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_952),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_848),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1058),
.Y(n_1226)
);

INVxp33_ASAP7_75t_SL g1227 ( 
.A(n_905),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_906),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_906),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_954),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_972),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1021),
.Y(n_1232)
);

INVxp33_ASAP7_75t_SL g1233 ( 
.A(n_846),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_975),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_906),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_977),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1107),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_983),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_990),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1001),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1114),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1152),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1188),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1210),
.Y(n_1244)
);

AOI22x1_ASAP7_75t_SL g1245 ( 
.A1(n_1199),
.A2(n_921),
.B1(n_925),
.B2(n_855),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1214),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1225),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1229),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1195),
.A2(n_994),
.B1(n_1009),
.B2(n_966),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1228),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1185),
.B(n_1146),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1235),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1187),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1198),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1189),
.B(n_1190),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1191),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1192),
.A2(n_863),
.B(n_842),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1194),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1196),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1233),
.B(n_956),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1197),
.Y(n_1261)
);

BUFx8_ASAP7_75t_L g1262 ( 
.A(n_1207),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1201),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1200),
.A2(n_1025),
.B1(n_1066),
.B2(n_1043),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1220),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1203),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1204),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1205),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1206),
.A2(n_883),
.B(n_869),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1195),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1193),
.A2(n_1074),
.B1(n_1109),
.B2(n_1080),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1242),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1208),
.B(n_1057),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1211),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1212),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1213),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1215),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1217),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1222),
.B(n_1237),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1219),
.B(n_884),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1209),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1222),
.B(n_889),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1232),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1221),
.Y(n_1284)
);

BUFx8_ASAP7_75t_L g1285 ( 
.A(n_1223),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1224),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1216),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1268),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1252),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1254),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1281),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1253),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1259),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1283),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1262),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1287),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1263),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1267),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1273),
.B(n_1227),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1260),
.A2(n_1218),
.B1(n_1202),
.B2(n_1186),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1272),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1272),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1252),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1286),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1265),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1265),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1271),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1249),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1266),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1270),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1274),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1270),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1264),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1275),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1279),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1277),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1284),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1285),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1245),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1258),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1256),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1261),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1261),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1251),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1248),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_R g1326 ( 
.A(n_1244),
.B(n_1241),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1282),
.B(n_1226),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1255),
.A2(n_893),
.B(n_888),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1276),
.B(n_1230),
.Y(n_1329)
);

NAND2xp33_ASAP7_75t_R g1330 ( 
.A(n_1257),
.B(n_968),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1243),
.B(n_1231),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1276),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1278),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1278),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1246),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1247),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1250),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1269),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1280),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1253),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1252),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1268),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1268),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1268),
.B(n_1129),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1268),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1270),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1253),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1253),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1268),
.Y(n_1349)
);

NOR2xp67_ASAP7_75t_L g1350 ( 
.A(n_1265),
.B(n_1234),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1268),
.Y(n_1351)
);

NOR2xp67_ASAP7_75t_L g1352 ( 
.A(n_1265),
.B(n_1236),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1293),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1301),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1321),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1302),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1290),
.B(n_1238),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1299),
.B(n_923),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1309),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1297),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1288),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1339),
.B(n_934),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1298),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1312),
.B(n_1094),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1311),
.B(n_914),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1314),
.B(n_881),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1310),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1320),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1322),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1296),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1323),
.Y(n_1371)
);

OAI21xp33_ASAP7_75t_L g1372 ( 
.A1(n_1300),
.A2(n_1317),
.B(n_1316),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1332),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1346),
.B(n_959),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1304),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1292),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1333),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1340),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1325),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1324),
.B(n_991),
.Y(n_1380)
);

INVx4_ASAP7_75t_SL g1381 ( 
.A(n_1327),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1342),
.Y(n_1382)
);

AO22x2_ASAP7_75t_L g1383 ( 
.A1(n_1308),
.A2(n_1005),
.B1(n_1132),
.B2(n_1069),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1344),
.B(n_1151),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1347),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1329),
.B(n_978),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1334),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1335),
.B(n_1179),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1348),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1331),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1343),
.B(n_847),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1289),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1336),
.B(n_1006),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1303),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1341),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1337),
.B(n_1158),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1338),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1289),
.Y(n_1398)
);

NAND3x1_ASAP7_75t_L g1399 ( 
.A(n_1307),
.B(n_1295),
.C(n_1345),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1349),
.B(n_1077),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1315),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1351),
.B(n_1172),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1289),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1326),
.B(n_1239),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1313),
.Y(n_1405)
);

NAND2x1_ASAP7_75t_L g1406 ( 
.A(n_1350),
.B(n_882),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1328),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1352),
.B(n_1240),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1291),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1328),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1294),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1305),
.B(n_969),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1306),
.B(n_998),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1318),
.B(n_1180),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1319),
.B(n_1033),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1330),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1301),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1301),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1321),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1301),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1339),
.B(n_1181),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1310),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1299),
.B(n_1184),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1302),
.B(n_1071),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1312),
.B(n_1137),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1312),
.B(n_1137),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1339),
.B(n_980),
.Y(n_1428)
);

INVx4_ASAP7_75t_L g1429 ( 
.A(n_1301),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1301),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1339),
.B(n_980),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1312),
.B(n_1153),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1339),
.B(n_980),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1312),
.B(n_1052),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1301),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1301),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1293),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1293),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1301),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1321),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1321),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1301),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1310),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1312),
.B(n_1176),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_1288),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1339),
.B(n_849),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1293),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1321),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1315),
.B(n_976),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1293),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1293),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1321),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1321),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1299),
.B(n_1166),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1302),
.B(n_1008),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1293),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1321),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1299),
.B(n_1170),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1293),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1312),
.B(n_1176),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1339),
.A2(n_927),
.B1(n_1049),
.B2(n_864),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1312),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1300),
.A2(n_852),
.B1(n_857),
.B2(n_854),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1299),
.B(n_858),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1355),
.Y(n_1466)
);

NOR3xp33_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1012),
.C(n_1010),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1359),
.Y(n_1468)
);

INVxp33_ASAP7_75t_L g1469 ( 
.A(n_1396),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1362),
.B(n_860),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1369),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1376),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1358),
.B(n_862),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1455),
.B(n_1015),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1378),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1459),
.B(n_1465),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1385),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1388),
.B(n_1016),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1353),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1390),
.B(n_1019),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1368),
.B(n_865),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1370),
.B(n_867),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1440),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1360),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1420),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1361),
.B(n_868),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1367),
.B(n_1028),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1446),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1404),
.B(n_1034),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1371),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1382),
.B(n_870),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1363),
.Y(n_1492)
);

O2A1O1Ixp5_ASAP7_75t_L g1493 ( 
.A1(n_1389),
.A2(n_1366),
.B(n_1442),
.C(n_1441),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1372),
.A2(n_1178),
.B1(n_916),
.B2(n_924),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1369),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1449),
.A2(n_875),
.B1(n_877),
.B2(n_876),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1453),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1375),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1463),
.B(n_878),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1454),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1458),
.Y(n_1501)
);

NAND2xp33_ASAP7_75t_L g1502 ( 
.A(n_1409),
.B(n_1399),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1464),
.A2(n_1056),
.B(n_1063),
.C(n_1039),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1397),
.A2(n_947),
.B(n_899),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1416),
.B(n_1428),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1431),
.B(n_1064),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1364),
.B(n_879),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1462),
.A2(n_981),
.B1(n_1013),
.B2(n_973),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1433),
.B(n_1070),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1417),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1384),
.B(n_1380),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1423),
.B(n_1076),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_SL g1514 ( 
.A1(n_1400),
.A2(n_887),
.B1(n_891),
.B2(n_885),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1426),
.B(n_1082),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1373),
.B(n_880),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1422),
.A2(n_1447),
.B(n_1365),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1393),
.B(n_1089),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1444),
.B(n_894),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1448),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1451),
.B(n_1095),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1452),
.B(n_1099),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1357),
.A2(n_903),
.B1(n_904),
.B2(n_897),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1377),
.B(n_907),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_L g1526 ( 
.A(n_1409),
.B(n_908),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1457),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1460),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1379),
.B(n_1113),
.Y(n_1529)
);

NAND2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1391),
.B(n_911),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1394),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1398),
.B(n_1118),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1398),
.B(n_1125),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1387),
.B(n_915),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_L g1535 ( 
.A(n_1403),
.B(n_917),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1395),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1386),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1403),
.B(n_1136),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1427),
.B(n_1139),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1356),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1392),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1410),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1445),
.B(n_918),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1461),
.B(n_1456),
.Y(n_1544)
);

NAND2xp33_ASAP7_75t_L g1545 ( 
.A(n_1402),
.B(n_922),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1407),
.Y(n_1546)
);

INVxp67_ASAP7_75t_SL g1547 ( 
.A(n_1401),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1443),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1408),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1406),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1434),
.B(n_1142),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1374),
.B(n_1157),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1450),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1354),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1418),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1421),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1432),
.B(n_1160),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1419),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1425),
.B(n_1167),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1430),
.B(n_1169),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1381),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1412),
.B(n_1171),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1429),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1435),
.B(n_932),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1413),
.B(n_1183),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1411),
.A2(n_1027),
.B1(n_1037),
.B2(n_1018),
.Y(n_1566)
);

NAND2x1p5_ASAP7_75t_L g1567 ( 
.A(n_1436),
.B(n_955),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1437),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1381),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1414),
.B(n_1415),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1405),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1450),
.B(n_1383),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1369),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1424),
.A2(n_937),
.B1(n_939),
.B2(n_935),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1355),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1355),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1389),
.A2(n_843),
.B(n_841),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1353),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1355),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1396),
.B(n_940),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1390),
.A2(n_1055),
.B(n_1038),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1358),
.B(n_942),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1358),
.B(n_945),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1424),
.A2(n_949),
.B1(n_953),
.B2(n_948),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1355),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1353),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1404),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1353),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1368),
.B(n_957),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_L g1590 ( 
.A(n_1382),
.B(n_958),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1355),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1396),
.B(n_960),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1355),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1358),
.B(n_964),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1368),
.B(n_970),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1353),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1358),
.B(n_979),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1358),
.B(n_984),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_L g1599 ( 
.A(n_1424),
.B(n_987),
.C(n_986),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1358),
.B(n_988),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1443),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1358),
.B(n_989),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1358),
.B(n_992),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1396),
.B(n_997),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1355),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1381),
.B(n_982),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1396),
.B(n_1002),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1358),
.B(n_1003),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1443),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1368),
.B(n_1011),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1358),
.B(n_1020),
.Y(n_1611)
);

AND2x6_ASAP7_75t_SL g1612 ( 
.A(n_1414),
.B(n_1093),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1358),
.B(n_1022),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1368),
.B(n_1024),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1404),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1358),
.B(n_1026),
.Y(n_1616)
);

AND2x6_ASAP7_75t_SL g1617 ( 
.A(n_1414),
.B(n_1105),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1358),
.B(n_1030),
.Y(n_1618)
);

OAI22x1_ASAP7_75t_R g1619 ( 
.A1(n_1382),
.A2(n_1174),
.B1(n_1164),
.B2(n_1036),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1465),
.A2(n_1127),
.B1(n_1131),
.B2(n_1123),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1396),
.B(n_1032),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1358),
.B(n_1040),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1358),
.B(n_1041),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1476),
.B(n_1044),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1469),
.B(n_1047),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1493),
.A2(n_1175),
.B(n_1163),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1479),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1473),
.B(n_1150),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1470),
.B(n_1154),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1580),
.B(n_1050),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1484),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

INVx4_ASAP7_75t_L g1633 ( 
.A(n_1490),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1466),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1474),
.A2(n_1182),
.B(n_1102),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1609),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1517),
.A2(n_890),
.B(n_851),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1512),
.B(n_1054),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1490),
.B(n_1059),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1553),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1581),
.A2(n_1504),
.B(n_1505),
.Y(n_1641)
);

AND2x2_ASAP7_75t_SL g1642 ( 
.A(n_1502),
.B(n_1075),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1587),
.B(n_1615),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1490),
.B(n_1031),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1468),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1480),
.A2(n_1098),
.B(n_1029),
.Y(n_1646)
);

BUFx8_ASAP7_75t_L g1647 ( 
.A(n_1571),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1620),
.A2(n_1583),
.B(n_1582),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1594),
.A2(n_1147),
.B(n_1112),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1592),
.B(n_1140),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1597),
.A2(n_1144),
.B(n_1143),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1604),
.B(n_1145),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1607),
.B(n_1060),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1598),
.A2(n_1155),
.B(n_1149),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1600),
.A2(n_1168),
.B(n_1161),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1483),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1514),
.B(n_1065),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1621),
.B(n_1068),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1599),
.A2(n_1072),
.B1(n_1078),
.B2(n_1073),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1568),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1602),
.B(n_1079),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1472),
.Y(n_1662)
);

NOR2xp67_ASAP7_75t_L g1663 ( 
.A(n_1488),
.B(n_1081),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1544),
.B(n_1483),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1475),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1603),
.A2(n_1126),
.B(n_1067),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1608),
.A2(n_1134),
.B(n_1128),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1611),
.A2(n_1177),
.B(n_1173),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1467),
.A2(n_965),
.B(n_1130),
.C(n_1085),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1613),
.A2(n_853),
.B(n_845),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1547),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1616),
.B(n_1156),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1618),
.A2(n_861),
.B(n_856),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1622),
.B(n_1083),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1492),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1623),
.A2(n_871),
.B(n_866),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1478),
.B(n_1116),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1577),
.A2(n_1120),
.B(n_886),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1515),
.B(n_1086),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1511),
.B(n_1087),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1537),
.A2(n_1485),
.B(n_1477),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1497),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1500),
.Y(n_1683)
);

AND2x6_ASAP7_75t_L g1684 ( 
.A(n_1561),
.B(n_882),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1501),
.A2(n_895),
.B(n_872),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1575),
.A2(n_1090),
.B1(n_1096),
.B2(n_1091),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1489),
.B(n_1576),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1498),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1543),
.B(n_1103),
.C(n_1097),
.Y(n_1689)
);

AOI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1506),
.A2(n_1035),
.B(n_882),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1579),
.A2(n_1104),
.B1(n_1108),
.B2(n_1106),
.Y(n_1691)
);

AOI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1509),
.A2(n_1035),
.B(n_1101),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1507),
.B(n_1111),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1585),
.A2(n_1115),
.B(n_929),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1591),
.A2(n_931),
.B(n_900),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1593),
.A2(n_1117),
.B1(n_1121),
.B2(n_1119),
.Y(n_1696)
);

A2O1A1Ixp33_ASAP7_75t_L g1697 ( 
.A1(n_1503),
.A2(n_1135),
.B(n_1122),
.C(n_1133),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1511),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1556),
.Y(n_1699)
);

AO21x1_ASAP7_75t_L g1700 ( 
.A1(n_1494),
.A2(n_1035),
.B(n_1077),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1605),
.B(n_1551),
.Y(n_1701)
);

CKINVDCx6p67_ASAP7_75t_R g1702 ( 
.A(n_1570),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1578),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1548),
.B(n_1075),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1518),
.A2(n_938),
.B(n_936),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1499),
.B(n_1519),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1508),
.A2(n_1124),
.B(n_1148),
.C(n_1138),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1520),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1556),
.Y(n_1709)
);

NOR2xp67_ASAP7_75t_L g1710 ( 
.A(n_1471),
.B(n_941),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1549),
.A2(n_1075),
.B1(n_1162),
.B2(n_1159),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1574),
.B(n_943),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1487),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1552),
.B(n_1159),
.Y(n_1714)
);

BUFx8_ASAP7_75t_L g1715 ( 
.A(n_1495),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1586),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1545),
.A2(n_1061),
.B(n_1051),
.Y(n_1717)
);

O2A1O1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1584),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1606),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1560),
.A2(n_1100),
.B(n_1088),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1566),
.A2(n_1162),
.B(n_1165),
.C(n_1159),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1540),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1612),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1516),
.A2(n_1110),
.B(n_951),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1525),
.A2(n_961),
.B(n_946),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1573),
.A2(n_1165),
.B1(n_1162),
.B2(n_1023),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1481),
.A2(n_985),
.B(n_974),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1524),
.B(n_993),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1588),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1590),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1530),
.A2(n_1165),
.B(n_1004),
.C(n_967),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1596),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1510),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1539),
.B(n_1513),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1521),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1589),
.A2(n_1048),
.B(n_1046),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1557),
.B(n_962),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1527),
.B(n_4),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1528),
.B(n_5),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1627),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1631),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1636),
.B(n_1569),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1713),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1699),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1641),
.A2(n_1542),
.B(n_1595),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1634),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1648),
.A2(n_1614),
.B(n_1610),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1706),
.B(n_1617),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1734),
.B(n_1559),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_SL g1750 ( 
.A(n_1624),
.B(n_1486),
.C(n_1491),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1635),
.A2(n_1534),
.B(n_1535),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1681),
.A2(n_1564),
.B(n_1523),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1645),
.Y(n_1753)
);

O2A1O1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1630),
.A2(n_1526),
.B(n_1482),
.C(n_1496),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1653),
.B(n_1572),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1660),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1658),
.B(n_1554),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1699),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1642),
.B(n_1541),
.Y(n_1759)
);

O2A1O1Ixp5_ASAP7_75t_L g1760 ( 
.A1(n_1712),
.A2(n_1533),
.B(n_1538),
.C(n_1532),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1656),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1640),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1675),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_SL g1764 ( 
.A(n_1719),
.B(n_1563),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1638),
.B(n_1562),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1688),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1656),
.Y(n_1767)
);

O2A1O1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1628),
.A2(n_1565),
.B(n_1555),
.C(n_1558),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1701),
.A2(n_1522),
.B(n_1546),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1632),
.Y(n_1770)
);

BUFx8_ASAP7_75t_L g1771 ( 
.A(n_1656),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1703),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_R g1773 ( 
.A(n_1647),
.B(n_1536),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1687),
.B(n_1531),
.Y(n_1774)
);

AOI222xp33_ASAP7_75t_L g1775 ( 
.A1(n_1723),
.A2(n_1619),
.B1(n_1529),
.B2(n_1550),
.C1(n_1000),
.C2(n_995),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1650),
.B(n_1567),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1652),
.A2(n_1101),
.B(n_996),
.Y(n_1777)
);

AOI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1693),
.A2(n_1084),
.B1(n_1014),
.B2(n_971),
.C(n_1101),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1716),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1629),
.A2(n_676),
.B(n_674),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1737),
.A2(n_5),
.B(n_6),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1671),
.B(n_1035),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1643),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1689),
.B(n_6),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1661),
.A2(n_678),
.B(n_677),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1679),
.B(n_7),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1722),
.B(n_1035),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1708),
.B(n_7),
.Y(n_1788)
);

INVx6_ASAP7_75t_L g1789 ( 
.A(n_1715),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1698),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1633),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1672),
.A2(n_681),
.B(n_680),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_R g1793 ( 
.A(n_1709),
.B(n_682),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1662),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1729),
.Y(n_1795)
);

CKINVDCx8_ASAP7_75t_R g1796 ( 
.A(n_1644),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1697),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1702),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1677),
.B(n_8),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1674),
.A2(n_1637),
.B(n_1626),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1651),
.A2(n_684),
.B(n_683),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1665),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1644),
.B(n_685),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1682),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1683),
.B(n_9),
.Y(n_1805)
);

O2A1O1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1669),
.A2(n_13),
.B(n_10),
.C(n_12),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1654),
.A2(n_689),
.B(n_688),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1733),
.Y(n_1808)
);

O2A1O1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1718),
.A2(n_15),
.B(n_12),
.C(n_14),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1730),
.A2(n_18),
.B(n_19),
.C(n_17),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1659),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1655),
.A2(n_692),
.B(n_690),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1732),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1664),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1735),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1667),
.A2(n_695),
.B(n_694),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1738),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1668),
.A2(n_698),
.B(n_696),
.Y(n_1818)
);

NAND2x1p5_ASAP7_75t_L g1819 ( 
.A(n_1704),
.B(n_1639),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1666),
.B(n_16),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1649),
.A2(n_22),
.B(n_23),
.C(n_21),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1707),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1646),
.A2(n_1705),
.B(n_1673),
.C(n_1676),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1657),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1824)
);

INVxp67_ASAP7_75t_SL g1825 ( 
.A(n_1739),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1684),
.Y(n_1826)
);

BUFx8_ASAP7_75t_L g1827 ( 
.A(n_1684),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1684),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1714),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1690),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1686),
.B(n_25),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1670),
.A2(n_1720),
.B(n_1731),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1691),
.B(n_26),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1692),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1726),
.Y(n_1835)
);

INVx6_ASAP7_75t_L g1836 ( 
.A(n_1663),
.Y(n_1836)
);

INVx6_ASAP7_75t_L g1837 ( 
.A(n_1710),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1721),
.A2(n_1685),
.B(n_1695),
.C(n_1694),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1680),
.Y(n_1839)
);

AOI21x1_ASAP7_75t_L g1840 ( 
.A1(n_1700),
.A2(n_1678),
.B(n_1717),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1625),
.A2(n_1696),
.B1(n_1728),
.B2(n_1727),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1736),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1725),
.A2(n_700),
.B(n_699),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1711),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1724),
.A2(n_703),
.B(n_701),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1641),
.A2(n_705),
.B(n_704),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1706),
.B(n_27),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1641),
.A2(n_708),
.B(n_707),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1634),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_SL g1850 ( 
.A(n_1642),
.B(n_709),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1706),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1851)
);

NAND2xp33_ASAP7_75t_SL g1852 ( 
.A(n_1650),
.B(n_29),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1627),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1627),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1706),
.B(n_30),
.Y(n_1855)
);

AND2x6_ASAP7_75t_L g1856 ( 
.A(n_1708),
.B(n_711),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1734),
.B(n_30),
.Y(n_1857)
);

O2A1O1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1706),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1734),
.B(n_33),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1734),
.B(n_34),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1634),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1706),
.B(n_34),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1636),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1634),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1636),
.B(n_713),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1706),
.B(n_35),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1749),
.B(n_35),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1815),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1855),
.B(n_36),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1859),
.B(n_36),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1862),
.A2(n_37),
.B(n_38),
.Y(n_1871)
);

AO31x2_ASAP7_75t_L g1872 ( 
.A1(n_1830),
.A2(n_715),
.A3(n_716),
.B(n_714),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1866),
.B(n_38),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1783),
.B(n_39),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1746),
.Y(n_1875)
);

AO32x2_ASAP7_75t_L g1876 ( 
.A1(n_1822),
.A2(n_42),
.A3(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1800),
.A2(n_718),
.B(n_717),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1758),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1834),
.A2(n_721),
.B(n_719),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1863),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1748),
.A2(n_1860),
.B1(n_1857),
.B2(n_1781),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1850),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1805),
.B(n_45),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1846),
.A2(n_45),
.B(n_46),
.Y(n_1884)
);

O2A1O1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1847),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1848),
.A2(n_723),
.B(n_722),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1743),
.B(n_47),
.Y(n_1887)
);

AO21x1_ASAP7_75t_L g1888 ( 
.A1(n_1820),
.A2(n_1852),
.B(n_1747),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1768),
.A2(n_50),
.B(n_51),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1762),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1863),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1786),
.B(n_51),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1745),
.A2(n_52),
.B(n_53),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1774),
.B(n_53),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1771),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1757),
.B(n_1756),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1740),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1840),
.A2(n_725),
.B(n_724),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1758),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1832),
.A2(n_727),
.B(n_726),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1753),
.Y(n_1901)
);

NAND3xp33_ASAP7_75t_L g1902 ( 
.A(n_1851),
.B(n_54),
.C(n_55),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1858),
.B(n_54),
.C(n_55),
.Y(n_1903)
);

OA21x2_ASAP7_75t_L g1904 ( 
.A1(n_1760),
.A2(n_56),
.B(n_57),
.Y(n_1904)
);

OAI21x1_ASAP7_75t_L g1905 ( 
.A1(n_1801),
.A2(n_729),
.B(n_728),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_L g1906 ( 
.A(n_1784),
.B(n_56),
.C(n_58),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1752),
.A2(n_58),
.B(n_59),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1765),
.B(n_59),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1755),
.B(n_60),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1823),
.A2(n_60),
.B(n_61),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1790),
.B(n_62),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1761),
.Y(n_1912)
);

NAND2xp33_ASAP7_75t_L g1913 ( 
.A(n_1750),
.B(n_62),
.Y(n_1913)
);

BUFx10_ASAP7_75t_L g1914 ( 
.A(n_1789),
.Y(n_1914)
);

OAI21x1_ASAP7_75t_L g1915 ( 
.A1(n_1807),
.A2(n_732),
.B(n_731),
.Y(n_1915)
);

OAI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1754),
.A2(n_63),
.B(n_64),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1796),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1833),
.B(n_63),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1761),
.Y(n_1919)
);

BUFx10_ASAP7_75t_L g1920 ( 
.A(n_1789),
.Y(n_1920)
);

NAND2x1p5_ASAP7_75t_L g1921 ( 
.A(n_1798),
.B(n_733),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1776),
.B(n_64),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1831),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_L g1924 ( 
.A1(n_1812),
.A2(n_735),
.B(n_734),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1794),
.Y(n_1925)
);

AO31x2_ASAP7_75t_L g1926 ( 
.A1(n_1829),
.A2(n_738),
.A3(n_740),
.B(n_736),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1825),
.B(n_65),
.Y(n_1927)
);

AO22x2_ASAP7_75t_L g1928 ( 
.A1(n_1817),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1769),
.A2(n_742),
.B(n_741),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1799),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1770),
.B(n_70),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1759),
.A2(n_1838),
.B(n_1782),
.Y(n_1932)
);

AO31x2_ASAP7_75t_L g1933 ( 
.A1(n_1808),
.A2(n_1810),
.A3(n_1763),
.B(n_1766),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1741),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1802),
.B(n_72),
.Y(n_1935)
);

AO32x2_ASAP7_75t_L g1936 ( 
.A1(n_1814),
.A2(n_74),
.A3(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_1936)
);

NAND2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1744),
.B(n_743),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1839),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1816),
.A2(n_745),
.B(n_744),
.Y(n_1939)
);

BUFx12f_ASAP7_75t_L g1940 ( 
.A(n_1827),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1751),
.A2(n_73),
.B(n_74),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1809),
.A2(n_75),
.B(n_77),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1797),
.A2(n_78),
.B(n_79),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1806),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_1944)
);

OA21x2_ASAP7_75t_L g1945 ( 
.A1(n_1785),
.A2(n_80),
.B(n_81),
.Y(n_1945)
);

AO22x2_ASAP7_75t_L g1946 ( 
.A1(n_1804),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_1946)
);

OAI21x1_ASAP7_75t_L g1947 ( 
.A1(n_1898),
.A2(n_1780),
.B(n_1843),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1875),
.Y(n_1948)
);

OAI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1869),
.A2(n_1873),
.B1(n_1871),
.B2(n_1881),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1880),
.Y(n_1950)
);

OAI21x1_ASAP7_75t_L g1951 ( 
.A1(n_1900),
.A2(n_1845),
.B(n_1818),
.Y(n_1951)
);

AO21x2_ASAP7_75t_L g1952 ( 
.A1(n_1910),
.A2(n_1777),
.B(n_1792),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1901),
.Y(n_1953)
);

O2A1O1Ixp5_ASAP7_75t_L g1954 ( 
.A1(n_1916),
.A2(n_1942),
.B(n_1882),
.C(n_1888),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1877),
.A2(n_1861),
.B(n_1849),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1940),
.Y(n_1956)
);

AO21x2_ASAP7_75t_L g1957 ( 
.A1(n_1932),
.A2(n_1787),
.B(n_1864),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1880),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1925),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1868),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1879),
.A2(n_1842),
.B(n_1819),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1897),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1886),
.A2(n_1788),
.B(n_1841),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1896),
.B(n_1836),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1891),
.B(n_1890),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1870),
.B(n_1835),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1913),
.A2(n_1844),
.B1(n_1837),
.B2(n_1775),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1934),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1878),
.B(n_1836),
.Y(n_1969)
);

OAI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1902),
.A2(n_1811),
.B(n_1821),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1884),
.A2(n_1828),
.B(n_1826),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_SL g1972 ( 
.A1(n_1935),
.A2(n_1824),
.B(n_1778),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1899),
.Y(n_1973)
);

AND2x4_ASAP7_75t_SL g1974 ( 
.A(n_1914),
.B(n_1865),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1895),
.B(n_1767),
.Y(n_1975)
);

NOR2xp67_ASAP7_75t_L g1976 ( 
.A(n_1927),
.B(n_1791),
.Y(n_1976)
);

CKINVDCx6p67_ASAP7_75t_R g1977 ( 
.A(n_1920),
.Y(n_1977)
);

OAI21x1_ASAP7_75t_L g1978 ( 
.A1(n_1905),
.A2(n_1779),
.B(n_1772),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1894),
.B(n_1795),
.Y(n_1979)
);

OA21x2_ASAP7_75t_L g1980 ( 
.A1(n_1907),
.A2(n_1853),
.B(n_1813),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1903),
.A2(n_1856),
.B(n_1803),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1867),
.B(n_1854),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1933),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1912),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1938),
.Y(n_1985)
);

AO21x2_ASAP7_75t_L g1986 ( 
.A1(n_1929),
.A2(n_1793),
.B(n_1773),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1893),
.A2(n_1764),
.B(n_1856),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1941),
.A2(n_1856),
.B(n_1742),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1889),
.A2(n_1837),
.B(n_85),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1933),
.Y(n_1990)
);

CKINVDCx6p67_ASAP7_75t_R g1991 ( 
.A(n_1911),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1874),
.Y(n_1992)
);

OAI22x1_ASAP7_75t_L g1993 ( 
.A1(n_1918),
.A2(n_1906),
.B1(n_1883),
.B2(n_1922),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1944),
.A2(n_82),
.B(n_84),
.Y(n_1994)
);

OAI21x1_ASAP7_75t_L g1995 ( 
.A1(n_1963),
.A2(n_1939),
.B(n_1924),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1960),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1948),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1965),
.Y(n_1998)
);

OAI21x1_ASAP7_75t_SL g1999 ( 
.A1(n_1981),
.A2(n_1885),
.B(n_1923),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1977),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1992),
.B(n_1931),
.Y(n_2001)
);

A2O1A1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1989),
.A2(n_1909),
.B(n_1908),
.C(n_1930),
.Y(n_2002)
);

BUFx12f_ASAP7_75t_L g2003 ( 
.A(n_1956),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_SL g2004 ( 
.A(n_1975),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_L g2005 ( 
.A1(n_1951),
.A2(n_1915),
.B(n_1904),
.Y(n_2005)
);

NAND2x1p5_ASAP7_75t_L g2006 ( 
.A(n_1950),
.B(n_1917),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1962),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1985),
.B(n_1912),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1987),
.A2(n_1954),
.B(n_1949),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1953),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1959),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1968),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1983),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1979),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1955),
.Y(n_2015)
);

INVx4_ASAP7_75t_L g2016 ( 
.A(n_1950),
.Y(n_2016)
);

OA21x2_ASAP7_75t_L g2017 ( 
.A1(n_1990),
.A2(n_1887),
.B(n_1892),
.Y(n_2017)
);

NAND2x1p5_ASAP7_75t_L g2018 ( 
.A(n_1984),
.B(n_1919),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1966),
.B(n_1928),
.Y(n_2019)
);

AND2x4_ASAP7_75t_L g2020 ( 
.A(n_1976),
.B(n_1926),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1982),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1967),
.A2(n_1946),
.B1(n_1921),
.B2(n_1945),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1957),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1973),
.B(n_85),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1958),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1978),
.Y(n_2026)
);

BUFx4f_ASAP7_75t_L g2027 ( 
.A(n_1991),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1980),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1980),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1961),
.Y(n_2030)
);

OAI21x1_ASAP7_75t_L g2031 ( 
.A1(n_1947),
.A2(n_1937),
.B(n_1943),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1993),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1970),
.A2(n_1936),
.B(n_1876),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1964),
.B(n_1971),
.Y(n_2034)
);

AOI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1952),
.A2(n_1936),
.B(n_1876),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1988),
.A2(n_1872),
.B(n_1926),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1974),
.B(n_1872),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1994),
.Y(n_2038)
);

AOI21xp33_ASAP7_75t_L g2039 ( 
.A1(n_1986),
.A2(n_86),
.B(n_87),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1994),
.A2(n_87),
.B(n_88),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_1969),
.B(n_88),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1972),
.Y(n_2042)
);

OAI21x1_ASAP7_75t_L g2043 ( 
.A1(n_1963),
.A2(n_748),
.B(n_746),
.Y(n_2043)
);

NAND2x1_ASAP7_75t_L g2044 ( 
.A(n_1948),
.B(n_89),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1966),
.B(n_89),
.Y(n_2045)
);

INVxp67_ASAP7_75t_L g2046 ( 
.A(n_2034),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1997),
.B(n_2010),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2011),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2014),
.B(n_91),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1996),
.Y(n_2050)
);

BUFx2_ASAP7_75t_L g2051 ( 
.A(n_2032),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2012),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_2017),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_2036),
.A2(n_92),
.B(n_93),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_2017),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2007),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2021),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_2013),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_2042),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2029),
.Y(n_2060)
);

NAND2x1_ASAP7_75t_L g2061 ( 
.A(n_2038),
.B(n_2015),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2023),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2001),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_SL g2064 ( 
.A1(n_2033),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_L g2065 ( 
.A(n_2027),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2008),
.B(n_94),
.Y(n_2066)
);

INVx8_ASAP7_75t_L g2067 ( 
.A(n_2003),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2028),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_2005),
.A2(n_1995),
.B(n_2031),
.Y(n_2069)
);

BUFx4f_ASAP7_75t_SL g2070 ( 
.A(n_2000),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1998),
.B(n_96),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2030),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2019),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2045),
.B(n_97),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_2026),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2020),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_2025),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2024),
.B(n_97),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2037),
.Y(n_2079)
);

AOI21x1_ASAP7_75t_L g2080 ( 
.A1(n_2009),
.A2(n_98),
.B(n_99),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2044),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2044),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2018),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2043),
.Y(n_2084)
);

OAI222xp33_ASAP7_75t_L g2085 ( 
.A1(n_2022),
.A2(n_101),
.B1(n_104),
.B2(n_99),
.C1(n_100),
.C2(n_102),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_2035),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2041),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2016),
.B(n_101),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2006),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1999),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_2004),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2040),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_2002),
.B(n_102),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1999),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2039),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1997),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1997),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1997),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1997),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1996),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1996),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1997),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1996),
.Y(n_2103)
);

OAI21x1_ASAP7_75t_L g2104 ( 
.A1(n_2036),
.A2(n_104),
.B(n_105),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1997),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1998),
.B(n_105),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1996),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1998),
.B(n_106),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1996),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1997),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1997),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_2032),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_2032),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1998),
.B(n_106),
.Y(n_2114)
);

AO21x2_ASAP7_75t_L g2115 ( 
.A1(n_2023),
.A2(n_107),
.B(n_108),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2034),
.B(n_108),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1996),
.Y(n_2117)
);

INVx2_ASAP7_75t_SL g2118 ( 
.A(n_1998),
.Y(n_2118)
);

OA21x2_ASAP7_75t_L g2119 ( 
.A1(n_2035),
.A2(n_109),
.B(n_110),
.Y(n_2119)
);

AO21x2_ASAP7_75t_L g2120 ( 
.A1(n_2023),
.A2(n_110),
.B(n_111),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_2003),
.Y(n_2121)
);

OAI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_2095),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.C(n_114),
.Y(n_2122)
);

AO21x2_ASAP7_75t_L g2123 ( 
.A1(n_2062),
.A2(n_114),
.B(n_115),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_SL g2124 ( 
.A1(n_2121),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_2124)
);

AOI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_2086),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2073),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2047),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2093),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_124),
.Y(n_2128)
);

OAI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_2092),
.A2(n_126),
.B1(n_123),
.B2(n_125),
.Y(n_2129)
);

AOI21xp5_ASAP7_75t_L g2130 ( 
.A1(n_2116),
.A2(n_125),
.B(n_126),
.Y(n_2130)
);

OAI21x1_ASAP7_75t_L g2131 ( 
.A1(n_2061),
.A2(n_127),
.B(n_128),
.Y(n_2131)
);

AOI211xp5_ASAP7_75t_L g2132 ( 
.A1(n_2085),
.A2(n_137),
.B(n_145),
.C(n_127),
.Y(n_2132)
);

AOI21xp33_ASAP7_75t_L g2133 ( 
.A1(n_2090),
.A2(n_2094),
.B(n_2119),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2048),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2046),
.B(n_129),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2068),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_2061),
.A2(n_129),
.B(n_130),
.Y(n_2137)
);

OAI211xp5_ASAP7_75t_L g2138 ( 
.A1(n_2064),
.A2(n_133),
.B(n_130),
.C(n_131),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2060),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2119),
.A2(n_134),
.B1(n_131),
.B2(n_133),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2096),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2118),
.B(n_134),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2097),
.Y(n_2143)
);

AOI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2112),
.A2(n_2113),
.B1(n_2051),
.B2(n_2087),
.C(n_2063),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2059),
.B(n_135),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_2091),
.Y(n_2146)
);

OAI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_2051),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_2147)
);

AOI21xp33_ASAP7_75t_L g2148 ( 
.A1(n_2082),
.A2(n_136),
.B(n_138),
.Y(n_2148)
);

OAI33xp33_ASAP7_75t_L g2149 ( 
.A1(n_2049),
.A2(n_140),
.A3(n_142),
.B1(n_138),
.B2(n_139),
.B3(n_141),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_2115),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_2091),
.Y(n_2151)
);

OA21x2_ASAP7_75t_L g2152 ( 
.A1(n_2053),
.A2(n_143),
.B(n_145),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2077),
.B(n_146),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2083),
.B(n_146),
.Y(n_2154)
);

A2O1A1Ixp33_ASAP7_75t_L g2155 ( 
.A1(n_2054),
.A2(n_155),
.B(n_164),
.C(n_147),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2081),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2098),
.B(n_148),
.Y(n_2157)
);

AOI221xp5_ASAP7_75t_L g2158 ( 
.A1(n_2120),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.C(n_153),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2076),
.A2(n_2108),
.B1(n_2079),
.B2(n_2089),
.Y(n_2159)
);

AOI221xp5_ASAP7_75t_L g2160 ( 
.A1(n_2055),
.A2(n_2052),
.B1(n_2078),
.B2(n_2072),
.C(n_2111),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2108),
.A2(n_153),
.B1(n_150),
.B2(n_152),
.Y(n_2161)
);

AOI22xp33_ASAP7_75t_SL g2162 ( 
.A1(n_2104),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2162)
);

OAI211xp5_ASAP7_75t_L g2163 ( 
.A1(n_2080),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_2067),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2057),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_2165)
);

OAI211xp5_ASAP7_75t_SL g2166 ( 
.A1(n_2066),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2099),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2058),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2084),
.A2(n_160),
.B(n_161),
.Y(n_2169)
);

BUFx3_ASAP7_75t_L g2170 ( 
.A(n_2067),
.Y(n_2170)
);

OAI21x1_ASAP7_75t_L g2171 ( 
.A1(n_2069),
.A2(n_163),
.B(n_164),
.Y(n_2171)
);

AOI222xp33_ASAP7_75t_L g2172 ( 
.A1(n_2074),
.A2(n_166),
.B1(n_168),
.B2(n_163),
.C1(n_165),
.C2(n_167),
.Y(n_2172)
);

AOI222xp33_ASAP7_75t_L g2173 ( 
.A1(n_2071),
.A2(n_170),
.B1(n_172),
.B2(n_166),
.C1(n_169),
.C2(n_171),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_2106),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2102),
.B(n_172),
.Y(n_2175)
);

BUFx4f_ASAP7_75t_SL g2176 ( 
.A(n_2065),
.Y(n_2176)
);

A2O1A1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_2114),
.A2(n_182),
.B(n_190),
.C(n_173),
.Y(n_2177)
);

OAI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_2080),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2105),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_2091),
.B(n_174),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_2056),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2181)
);

AOI221xp5_ASAP7_75t_L g2182 ( 
.A1(n_2110),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.C(n_180),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2050),
.A2(n_2100),
.B1(n_2103),
.B2(n_2101),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2107),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2109),
.Y(n_2185)
);

OAI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2117),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_2186)
);

INVx8_ASAP7_75t_L g2187 ( 
.A(n_2065),
.Y(n_2187)
);

AOI221xp5_ASAP7_75t_L g2188 ( 
.A1(n_2075),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.C(n_187),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2088),
.B(n_185),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2070),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2093),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2070),
.B(n_191),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2059),
.B(n_192),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2068),
.Y(n_2194)
);

CKINVDCx11_ASAP7_75t_R g2195 ( 
.A(n_2121),
.Y(n_2195)
);

OAI211xp5_ASAP7_75t_L g2196 ( 
.A1(n_2093),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_2196)
);

OAI211xp5_ASAP7_75t_SL g2197 ( 
.A1(n_2094),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2046),
.B(n_195),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2047),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_2118),
.B(n_196),
.Y(n_2200)
);

AOI22xp33_ASAP7_75t_L g2201 ( 
.A1(n_2086),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_2201)
);

INVx3_ASAP7_75t_L g2202 ( 
.A(n_2091),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2086),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_2203)
);

AOI22xp33_ASAP7_75t_L g2204 ( 
.A1(n_2086),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2204)
);

AOI221xp5_ASAP7_75t_L g2205 ( 
.A1(n_2086),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.C(n_205),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_2061),
.A2(n_202),
.B(n_203),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2046),
.B(n_204),
.Y(n_2207)
);

AOI211xp5_ASAP7_75t_L g2208 ( 
.A1(n_2093),
.A2(n_214),
.B(n_222),
.C(n_206),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_2094),
.B(n_206),
.C(n_207),
.Y(n_2209)
);

OA21x2_ASAP7_75t_L g2210 ( 
.A1(n_2062),
.A2(n_207),
.B(n_208),
.Y(n_2210)
);

OAI211xp5_ASAP7_75t_L g2211 ( 
.A1(n_2093),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_2211)
);

AOI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_2086),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2086),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_2213)
);

OAI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2093),
.A2(n_212),
.B(n_213),
.Y(n_2214)
);

OAI211xp5_ASAP7_75t_L g2215 ( 
.A1(n_2093),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2086),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2046),
.B(n_219),
.Y(n_2217)
);

OAI21xp5_ASAP7_75t_SL g2218 ( 
.A1(n_2093),
.A2(n_219),
.B(n_220),
.Y(n_2218)
);

AOI22xp33_ASAP7_75t_L g2219 ( 
.A1(n_2086),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2127),
.B(n_221),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2199),
.B(n_223),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_2152),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2134),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2160),
.B(n_223),
.Y(n_2224)
);

NOR2x1_ASAP7_75t_L g2225 ( 
.A(n_2146),
.B(n_224),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2151),
.B(n_224),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2141),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_L g2228 ( 
.A(n_2195),
.B(n_225),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2135),
.B(n_225),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2149),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2202),
.B(n_226),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2152),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2143),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2167),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2144),
.B(n_228),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2179),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2218),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2139),
.Y(n_2238)
);

AOI222xp33_ASAP7_75t_L g2239 ( 
.A1(n_2214),
.A2(n_231),
.B1(n_233),
.B2(n_229),
.C1(n_230),
.C2(n_232),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2207),
.B(n_232),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2145),
.B(n_233),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2136),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2194),
.Y(n_2243)
);

AND2x4_ASAP7_75t_SL g2244 ( 
.A(n_2142),
.B(n_234),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2193),
.B(n_235),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2198),
.B(n_235),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2157),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2175),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2170),
.B(n_236),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2185),
.Y(n_2250)
);

INVx2_ASAP7_75t_SL g2251 ( 
.A(n_2187),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2133),
.B(n_2189),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2210),
.B(n_237),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2210),
.Y(n_2254)
);

BUFx3_ASAP7_75t_L g2255 ( 
.A(n_2176),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2159),
.Y(n_2256)
);

OAI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2191),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2257)
);

BUFx3_ASAP7_75t_L g2258 ( 
.A(n_2187),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_2200),
.B(n_239),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2168),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2123),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_2154),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2140),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2153),
.B(n_243),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2131),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2183),
.B(n_243),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2164),
.B(n_244),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2217),
.B(n_245),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2171),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2130),
.B(n_245),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2192),
.B(n_246),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2137),
.B(n_2206),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2174),
.B(n_2180),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2161),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2209),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2178),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2125),
.B(n_247),
.Y(n_2277)
);

BUFx3_ASAP7_75t_L g2278 ( 
.A(n_2124),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2201),
.B(n_248),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2147),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2163),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2205),
.B(n_249),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_2156),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2129),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2122),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2177),
.B(n_250),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2169),
.B(n_250),
.Y(n_2287)
);

NAND2x1p5_ASAP7_75t_SL g2288 ( 
.A(n_2208),
.B(n_2166),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2203),
.B(n_251),
.Y(n_2289)
);

HB1xp67_ASAP7_75t_L g2290 ( 
.A(n_2155),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2158),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2186),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2126),
.B(n_252),
.Y(n_2293)
);

BUFx6f_ASAP7_75t_L g2294 ( 
.A(n_2196),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2204),
.Y(n_2295)
);

AOI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_2211),
.A2(n_256),
.B1(n_253),
.B2(n_254),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_2215),
.Y(n_2297)
);

AND2x4_ASAP7_75t_SL g2298 ( 
.A(n_2219),
.B(n_254),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2212),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2213),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2148),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2216),
.Y(n_2302)
);

INVxp67_ASAP7_75t_SL g2303 ( 
.A(n_2150),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2165),
.B(n_256),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2162),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2188),
.B(n_257),
.Y(n_2306)
);

AOI21xp33_ASAP7_75t_SL g2307 ( 
.A1(n_2172),
.A2(n_257),
.B(n_258),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2190),
.B(n_258),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2197),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2173),
.B(n_259),
.Y(n_2310)
);

HB1xp67_ASAP7_75t_L g2311 ( 
.A(n_2182),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2181),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2128),
.B(n_259),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2184),
.B(n_260),
.Y(n_2314)
);

INVx1_ASAP7_75t_SL g2315 ( 
.A(n_2132),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2138),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2139),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2127),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2127),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_2152),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2127),
.B(n_261),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2127),
.B(n_261),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2127),
.Y(n_2323)
);

NOR2x1_ASAP7_75t_L g2324 ( 
.A(n_2146),
.B(n_262),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2127),
.B(n_262),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2127),
.B(n_263),
.Y(n_2326)
);

AND2x4_ASAP7_75t_L g2327 ( 
.A(n_2146),
.B(n_263),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_SL g2328 ( 
.A(n_2145),
.B(n_264),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2195),
.B(n_264),
.Y(n_2329)
);

BUFx2_ASAP7_75t_L g2330 ( 
.A(n_2152),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2127),
.B(n_265),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2127),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2127),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2195),
.B(n_265),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2127),
.B(n_266),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2127),
.Y(n_2336)
);

OAI222xp33_ASAP7_75t_L g2337 ( 
.A1(n_2159),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.C1(n_268),
.C2(n_270),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2139),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2290),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_2232),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2222),
.B(n_2330),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_2222),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2252),
.B(n_266),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2269),
.B(n_271),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2262),
.B(n_272),
.Y(n_2345)
);

INVx1_ASAP7_75t_SL g2346 ( 
.A(n_2255),
.Y(n_2346)
);

AOI22xp33_ASAP7_75t_SL g2347 ( 
.A1(n_2330),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2254),
.B(n_273),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2276),
.B(n_274),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2247),
.B(n_277),
.Y(n_2350)
);

INVxp67_ASAP7_75t_SL g2351 ( 
.A(n_2320),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2248),
.B(n_278),
.Y(n_2352)
);

AND2x4_ASAP7_75t_SL g2353 ( 
.A(n_2259),
.B(n_279),
.Y(n_2353)
);

INVx1_ASAP7_75t_SL g2354 ( 
.A(n_2258),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2280),
.B(n_279),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2223),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2318),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2319),
.B(n_280),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2227),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2323),
.B(n_280),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2332),
.B(n_281),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2272),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2333),
.B(n_281),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_2336),
.B(n_282),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2265),
.B(n_282),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2253),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2311),
.A2(n_283),
.B(n_284),
.Y(n_2367)
);

INVx1_ASAP7_75t_SL g2368 ( 
.A(n_2244),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_2233),
.B(n_283),
.Y(n_2369)
);

OR2x2_ASAP7_75t_L g2370 ( 
.A(n_2234),
.B(n_285),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2238),
.Y(n_2371)
);

OR2x2_ASAP7_75t_L g2372 ( 
.A(n_2236),
.B(n_2220),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2261),
.B(n_286),
.Y(n_2373)
);

HB1xp67_ASAP7_75t_L g2374 ( 
.A(n_2284),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2275),
.B(n_286),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2250),
.Y(n_2376)
);

NAND2x1p5_ASAP7_75t_L g2377 ( 
.A(n_2225),
.B(n_287),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2292),
.Y(n_2378)
);

OR2x2_ASAP7_75t_L g2379 ( 
.A(n_2326),
.B(n_288),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2260),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2221),
.B(n_288),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2322),
.B(n_289),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2325),
.B(n_289),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2321),
.B(n_290),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2317),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2331),
.B(n_290),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2335),
.B(n_291),
.Y(n_2387)
);

OAI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2237),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2235),
.B(n_292),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2241),
.B(n_293),
.Y(n_2390)
);

CKINVDCx16_ASAP7_75t_R g2391 ( 
.A(n_2278),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2281),
.B(n_294),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2251),
.B(n_294),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2301),
.B(n_295),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2266),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2327),
.B(n_2226),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2338),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2224),
.B(n_296),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2231),
.B(n_296),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2243),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2273),
.B(n_297),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2264),
.B(n_297),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2271),
.B(n_298),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2249),
.B(n_298),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2245),
.B(n_299),
.Y(n_2405)
);

INVx4_ASAP7_75t_L g2406 ( 
.A(n_2268),
.Y(n_2406)
);

AND2x4_ASAP7_75t_SL g2407 ( 
.A(n_2228),
.B(n_299),
.Y(n_2407)
);

NAND2x1_ASAP7_75t_L g2408 ( 
.A(n_2324),
.B(n_300),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2283),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2295),
.B(n_301),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2242),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2299),
.B(n_302),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2246),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2256),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2300),
.B(n_303),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2302),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2274),
.B(n_2303),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2312),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2309),
.B(n_304),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_L g2420 ( 
.A(n_2294),
.B(n_304),
.C(n_305),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2305),
.Y(n_2421)
);

OR2x2_ASAP7_75t_L g2422 ( 
.A(n_2288),
.B(n_306),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2287),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2286),
.B(n_2316),
.Y(n_2424)
);

AND2x4_ASAP7_75t_SL g2425 ( 
.A(n_2329),
.B(n_306),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2334),
.B(n_2229),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2294),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2240),
.B(n_307),
.Y(n_2428)
);

INVxp67_ASAP7_75t_SL g2429 ( 
.A(n_2285),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2315),
.B(n_2270),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2267),
.B(n_307),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2297),
.B(n_308),
.Y(n_2432)
);

OR2x2_ASAP7_75t_L g2433 ( 
.A(n_2306),
.B(n_308),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2297),
.B(n_309),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2328),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2282),
.Y(n_2436)
);

OR2x2_ASAP7_75t_L g2437 ( 
.A(n_2293),
.B(n_309),
.Y(n_2437)
);

OAI221xp5_ASAP7_75t_L g2438 ( 
.A1(n_2230),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.C(n_313),
.Y(n_2438)
);

NAND2x1p5_ASAP7_75t_L g2439 ( 
.A(n_2304),
.B(n_310),
.Y(n_2439)
);

AND2x4_ASAP7_75t_L g2440 ( 
.A(n_2298),
.B(n_311),
.Y(n_2440)
);

HB1xp67_ASAP7_75t_L g2441 ( 
.A(n_2257),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2313),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2277),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2308),
.B(n_312),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2279),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_2310),
.B(n_313),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2289),
.B(n_314),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2239),
.B(n_314),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2314),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2296),
.B(n_2291),
.Y(n_2450)
);

INVx2_ASAP7_75t_SL g2451 ( 
.A(n_2337),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2307),
.B(n_315),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2263),
.B(n_315),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_SL g2454 ( 
.A1(n_2222),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2454)
);

INVxp67_ASAP7_75t_SL g2455 ( 
.A(n_2290),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2223),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_2258),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2222),
.B(n_316),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2262),
.B(n_317),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2252),
.B(n_318),
.Y(n_2460)
);

AND2x4_ASAP7_75t_SL g2461 ( 
.A(n_2259),
.B(n_319),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2262),
.B(n_319),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2318),
.B(n_320),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2223),
.Y(n_2464)
);

AOI221xp5_ASAP7_75t_L g2465 ( 
.A1(n_2222),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.C(n_324),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2252),
.B(n_322),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2272),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2252),
.B(n_323),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2272),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2318),
.B(n_324),
.Y(n_2470)
);

OR2x6_ASAP7_75t_L g2471 ( 
.A(n_2327),
.B(n_325),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2272),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2223),
.Y(n_2473)
);

NAND2x1p5_ASAP7_75t_L g2474 ( 
.A(n_2225),
.B(n_325),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2223),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2222),
.B(n_326),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2223),
.Y(n_2477)
);

OR2x2_ASAP7_75t_L g2478 ( 
.A(n_2318),
.B(n_326),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2252),
.B(n_327),
.Y(n_2479)
);

AND2x4_ASAP7_75t_SL g2480 ( 
.A(n_2259),
.B(n_327),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2318),
.B(n_328),
.Y(n_2481)
);

INVx3_ASAP7_75t_L g2482 ( 
.A(n_2258),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2252),
.B(n_328),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2222),
.B(n_329),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2223),
.Y(n_2485)
);

OR2x2_ASAP7_75t_L g2486 ( 
.A(n_2318),
.B(n_329),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2272),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2252),
.B(n_330),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2252),
.B(n_330),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2223),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2255),
.B(n_331),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2272),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2252),
.B(n_331),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2252),
.B(n_332),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_2318),
.B(n_332),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2223),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2223),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2252),
.B(n_333),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2223),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2223),
.Y(n_2500)
);

AND2x4_ASAP7_75t_L g2501 ( 
.A(n_2262),
.B(n_334),
.Y(n_2501)
);

OAI211xp5_ASAP7_75t_SL g2502 ( 
.A1(n_2267),
.A2(n_337),
.B(n_335),
.C(n_336),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2222),
.B(n_335),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2223),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2318),
.B(n_336),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2252),
.B(n_337),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2252),
.B(n_338),
.Y(n_2507)
);

INVxp67_ASAP7_75t_SL g2508 ( 
.A(n_2290),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2223),
.Y(n_2509)
);

NAND2x1_ASAP7_75t_L g2510 ( 
.A(n_2222),
.B(n_338),
.Y(n_2510)
);

NAND3xp33_ASAP7_75t_L g2511 ( 
.A(n_2339),
.B(n_339),
.C(n_340),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2510),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2374),
.B(n_340),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2427),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2423),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2362),
.B(n_341),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2451),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_SL g2518 ( 
.A(n_2435),
.B(n_2342),
.C(n_2367),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2467),
.B(n_342),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2455),
.B(n_343),
.Y(n_2520)
);

INVx5_ASAP7_75t_L g2521 ( 
.A(n_2434),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2469),
.B(n_2472),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2487),
.B(n_344),
.Y(n_2523)
);

AOI22xp33_ASAP7_75t_L g2524 ( 
.A1(n_2395),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_2524)
);

OAI221xp5_ASAP7_75t_SL g2525 ( 
.A1(n_2508),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2357),
.Y(n_2526)
);

OR2x2_ASAP7_75t_L g2527 ( 
.A(n_2413),
.B(n_348),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2492),
.B(n_349),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2396),
.B(n_349),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_L g2530 ( 
.A1(n_2436),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_2530)
);

OAI31xp33_ASAP7_75t_L g2531 ( 
.A1(n_2342),
.A2(n_353),
.A3(n_350),
.B(n_352),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2391),
.B(n_353),
.Y(n_2532)
);

NAND3xp33_ASAP7_75t_L g2533 ( 
.A(n_2341),
.B(n_354),
.C(n_355),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2340),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2482),
.B(n_354),
.Y(n_2535)
);

NAND3xp33_ASAP7_75t_L g2536 ( 
.A(n_2465),
.B(n_357),
.C(n_358),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2378),
.Y(n_2537)
);

AOI211x1_ASAP7_75t_SL g2538 ( 
.A1(n_2409),
.A2(n_2458),
.B(n_2484),
.C(n_2476),
.Y(n_2538)
);

NAND3xp33_ASAP7_75t_SL g2539 ( 
.A(n_2408),
.B(n_358),
.C(n_359),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2426),
.B(n_360),
.Y(n_2540)
);

NAND4xp25_ASAP7_75t_L g2541 ( 
.A(n_2422),
.B(n_363),
.C(n_360),
.D(n_361),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2366),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2416),
.A2(n_364),
.B1(n_361),
.B2(n_363),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2356),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2359),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2457),
.B(n_364),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2372),
.B(n_365),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2441),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2503),
.B(n_2343),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2377),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2456),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2460),
.B(n_365),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2466),
.B(n_367),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2474),
.Y(n_2554)
);

OAI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2351),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2555)
);

NAND4xp25_ASAP7_75t_L g2556 ( 
.A(n_2354),
.B(n_370),
.C(n_368),
.D(n_369),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2468),
.B(n_370),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_L g2558 ( 
.A(n_2346),
.B(n_371),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2479),
.B(n_371),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2348),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2406),
.B(n_372),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2464),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2408),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2473),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2418),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2424),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2345),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2475),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2477),
.Y(n_2569)
);

INVx5_ASAP7_75t_L g2570 ( 
.A(n_2419),
.Y(n_2570)
);

BUFx2_ASAP7_75t_L g2571 ( 
.A(n_2471),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2483),
.B(n_373),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2488),
.B(n_375),
.Y(n_2573)
);

NAND2xp33_ASAP7_75t_R g2574 ( 
.A(n_2489),
.B(n_375),
.Y(n_2574)
);

AOI21xp33_ASAP7_75t_L g2575 ( 
.A1(n_2373),
.A2(n_376),
.B(n_377),
.Y(n_2575)
);

OR2x2_ASAP7_75t_L g2576 ( 
.A(n_2360),
.B(n_376),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2493),
.B(n_377),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_2421),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2494),
.B(n_378),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2353),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2498),
.B(n_2506),
.Y(n_2581)
);

INVx3_ASAP7_75t_L g2582 ( 
.A(n_2459),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2462),
.Y(n_2583)
);

OAI31xp33_ASAP7_75t_L g2584 ( 
.A1(n_2450),
.A2(n_381),
.A3(n_379),
.B(n_380),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2507),
.B(n_382),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2501),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2349),
.B(n_382),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2365),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2442),
.B(n_383),
.Y(n_2589)
);

INVx6_ASAP7_75t_L g2590 ( 
.A(n_2471),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2399),
.B(n_384),
.Y(n_2591)
);

INVxp67_ASAP7_75t_SL g2592 ( 
.A(n_2430),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_SL g2593 ( 
.A(n_2344),
.B(n_385),
.Y(n_2593)
);

NAND2x1p5_ASAP7_75t_L g2594 ( 
.A(n_2440),
.B(n_385),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2485),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2350),
.B(n_386),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2401),
.B(n_386),
.Y(n_2597)
);

OAI33xp33_ASAP7_75t_L g2598 ( 
.A1(n_2452),
.A2(n_390),
.A3(n_392),
.B1(n_387),
.B2(n_388),
.B3(n_391),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2352),
.B(n_387),
.Y(n_2599)
);

AND2x4_ASAP7_75t_L g2600 ( 
.A(n_2368),
.B(n_390),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2490),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2496),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2371),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2355),
.B(n_391),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2380),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2358),
.B(n_393),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2361),
.B(n_393),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2497),
.Y(n_2608)
);

HB1xp67_ASAP7_75t_L g2609 ( 
.A(n_2499),
.Y(n_2609)
);

AND2x4_ASAP7_75t_L g2610 ( 
.A(n_2387),
.B(n_394),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2500),
.B(n_395),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2504),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2385),
.Y(n_2613)
);

AOI221xp5_ASAP7_75t_L g2614 ( 
.A1(n_2438),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.C(n_398),
.Y(n_2614)
);

AND2x4_ASAP7_75t_L g2615 ( 
.A(n_2403),
.B(n_396),
.Y(n_2615)
);

OAI221xp5_ASAP7_75t_L g2616 ( 
.A1(n_2417),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.C(n_400),
.Y(n_2616)
);

BUFx6f_ASAP7_75t_L g2617 ( 
.A(n_2393),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2509),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_2461),
.Y(n_2619)
);

AOI32xp33_ASAP7_75t_L g2620 ( 
.A1(n_2448),
.A2(n_401),
.A3(n_404),
.B1(n_400),
.B2(n_402),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2376),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2480),
.Y(n_2622)
);

INVxp67_ASAP7_75t_SL g2623 ( 
.A(n_2394),
.Y(n_2623)
);

OAI31xp33_ASAP7_75t_L g2624 ( 
.A1(n_2439),
.A2(n_404),
.A3(n_399),
.B(n_401),
.Y(n_2624)
);

AOI21xp5_ASAP7_75t_L g2625 ( 
.A1(n_2398),
.A2(n_405),
.B(n_406),
.Y(n_2625)
);

OAI33xp33_ASAP7_75t_L g2626 ( 
.A1(n_2389),
.A2(n_407),
.A3(n_409),
.B1(n_405),
.B2(n_406),
.B3(n_408),
.Y(n_2626)
);

AO21x2_ASAP7_75t_L g2627 ( 
.A1(n_2412),
.A2(n_407),
.B(n_410),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2400),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2363),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2364),
.Y(n_2630)
);

OAI221xp5_ASAP7_75t_L g2631 ( 
.A1(n_2429),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.C(n_415),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2397),
.Y(n_2632)
);

INVx1_ASAP7_75t_SL g2633 ( 
.A(n_2407),
.Y(n_2633)
);

OR2x6_ASAP7_75t_L g2634 ( 
.A(n_2590),
.B(n_2404),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2566),
.B(n_2491),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2617),
.B(n_2431),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2548),
.B(n_2463),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2569),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2609),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2617),
.B(n_2581),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2590),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2567),
.B(n_2428),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2570),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2580),
.B(n_2582),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2512),
.B(n_2405),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2630),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2570),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2538),
.B(n_2375),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2537),
.Y(n_2649)
);

NAND4xp75_ASAP7_75t_L g2650 ( 
.A(n_2584),
.B(n_2453),
.C(n_2447),
.D(n_2444),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2592),
.B(n_2623),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2629),
.B(n_2449),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2544),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2545),
.Y(n_2654)
);

INVx1_ASAP7_75t_SL g2655 ( 
.A(n_2532),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2551),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2571),
.B(n_2633),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2540),
.B(n_2443),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2562),
.Y(n_2659)
);

AND2x4_ASAP7_75t_SL g2660 ( 
.A(n_2529),
.B(n_2390),
.Y(n_2660)
);

AND2x4_ASAP7_75t_SL g2661 ( 
.A(n_2615),
.B(n_2402),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2619),
.B(n_2425),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2564),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2568),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_L g2665 ( 
.A1(n_2518),
.A2(n_2446),
.B1(n_2445),
.B2(n_2411),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2595),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2622),
.B(n_2381),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2601),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2602),
.Y(n_2669)
);

INVxp67_ASAP7_75t_SL g2670 ( 
.A(n_2574),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2521),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2522),
.B(n_2382),
.Y(n_2672)
);

AOI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2598),
.A2(n_2388),
.B1(n_2420),
.B2(n_2437),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2608),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2611),
.B(n_2383),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2612),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2618),
.Y(n_2677)
);

INVx4_ASAP7_75t_L g2678 ( 
.A(n_2546),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2589),
.B(n_2386),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2621),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2521),
.Y(n_2681)
);

INVx1_ASAP7_75t_SL g2682 ( 
.A(n_2552),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2628),
.Y(n_2683)
);

NAND5xp2_ASAP7_75t_L g2684 ( 
.A(n_2534),
.B(n_2454),
.C(n_2347),
.D(n_2392),
.E(n_2432),
.Y(n_2684)
);

OR2x2_ASAP7_75t_L g2685 ( 
.A(n_2547),
.B(n_2486),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2535),
.B(n_2369),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2583),
.B(n_2370),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2527),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2626),
.A2(n_2410),
.B1(n_2414),
.B2(n_2433),
.Y(n_2689)
);

OR2x2_ASAP7_75t_L g2690 ( 
.A(n_2549),
.B(n_2470),
.Y(n_2690)
);

BUFx3_ASAP7_75t_L g2691 ( 
.A(n_2594),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2627),
.B(n_2478),
.Y(n_2692)
);

INVx1_ASAP7_75t_SL g2693 ( 
.A(n_2553),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2640),
.B(n_2667),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2634),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2652),
.Y(n_2696)
);

AO22x1_ASAP7_75t_L g2697 ( 
.A1(n_2670),
.A2(n_2561),
.B1(n_2520),
.B2(n_2563),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2634),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2657),
.B(n_2526),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2644),
.B(n_2586),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2662),
.B(n_2558),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2646),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2635),
.B(n_2514),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2678),
.B(n_2516),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2682),
.B(n_2625),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2693),
.B(n_2513),
.Y(n_2706)
);

OR2x2_ASAP7_75t_L g2707 ( 
.A(n_2690),
.B(n_2515),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2655),
.B(n_2620),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2651),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2679),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2642),
.B(n_2519),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2688),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2675),
.B(n_2557),
.Y(n_2713)
);

HB1xp67_ASAP7_75t_L g2714 ( 
.A(n_2672),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2643),
.B(n_2647),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2649),
.Y(n_2716)
);

O2A1O1Ixp33_ASAP7_75t_L g2717 ( 
.A1(n_2648),
.A2(n_2541),
.B(n_2556),
.C(n_2525),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2637),
.B(n_2576),
.Y(n_2718)
);

INVxp67_ASAP7_75t_L g2719 ( 
.A(n_2641),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2671),
.B(n_2523),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2660),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2661),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2653),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2654),
.Y(n_2724)
);

BUFx2_ASAP7_75t_L g2725 ( 
.A(n_2691),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2708),
.A2(n_2650),
.B1(n_2673),
.B2(n_2665),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2714),
.Y(n_2727)
);

AOI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2717),
.A2(n_2697),
.B(n_2684),
.Y(n_2728)
);

OAI221xp5_ASAP7_75t_L g2729 ( 
.A1(n_2705),
.A2(n_2692),
.B1(n_2689),
.B2(n_2517),
.C(n_2681),
.Y(n_2729)
);

INVx1_ASAP7_75t_SL g2730 ( 
.A(n_2701),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2703),
.B(n_2686),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2694),
.B(n_2645),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2710),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_2725),
.Y(n_2734)
);

AOI31xp33_ASAP7_75t_L g2735 ( 
.A1(n_2699),
.A2(n_2638),
.A3(n_2639),
.B(n_2636),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2706),
.B(n_2658),
.Y(n_2736)
);

NAND4xp25_ASAP7_75t_L g2737 ( 
.A(n_2715),
.B(n_2656),
.C(n_2663),
.D(n_2659),
.Y(n_2737)
);

OAI21xp5_ASAP7_75t_SL g2738 ( 
.A1(n_2700),
.A2(n_2713),
.B(n_2704),
.Y(n_2738)
);

OAI21xp33_ASAP7_75t_L g2739 ( 
.A1(n_2722),
.A2(n_2666),
.B(n_2664),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2711),
.B(n_2697),
.Y(n_2740)
);

INVxp67_ASAP7_75t_L g2741 ( 
.A(n_2695),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2719),
.B(n_2687),
.Y(n_2742)
);

O2A1O1Ixp33_ASAP7_75t_L g2743 ( 
.A1(n_2709),
.A2(n_2616),
.B(n_2575),
.C(n_2702),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2718),
.B(n_2685),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2696),
.B(n_2572),
.Y(n_2745)
);

AOI31xp33_ASAP7_75t_L g2746 ( 
.A1(n_2730),
.A2(n_2721),
.A3(n_2712),
.B(n_2720),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2726),
.A2(n_2650),
.B1(n_2698),
.B2(n_2707),
.Y(n_2747)
);

OR2x2_ASAP7_75t_L g2748 ( 
.A(n_2744),
.B(n_2734),
.Y(n_2748)
);

NOR2xp67_ASAP7_75t_SL g2749 ( 
.A(n_2733),
.B(n_2511),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2736),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2732),
.Y(n_2751)
);

OAI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2728),
.A2(n_2624),
.B1(n_2531),
.B2(n_2533),
.C(n_2536),
.Y(n_2752)
);

INVx2_ASAP7_75t_SL g2753 ( 
.A(n_2731),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2742),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2745),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2748),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2747),
.A2(n_2740),
.B1(n_2729),
.B2(n_2741),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2746),
.B(n_2738),
.Y(n_2758)
);

O2A1O1Ixp5_ASAP7_75t_L g2759 ( 
.A1(n_2751),
.A2(n_2727),
.B(n_2723),
.C(n_2724),
.Y(n_2759)
);

OAI221xp5_ASAP7_75t_L g2760 ( 
.A1(n_2752),
.A2(n_2743),
.B1(n_2737),
.B2(n_2739),
.C(n_2735),
.Y(n_2760)
);

OR2x2_ASAP7_75t_L g2761 ( 
.A(n_2753),
.B(n_2716),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2749),
.A2(n_2542),
.B1(n_2528),
.B2(n_2550),
.Y(n_2762)
);

OAI32xp33_ASAP7_75t_L g2763 ( 
.A1(n_2750),
.A2(n_2754),
.A3(n_2723),
.B1(n_2755),
.B2(n_2669),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2748),
.Y(n_2764)
);

OAI221xp5_ASAP7_75t_L g2765 ( 
.A1(n_2757),
.A2(n_2560),
.B1(n_2668),
.B2(n_2676),
.C(n_2674),
.Y(n_2765)
);

AOI221xp5_ASAP7_75t_L g2766 ( 
.A1(n_2760),
.A2(n_2683),
.B1(n_2680),
.B2(n_2677),
.C(n_2555),
.Y(n_2766)
);

AOI221xp5_ASAP7_75t_L g2767 ( 
.A1(n_2763),
.A2(n_2539),
.B1(n_2631),
.B2(n_2593),
.C(n_2607),
.Y(n_2767)
);

OAI221xp5_ASAP7_75t_L g2768 ( 
.A1(n_2762),
.A2(n_2554),
.B1(n_2559),
.B2(n_2614),
.C(n_2597),
.Y(n_2768)
);

AOI311xp33_ASAP7_75t_L g2769 ( 
.A1(n_2756),
.A2(n_2606),
.A3(n_2604),
.B(n_2600),
.C(n_2502),
.Y(n_2769)
);

O2A1O1Ixp33_ASAP7_75t_L g2770 ( 
.A1(n_2758),
.A2(n_2384),
.B(n_2587),
.C(n_2577),
.Y(n_2770)
);

AOI21xp33_ASAP7_75t_SL g2771 ( 
.A1(n_2764),
.A2(n_2761),
.B(n_2579),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2759),
.Y(n_2772)
);

NAND4xp25_ASAP7_75t_L g2773 ( 
.A(n_2758),
.B(n_2573),
.C(n_2585),
.D(n_2524),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2764),
.B(n_2588),
.Y(n_2774)
);

OAI31xp33_ASAP7_75t_L g2775 ( 
.A1(n_2760),
.A2(n_2599),
.A3(n_2596),
.B(n_2379),
.Y(n_2775)
);

OAI221xp5_ASAP7_75t_SL g2776 ( 
.A1(n_2757),
.A2(n_2530),
.B1(n_2543),
.B2(n_2578),
.C(n_2495),
.Y(n_2776)
);

OAI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2764),
.A2(n_2481),
.B1(n_2505),
.B2(n_2610),
.Y(n_2777)
);

OAI221xp5_ASAP7_75t_SL g2778 ( 
.A1(n_2757),
.A2(n_2415),
.B1(n_2565),
.B2(n_2605),
.C(n_2603),
.Y(n_2778)
);

O2A1O1Ixp33_ASAP7_75t_L g2779 ( 
.A1(n_2758),
.A2(n_2591),
.B(n_2632),
.C(n_2613),
.Y(n_2779)
);

OAI33xp33_ASAP7_75t_L g2780 ( 
.A1(n_2758),
.A2(n_416),
.A3(n_418),
.B1(n_412),
.B2(n_415),
.B3(n_417),
.Y(n_2780)
);

AO221x1_ASAP7_75t_L g2781 ( 
.A1(n_2756),
.A2(n_419),
.B1(n_416),
.B2(n_417),
.C(n_420),
.Y(n_2781)
);

NAND4xp75_ASAP7_75t_L g2782 ( 
.A(n_2758),
.B(n_421),
.C(n_419),
.D(n_420),
.Y(n_2782)
);

AOI221xp5_ASAP7_75t_L g2783 ( 
.A1(n_2772),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_2783)
);

OAI221xp5_ASAP7_75t_SL g2784 ( 
.A1(n_2775),
.A2(n_424),
.B1(n_426),
.B2(n_423),
.C(n_425),
.Y(n_2784)
);

A2O1A1Ixp33_ASAP7_75t_L g2785 ( 
.A1(n_2770),
.A2(n_426),
.B(n_422),
.C(n_425),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2781),
.B(n_427),
.Y(n_2786)
);

OAI21xp5_ASAP7_75t_SL g2787 ( 
.A1(n_2771),
.A2(n_427),
.B(n_428),
.Y(n_2787)
);

AOI221xp5_ASAP7_75t_L g2788 ( 
.A1(n_2765),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.C(n_431),
.Y(n_2788)
);

OAI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2773),
.A2(n_2768),
.B1(n_2774),
.B2(n_2777),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2779),
.A2(n_429),
.B(n_430),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2782),
.Y(n_2791)
);

OAI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2766),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_2792)
);

AOI221xp5_ASAP7_75t_L g2793 ( 
.A1(n_2767),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.C(n_435),
.Y(n_2793)
);

BUFx2_ASAP7_75t_L g2794 ( 
.A(n_2769),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2778),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2776),
.Y(n_2796)
);

OAI21xp5_ASAP7_75t_SL g2797 ( 
.A1(n_2780),
.A2(n_435),
.B(n_436),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2781),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2772),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2799)
);

AOI221xp5_ASAP7_75t_L g2800 ( 
.A1(n_2772),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.C(n_440),
.Y(n_2800)
);

OAI322xp33_ASAP7_75t_L g2801 ( 
.A1(n_2772),
.A2(n_445),
.A3(n_444),
.B1(n_442),
.B2(n_440),
.C1(n_441),
.C2(n_443),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2781),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2798),
.Y(n_2803)
);

OA22x2_ASAP7_75t_L g2804 ( 
.A1(n_2787),
.A2(n_2797),
.B1(n_2802),
.B2(n_2795),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2786),
.Y(n_2805)
);

AOI221xp5_ASAP7_75t_L g2806 ( 
.A1(n_2801),
.A2(n_446),
.B1(n_442),
.B2(n_443),
.C(n_447),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2791),
.B(n_446),
.Y(n_2807)
);

AOI32xp33_ASAP7_75t_L g2808 ( 
.A1(n_2799),
.A2(n_449),
.A3(n_447),
.B1(n_448),
.B2(n_450),
.Y(n_2808)
);

AOI21xp33_ASAP7_75t_L g2809 ( 
.A1(n_2789),
.A2(n_448),
.B(n_449),
.Y(n_2809)
);

OAI221xp5_ASAP7_75t_L g2810 ( 
.A1(n_2783),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.C(n_454),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2794),
.B(n_451),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2785),
.B(n_453),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2792),
.Y(n_2813)
);

XOR2xp5_ASAP7_75t_L g2814 ( 
.A(n_2796),
.B(n_455),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2800),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2784),
.A2(n_457),
.B(n_458),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2788),
.B(n_458),
.Y(n_2817)
);

OAI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2790),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_2818)
);

OAI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2793),
.A2(n_462),
.B1(n_459),
.B2(n_461),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2797),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_2820)
);

AOI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2797),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_2821)
);

OAI211xp5_ASAP7_75t_SL g2822 ( 
.A1(n_2799),
.A2(n_467),
.B(n_465),
.C(n_466),
.Y(n_2822)
);

AOI221xp5_ASAP7_75t_L g2823 ( 
.A1(n_2805),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.C(n_470),
.Y(n_2823)
);

OAI211xp5_ASAP7_75t_L g2824 ( 
.A1(n_2811),
.A2(n_472),
.B(n_468),
.C(n_471),
.Y(n_2824)
);

AOI221xp5_ASAP7_75t_L g2825 ( 
.A1(n_2809),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.C(n_475),
.Y(n_2825)
);

NAND3xp33_ASAP7_75t_SL g2826 ( 
.A(n_2820),
.B(n_473),
.C(n_476),
.Y(n_2826)
);

OAI211xp5_ASAP7_75t_SL g2827 ( 
.A1(n_2803),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_2827)
);

AOI31xp33_ASAP7_75t_L g2828 ( 
.A1(n_2807),
.A2(n_2821),
.A3(n_2806),
.B(n_2812),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2804),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2808),
.B(n_477),
.Y(n_2830)
);

NOR2x1_ASAP7_75t_L g2831 ( 
.A(n_2814),
.B(n_478),
.Y(n_2831)
);

NAND4xp25_ASAP7_75t_SL g2832 ( 
.A(n_2816),
.B(n_481),
.C(n_479),
.D(n_480),
.Y(n_2832)
);

AOI22xp33_ASAP7_75t_SL g2833 ( 
.A1(n_2813),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_2833)
);

OAI211xp5_ASAP7_75t_L g2834 ( 
.A1(n_2817),
.A2(n_486),
.B(n_484),
.C(n_485),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2815),
.A2(n_484),
.B(n_486),
.Y(n_2835)
);

NAND3xp33_ASAP7_75t_L g2836 ( 
.A(n_2819),
.B(n_489),
.C(n_488),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2822),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2818),
.Y(n_2838)
);

AOI322xp5_ASAP7_75t_L g2839 ( 
.A1(n_2810),
.A2(n_495),
.A3(n_494),
.B1(n_492),
.B2(n_487),
.C1(n_491),
.C2(n_493),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_2803),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2805),
.A2(n_494),
.B1(n_491),
.B2(n_492),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2820),
.B(n_495),
.Y(n_2842)
);

NAND2x1_ASAP7_75t_L g2843 ( 
.A(n_2803),
.B(n_496),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2811),
.B(n_496),
.Y(n_2844)
);

OR2x2_ASAP7_75t_L g2845 ( 
.A(n_2811),
.B(n_497),
.Y(n_2845)
);

NOR4xp25_ASAP7_75t_L g2846 ( 
.A(n_2809),
.B(n_499),
.C(n_497),
.D(n_498),
.Y(n_2846)
);

NOR2x1_ASAP7_75t_L g2847 ( 
.A(n_2811),
.B(n_498),
.Y(n_2847)
);

AOI221xp5_ASAP7_75t_L g2848 ( 
.A1(n_2805),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.C(n_503),
.Y(n_2848)
);

AOI211xp5_ASAP7_75t_SL g2849 ( 
.A1(n_2811),
.A2(n_503),
.B(n_500),
.C(n_502),
.Y(n_2849)
);

OAI322xp33_ASAP7_75t_L g2850 ( 
.A1(n_2811),
.A2(n_509),
.A3(n_508),
.B1(n_506),
.B2(n_504),
.C1(n_505),
.C2(n_507),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2812),
.Y(n_2851)
);

AOI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2805),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2805),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.Y(n_2853)
);

XNOR2xp5_ASAP7_75t_L g2854 ( 
.A(n_2814),
.B(n_510),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2804),
.Y(n_2855)
);

NOR2x1_ASAP7_75t_L g2856 ( 
.A(n_2829),
.B(n_510),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2855),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_2857)
);

INVxp67_ASAP7_75t_SL g2858 ( 
.A(n_2854),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2847),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2851),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_2860)
);

NOR2x1_ASAP7_75t_L g2861 ( 
.A(n_2840),
.B(n_514),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2831),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2845),
.Y(n_2863)
);

INVxp33_ASAP7_75t_SL g2864 ( 
.A(n_2844),
.Y(n_2864)
);

NOR4xp25_ASAP7_75t_L g2865 ( 
.A(n_2828),
.B(n_517),
.C(n_515),
.D(n_516),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2843),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2840),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2840),
.Y(n_2868)
);

INVxp33_ASAP7_75t_L g2869 ( 
.A(n_2846),
.Y(n_2869)
);

AOI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2826),
.A2(n_2842),
.B1(n_2832),
.B2(n_2827),
.Y(n_2870)
);

NOR2x1_ASAP7_75t_L g2871 ( 
.A(n_2850),
.B(n_515),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2837),
.Y(n_2872)
);

HB1xp67_ASAP7_75t_L g2873 ( 
.A(n_2849),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2838),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2833),
.B(n_516),
.Y(n_2875)
);

NOR2x1_ASAP7_75t_L g2876 ( 
.A(n_2830),
.B(n_517),
.Y(n_2876)
);

NAND3xp33_ASAP7_75t_L g2877 ( 
.A(n_2825),
.B(n_518),
.C(n_519),
.Y(n_2877)
);

OR2x2_ASAP7_75t_L g2878 ( 
.A(n_2836),
.B(n_518),
.Y(n_2878)
);

AOI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2834),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2841),
.B(n_520),
.Y(n_2880)
);

NOR2xp67_ASAP7_75t_L g2881 ( 
.A(n_2853),
.B(n_522),
.Y(n_2881)
);

NOR2x1_ASAP7_75t_L g2882 ( 
.A(n_2824),
.B(n_522),
.Y(n_2882)
);

AOI22xp33_ASAP7_75t_SL g2883 ( 
.A1(n_2835),
.A2(n_2839),
.B1(n_2852),
.B2(n_2848),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2823),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2847),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2847),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2840),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2855),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.Y(n_2888)
);

NOR2x1_ASAP7_75t_L g2889 ( 
.A(n_2829),
.B(n_524),
.Y(n_2889)
);

NOR2x1p5_ASAP7_75t_L g2890 ( 
.A(n_2829),
.B(n_525),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2849),
.B(n_526),
.Y(n_2891)
);

AOI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2855),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_2892)
);

OAI211xp5_ASAP7_75t_SL g2893 ( 
.A1(n_2829),
.A2(n_530),
.B(n_527),
.C(n_528),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2847),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2847),
.Y(n_2895)
);

NOR2x1_ASAP7_75t_L g2896 ( 
.A(n_2829),
.B(n_530),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2873),
.Y(n_2897)
);

NOR2x1_ASAP7_75t_L g2898 ( 
.A(n_2868),
.B(n_531),
.Y(n_2898)
);

OR2x2_ASAP7_75t_L g2899 ( 
.A(n_2887),
.B(n_532),
.Y(n_2899)
);

NOR2x1_ASAP7_75t_L g2900 ( 
.A(n_2867),
.B(n_532),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2865),
.B(n_533),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2869),
.B(n_533),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2890),
.B(n_534),
.Y(n_2903)
);

NOR2x1p5_ASAP7_75t_L g2904 ( 
.A(n_2875),
.B(n_534),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2861),
.B(n_535),
.Y(n_2905)
);

NAND4xp75_ASAP7_75t_L g2906 ( 
.A(n_2856),
.B(n_537),
.C(n_535),
.D(n_536),
.Y(n_2906)
);

NAND4xp75_ASAP7_75t_L g2907 ( 
.A(n_2889),
.B(n_538),
.C(n_536),
.D(n_537),
.Y(n_2907)
);

XNOR2xp5_ASAP7_75t_L g2908 ( 
.A(n_2870),
.B(n_539),
.Y(n_2908)
);

XNOR2xp5_ASAP7_75t_L g2909 ( 
.A(n_2864),
.B(n_539),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2896),
.B(n_540),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2862),
.B(n_540),
.Y(n_2911)
);

NAND4xp75_ASAP7_75t_L g2912 ( 
.A(n_2876),
.B(n_544),
.C(n_542),
.D(n_543),
.Y(n_2912)
);

NOR2x1_ASAP7_75t_L g2913 ( 
.A(n_2878),
.B(n_542),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2871),
.B(n_545),
.Y(n_2914)
);

NOR3xp33_ASAP7_75t_L g2915 ( 
.A(n_2858),
.B(n_545),
.C(n_546),
.Y(n_2915)
);

NOR2x1_ASAP7_75t_L g2916 ( 
.A(n_2893),
.B(n_546),
.Y(n_2916)
);

AND5x1_ASAP7_75t_L g2917 ( 
.A(n_2879),
.B(n_2892),
.C(n_2888),
.D(n_2857),
.E(n_2883),
.Y(n_2917)
);

NAND4xp75_ASAP7_75t_L g2918 ( 
.A(n_2882),
.B(n_550),
.C(n_547),
.D(n_549),
.Y(n_2918)
);

NAND4xp75_ASAP7_75t_L g2919 ( 
.A(n_2859),
.B(n_551),
.C(n_547),
.D(n_549),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2885),
.B(n_551),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2866),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2886),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2891),
.Y(n_2923)
);

AND3x2_ASAP7_75t_L g2924 ( 
.A(n_2894),
.B(n_2895),
.C(n_2874),
.Y(n_2924)
);

INVxp33_ASAP7_75t_L g2925 ( 
.A(n_2881),
.Y(n_2925)
);

NOR2x1_ASAP7_75t_L g2926 ( 
.A(n_2877),
.B(n_552),
.Y(n_2926)
);

AND2x2_ASAP7_75t_SL g2927 ( 
.A(n_2880),
.B(n_552),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2860),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_2863),
.Y(n_2929)
);

NAND2x1p5_ASAP7_75t_L g2930 ( 
.A(n_2884),
.B(n_555),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2872),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2873),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2887),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2858),
.A2(n_560),
.B1(n_557),
.B2(n_559),
.Y(n_2934)
);

NAND4xp75_ASAP7_75t_L g2935 ( 
.A(n_2856),
.B(n_562),
.C(n_560),
.D(n_561),
.Y(n_2935)
);

NAND4xp75_ASAP7_75t_L g2936 ( 
.A(n_2856),
.B(n_564),
.C(n_562),
.D(n_563),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2887),
.B(n_563),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2873),
.Y(n_2938)
);

NOR2x1_ASAP7_75t_L g2939 ( 
.A(n_2868),
.B(n_564),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2873),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2887),
.B(n_565),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2861),
.Y(n_2942)
);

XOR2xp5_ASAP7_75t_L g2943 ( 
.A(n_2873),
.B(n_565),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2873),
.Y(n_2944)
);

OR3x2_ASAP7_75t_L g2945 ( 
.A(n_2897),
.B(n_566),
.C(n_567),
.Y(n_2945)
);

AOI22xp5_ASAP7_75t_L g2946 ( 
.A1(n_2922),
.A2(n_2923),
.B1(n_2938),
.B2(n_2932),
.Y(n_2946)
);

O2A1O1Ixp33_ASAP7_75t_L g2947 ( 
.A1(n_2940),
.A2(n_569),
.B(n_566),
.C(n_568),
.Y(n_2947)
);

AND3x4_ASAP7_75t_L g2948 ( 
.A(n_2916),
.B(n_568),
.C(n_569),
.Y(n_2948)
);

OAI21xp33_ASAP7_75t_SL g2949 ( 
.A1(n_2944),
.A2(n_570),
.B(n_571),
.Y(n_2949)
);

O2A1O1Ixp5_ASAP7_75t_L g2950 ( 
.A1(n_2921),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_2950)
);

AOI211xp5_ASAP7_75t_SL g2951 ( 
.A1(n_2902),
.A2(n_574),
.B(n_572),
.C(n_573),
.Y(n_2951)
);

OAI211xp5_ASAP7_75t_SL g2952 ( 
.A1(n_2929),
.A2(n_575),
.B(n_573),
.C(n_574),
.Y(n_2952)
);

AOI221xp5_ASAP7_75t_L g2953 ( 
.A1(n_2914),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.C(n_578),
.Y(n_2953)
);

INVx1_ASAP7_75t_SL g2954 ( 
.A(n_2901),
.Y(n_2954)
);

NAND3xp33_ASAP7_75t_L g2955 ( 
.A(n_2924),
.B(n_576),
.C(n_577),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2910),
.Y(n_2956)
);

AND4x1_ASAP7_75t_L g2957 ( 
.A(n_2898),
.B(n_581),
.C(n_579),
.D(n_580),
.Y(n_2957)
);

OA22x2_ASAP7_75t_L g2958 ( 
.A1(n_2943),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_2958)
);

OAI221xp5_ASAP7_75t_L g2959 ( 
.A1(n_2939),
.A2(n_584),
.B1(n_582),
.B2(n_583),
.C(n_585),
.Y(n_2959)
);

AOI221xp5_ASAP7_75t_L g2960 ( 
.A1(n_2903),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.C(n_588),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2905),
.A2(n_586),
.B(n_588),
.Y(n_2961)
);

NAND4xp25_ASAP7_75t_L g2962 ( 
.A(n_2900),
.B(n_591),
.C(n_589),
.D(n_590),
.Y(n_2962)
);

A2O1A1Ixp33_ASAP7_75t_L g2963 ( 
.A1(n_2920),
.A2(n_591),
.B(n_589),
.C(n_590),
.Y(n_2963)
);

OAI32xp33_ASAP7_75t_L g2964 ( 
.A1(n_2899),
.A2(n_595),
.A3(n_592),
.B1(n_593),
.B2(n_596),
.Y(n_2964)
);

O2A1O1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2942),
.A2(n_596),
.B(n_593),
.C(n_595),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2913),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_2966)
);

AND4x1_ASAP7_75t_L g2967 ( 
.A(n_2911),
.B(n_601),
.C(n_599),
.D(n_600),
.Y(n_2967)
);

AOI322xp5_ASAP7_75t_L g2968 ( 
.A1(n_2926),
.A2(n_606),
.A3(n_605),
.B1(n_603),
.B2(n_601),
.C1(n_602),
.C2(n_604),
.Y(n_2968)
);

AOI222xp33_ASAP7_75t_L g2969 ( 
.A1(n_2927),
.A2(n_605),
.B1(n_608),
.B2(n_603),
.C1(n_604),
.C2(n_606),
.Y(n_2969)
);

OAI211xp5_ASAP7_75t_L g2970 ( 
.A1(n_2934),
.A2(n_610),
.B(n_608),
.C(n_609),
.Y(n_2970)
);

XOR2xp5_ASAP7_75t_L g2971 ( 
.A(n_2909),
.B(n_609),
.Y(n_2971)
);

AOI221x1_ASAP7_75t_L g2972 ( 
.A1(n_2915),
.A2(n_612),
.B1(n_610),
.B2(n_611),
.C(n_613),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2906),
.B(n_612),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2904),
.A2(n_616),
.B1(n_614),
.B2(n_615),
.Y(n_2974)
);

XNOR2xp5_ASAP7_75t_L g2975 ( 
.A(n_2908),
.B(n_614),
.Y(n_2975)
);

OAI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2930),
.A2(n_2918),
.B1(n_2935),
.B2(n_2907),
.Y(n_2976)
);

AOI211xp5_ASAP7_75t_L g2977 ( 
.A1(n_2928),
.A2(n_617),
.B(n_615),
.C(n_616),
.Y(n_2977)
);

NAND3xp33_ASAP7_75t_SL g2978 ( 
.A(n_2925),
.B(n_618),
.C(n_619),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2937),
.A2(n_621),
.B(n_618),
.C(n_620),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2933),
.A2(n_620),
.B(n_621),
.Y(n_2980)
);

O2A1O1Ixp5_ASAP7_75t_L g2981 ( 
.A1(n_2931),
.A2(n_624),
.B(n_622),
.C(n_623),
.Y(n_2981)
);

AOI221xp5_ASAP7_75t_L g2982 ( 
.A1(n_2941),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.C(n_625),
.Y(n_2982)
);

AOI221xp5_ASAP7_75t_L g2983 ( 
.A1(n_2917),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.C(n_628),
.Y(n_2983)
);

AOI211x1_ASAP7_75t_L g2984 ( 
.A1(n_2936),
.A2(n_629),
.B(n_626),
.C(n_628),
.Y(n_2984)
);

NOR3xp33_ASAP7_75t_L g2985 ( 
.A(n_2912),
.B(n_2919),
.C(n_629),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2910),
.Y(n_2986)
);

AOI211xp5_ASAP7_75t_SL g2987 ( 
.A1(n_2897),
.A2(n_632),
.B(n_630),
.C(n_631),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2957),
.Y(n_2988)
);

BUFx2_ASAP7_75t_L g2989 ( 
.A(n_2949),
.Y(n_2989)
);

AND2x4_ASAP7_75t_L g2990 ( 
.A(n_2946),
.B(n_631),
.Y(n_2990)
);

NOR2x1_ASAP7_75t_L g2991 ( 
.A(n_2955),
.B(n_632),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2958),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2945),
.Y(n_2993)
);

NOR2x1_ASAP7_75t_L g2994 ( 
.A(n_2978),
.B(n_633),
.Y(n_2994)
);

AOI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2954),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_2995)
);

INVx5_ASAP7_75t_L g2996 ( 
.A(n_2967),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2959),
.A2(n_2966),
.B1(n_2974),
.B2(n_2971),
.Y(n_2997)
);

INVx4_ASAP7_75t_L g2998 ( 
.A(n_2956),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2948),
.Y(n_2999)
);

HB1xp67_ASAP7_75t_L g3000 ( 
.A(n_2986),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2962),
.B(n_634),
.Y(n_3001)
);

NOR2xp33_ASAP7_75t_L g3002 ( 
.A(n_2952),
.B(n_635),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2984),
.Y(n_3003)
);

HB1xp67_ASAP7_75t_L g3004 ( 
.A(n_2975),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2987),
.B(n_636),
.Y(n_3005)
);

NAND3x1_ASAP7_75t_L g3006 ( 
.A(n_2985),
.B(n_2973),
.C(n_2983),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2976),
.Y(n_3007)
);

AND3x2_ASAP7_75t_L g3008 ( 
.A(n_2977),
.B(n_2953),
.C(n_2960),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2951),
.B(n_636),
.Y(n_3009)
);

XNOR2x1_ASAP7_75t_L g3010 ( 
.A(n_2969),
.B(n_637),
.Y(n_3010)
);

AND2x4_ASAP7_75t_L g3011 ( 
.A(n_2980),
.B(n_637),
.Y(n_3011)
);

NAND3xp33_ASAP7_75t_L g3012 ( 
.A(n_2968),
.B(n_638),
.C(n_639),
.Y(n_3012)
);

AND2x4_ASAP7_75t_L g3013 ( 
.A(n_2972),
.B(n_638),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2979),
.B(n_639),
.Y(n_3014)
);

OR2x6_ASAP7_75t_L g3015 ( 
.A(n_2961),
.B(n_640),
.Y(n_3015)
);

NOR2x1_ASAP7_75t_L g3016 ( 
.A(n_2947),
.B(n_2963),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2950),
.B(n_640),
.Y(n_3017)
);

INVxp67_ASAP7_75t_L g3018 ( 
.A(n_2970),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2981),
.B(n_641),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2989),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_3000),
.A2(n_2965),
.B(n_2964),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_3013),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2988),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2996),
.B(n_2982),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2996),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_3005),
.Y(n_3026)
);

AND2x2_ASAP7_75t_L g3027 ( 
.A(n_2998),
.B(n_641),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2994),
.Y(n_3028)
);

INVx3_ASAP7_75t_L g3029 ( 
.A(n_2990),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_3003),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_3009),
.Y(n_3031)
);

NAND3xp33_ASAP7_75t_L g3032 ( 
.A(n_3007),
.B(n_3004),
.C(n_2992),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_3019),
.Y(n_3033)
);

HB1xp67_ASAP7_75t_L g3034 ( 
.A(n_2999),
.Y(n_3034)
);

INVx3_ASAP7_75t_L g3035 ( 
.A(n_3011),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_3017),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_3015),
.Y(n_3037)
);

INVx3_ASAP7_75t_L g3038 ( 
.A(n_3015),
.Y(n_3038)
);

NAND3xp33_ASAP7_75t_SL g3039 ( 
.A(n_2993),
.B(n_642),
.C(n_643),
.Y(n_3039)
);

OR2x2_ASAP7_75t_L g3040 ( 
.A(n_3010),
.B(n_3018),
.Y(n_3040)
);

INVx2_ASAP7_75t_SL g3041 ( 
.A(n_2991),
.Y(n_3041)
);

INVx1_ASAP7_75t_SL g3042 ( 
.A(n_3014),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_3006),
.Y(n_3043)
);

AND3x4_ASAP7_75t_L g3044 ( 
.A(n_3016),
.B(n_643),
.C(n_644),
.Y(n_3044)
);

XNOR2xp5_ASAP7_75t_L g3045 ( 
.A(n_2997),
.B(n_3008),
.Y(n_3045)
);

HB1xp67_ASAP7_75t_L g3046 ( 
.A(n_3044),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_3022),
.Y(n_3047)
);

XNOR2xp5_ASAP7_75t_L g3048 ( 
.A(n_3045),
.B(n_3012),
.Y(n_3048)
);

BUFx2_ASAP7_75t_L g3049 ( 
.A(n_3020),
.Y(n_3049)
);

XNOR2xp5_ASAP7_75t_L g3050 ( 
.A(n_3032),
.B(n_2995),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_3038),
.B(n_3002),
.Y(n_3051)
);

INVxp67_ASAP7_75t_L g3052 ( 
.A(n_3027),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_3028),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_3025),
.B(n_3033),
.Y(n_3054)
);

HB1xp67_ASAP7_75t_L g3055 ( 
.A(n_3034),
.Y(n_3055)
);

AOI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_3043),
.A2(n_3001),
.B1(n_647),
.B2(n_645),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_3036),
.Y(n_3057)
);

INVx1_ASAP7_75t_SL g3058 ( 
.A(n_3055),
.Y(n_3058)
);

OAI22xp5_ASAP7_75t_SL g3059 ( 
.A1(n_3049),
.A2(n_3023),
.B1(n_3041),
.B2(n_3030),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_3046),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_3047),
.Y(n_3061)
);

OAI22xp33_ASAP7_75t_L g3062 ( 
.A1(n_3054),
.A2(n_3040),
.B1(n_3024),
.B2(n_3026),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_3053),
.A2(n_3039),
.B1(n_3031),
.B2(n_3042),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_3052),
.B(n_3037),
.Y(n_3064)
);

AO22x1_ASAP7_75t_L g3065 ( 
.A1(n_3057),
.A2(n_3035),
.B1(n_3029),
.B2(n_3021),
.Y(n_3065)
);

OAI22xp5_ASAP7_75t_L g3066 ( 
.A1(n_3050),
.A2(n_647),
.B1(n_645),
.B2(n_646),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_SL g3067 ( 
.A(n_3058),
.B(n_3048),
.Y(n_3067)
);

OAI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_3060),
.A2(n_3056),
.B1(n_3051),
.B2(n_649),
.Y(n_3068)
);

OAI22xp5_ASAP7_75t_L g3069 ( 
.A1(n_3062),
.A2(n_650),
.B1(n_646),
.B2(n_648),
.Y(n_3069)
);

OAI22xp5_ASAP7_75t_SL g3070 ( 
.A1(n_3059),
.A2(n_3061),
.B1(n_3063),
.B2(n_3064),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3065),
.Y(n_3071)
);

NAND2x1p5_ASAP7_75t_L g3072 ( 
.A(n_3066),
.B(n_648),
.Y(n_3072)
);

HB1xp67_ASAP7_75t_L g3073 ( 
.A(n_3058),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_3058),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_3073),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3070),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_3074),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_3071),
.B(n_651),
.Y(n_3078)
);

CKINVDCx20_ASAP7_75t_R g3079 ( 
.A(n_3067),
.Y(n_3079)
);

OAI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_3069),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_3072),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_3068),
.Y(n_3082)
);

OAI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_3079),
.A2(n_653),
.B(n_654),
.Y(n_3083)
);

AOI21xp5_ASAP7_75t_L g3084 ( 
.A1(n_3075),
.A2(n_655),
.B(n_656),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3076),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3081),
.Y(n_3086)
);

OAI21x1_ASAP7_75t_SL g3087 ( 
.A1(n_3078),
.A2(n_656),
.B(n_657),
.Y(n_3087)
);

XNOR2xp5_ASAP7_75t_L g3088 ( 
.A(n_3085),
.B(n_3082),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_3086),
.B(n_3080),
.Y(n_3089)
);

AOI21xp33_ASAP7_75t_SL g3090 ( 
.A1(n_3087),
.A2(n_3077),
.B(n_657),
.Y(n_3090)
);

AOI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_3088),
.A2(n_3083),
.B1(n_3084),
.B2(n_660),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_L g3092 ( 
.A1(n_3089),
.A2(n_661),
.B1(n_658),
.B2(n_659),
.Y(n_3092)
);

OA21x2_ASAP7_75t_L g3093 ( 
.A1(n_3092),
.A2(n_3090),
.B(n_658),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_3093),
.A2(n_3091),
.B(n_661),
.Y(n_3094)
);

AOI211xp5_ASAP7_75t_L g3095 ( 
.A1(n_3094),
.A2(n_664),
.B(n_662),
.C(n_663),
.Y(n_3095)
);


endmodule