module fake_jpeg_30773_n_60 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_20),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_23),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_18),
.B(n_7),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_1),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_27),
.B(n_25),
.C(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_43),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_17),
.B1(n_15),
.B2(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.C(n_40),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_49),
.C(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_53),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_44),
.B(n_57),
.C(n_52),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_36),
.B(n_48),
.Y(n_60)
);


endmodule