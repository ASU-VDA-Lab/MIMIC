module fake_jpeg_1777_n_86 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_33),
.Y(n_36)
);

OR2x2_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_45),
.Y(n_55)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_28),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_37),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_56),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_39),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_40),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_28),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_12),
.C(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_27),
.B1(n_26),
.B2(n_4),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_2),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_3),
.B(n_4),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_63),
.C(n_58),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_58),
.B1(n_6),
.B2(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

BUFx12f_ASAP7_75t_SL g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.Y(n_79)
);

OA21x2_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_5),
.B(n_7),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_71),
.B1(n_9),
.B2(n_11),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_79),
.C(n_13),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_8),
.CI(n_15),
.CON(n_85),
.SN(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_16),
.Y(n_86)
);


endmodule