module fake_jpeg_15572_n_199 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_25),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_30),
.Y(n_45)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_14),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_17),
.C(n_14),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_19),
.C(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_54),
.B1(n_46),
.B2(n_29),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_67),
.B1(n_30),
.B2(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_45),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_53),
.Y(n_75)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_29),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_68),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_40),
.B(n_49),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_74),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_53),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_75),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_38),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_82),
.B1(n_57),
.B2(n_47),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_39),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_59),
.B1(n_44),
.B2(n_37),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_86),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_47),
.B1(n_41),
.B2(n_34),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_56),
.B1(n_29),
.B2(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_92),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_60),
.A3(n_64),
.B1(n_56),
.B2(n_70),
.C1(n_62),
.C2(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_102),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_103),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_67),
.B1(n_54),
.B2(n_60),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_100),
.B(n_79),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_71),
.B1(n_47),
.B2(n_59),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_45),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_61),
.B1(n_44),
.B2(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_77),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_112),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_121),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_101),
.B1(n_98),
.B2(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_104),
.B1(n_95),
.B2(n_100),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_82),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_74),
.B(n_78),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_22),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_76),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_94),
.C(n_104),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.C(n_134),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_94),
.C(n_75),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_133),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_48),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_100),
.B1(n_82),
.B2(n_78),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_138),
.B(n_117),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_37),
.C(n_52),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_22),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_52),
.B1(n_0),
.B2(n_3),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_130),
.B(n_132),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_22),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_122),
.C(n_111),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_114),
.C(n_22),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_107),
.B(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_37),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_109),
.C(n_107),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_126),
.C(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_142),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_124),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_154),
.C(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_109),
.C(n_138),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_146),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_1),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_158),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_37),
.C(n_22),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_141),
.C(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_173),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_145),
.B1(n_151),
.B2(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_174),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_152),
.C(n_143),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.C(n_5),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_159),
.C(n_163),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_174)
);

OAI21x1_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_173),
.B(n_168),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_9),
.B(n_10),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

AOI31xp67_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_6),
.C(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_185),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_181),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_9),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_177),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_184),
.B(n_11),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_10),
.B(n_11),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_191),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_195),
.B(n_11),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_R g196 ( 
.A(n_194),
.B(n_189),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.C(n_12),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_12),
.Y(n_199)
);


endmodule