module fake_jpeg_8621_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_31),
.B1(n_32),
.B2(n_28),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_59),
.B1(n_61),
.B2(n_42),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_31),
.B1(n_32),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_31),
.B1(n_32),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_24),
.B1(n_30),
.B2(n_28),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_18),
.B(n_23),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_41),
.B(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_39),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_17),
.B1(n_41),
.B2(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_17),
.B1(n_18),
.B2(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_72),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_34),
.B(n_20),
.Y(n_103)
);

OAI22x1_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_87),
.B1(n_20),
.B2(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_78),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_34),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_13),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_1),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_44),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_44),
.B1(n_29),
.B2(n_57),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_57),
.B(n_40),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_40),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_52),
.B1(n_57),
.B2(n_38),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_102),
.B1(n_79),
.B2(n_92),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_80),
.B(n_90),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_107),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_38),
.B1(n_29),
.B2(n_35),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_114),
.B1(n_75),
.B2(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_38),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_40),
.B(n_35),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_112),
.B(n_113),
.Y(n_132)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_88),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_38),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_122),
.B1(n_128),
.B2(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_71),
.B1(n_86),
.B2(n_66),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_126),
.A2(n_139),
.B(n_40),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_66),
.B1(n_91),
.B2(n_88),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_91),
.C(n_89),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_135),
.C(n_40),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_131),
.B1(n_147),
.B2(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_91),
.B1(n_83),
.B2(n_38),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_112),
.B1(n_113),
.B2(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_27),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_40),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_27),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_35),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_141),
.B(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_67),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_40),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_15),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_40),
.B1(n_54),
.B2(n_46),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_13),
.C(n_4),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_145),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_94),
.A2(n_40),
.B(n_4),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_119),
.B(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_54),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_163),
.B(n_144),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_103),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_132),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_152),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_96),
.B1(n_104),
.B2(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_96),
.B1(n_97),
.B2(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_167),
.C(n_129),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_126),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_97),
.B1(n_46),
.B2(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_46),
.B1(n_110),
.B2(n_7),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_166),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_141),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_171),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_150),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_190),
.C(n_199),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_201),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_165),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_130),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_133),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_161),
.B1(n_177),
.B2(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_156),
.B1(n_175),
.B2(n_149),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_178),
.B1(n_191),
.B2(n_201),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_186),
.C(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_216),
.C(n_220),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_151),
.B1(n_120),
.B2(n_149),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_178),
.B1(n_179),
.B2(n_199),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_163),
.C(n_155),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_155),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_217),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_197),
.B1(n_192),
.B2(n_185),
.C(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_159),
.C(n_110),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_1),
.B1(n_6),
.B2(n_8),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_187),
.C(n_184),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_233),
.C(n_236),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_10),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_208),
.B1(n_209),
.B2(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_217),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_201),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_179),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_189),
.C(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_203),
.B1(n_212),
.B2(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_227),
.B1(n_228),
.B2(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_220),
.C(n_216),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.C(n_225),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_207),
.C(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_6),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_249),
.Y(n_250)
);

NOR2x1_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_247),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_6),
.B(n_8),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_10),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_222),
.C(n_236),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_257),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_259),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_232),
.C(n_229),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_244),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_258),
.B1(n_246),
.B2(n_12),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_258),
.B(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_11),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_10),
.B(n_11),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_261),
.C(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_12),
.B1(n_270),
.B2(n_271),
.C(n_274),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_276),
.Y(n_279)
);


endmodule