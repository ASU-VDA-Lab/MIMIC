module fake_aes_567_n_43 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_43);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_9), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
AOI22x1_ASAP7_75t_L g20 ( .A1(n_12), .A2(n_10), .B1(n_2), .B2(n_3), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_12), .B(n_0), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_15), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_14), .B(n_2), .Y(n_23) );
AOI22xp33_ASAP7_75t_SL g24 ( .A1(n_20), .A2(n_17), .B1(n_16), .B2(n_13), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_16), .B1(n_5), .B2(n_6), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_18), .B(n_3), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_19), .B(n_18), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_24), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_21), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_30), .B(n_23), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_28), .B(n_19), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_29), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_25), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
A2O1A1Ixp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_20), .B(n_6), .C(n_7), .Y(n_36) );
AND2x2_ASAP7_75t_L g37 ( .A(n_33), .B(n_5), .Y(n_37) );
AND2x2_ASAP7_75t_L g38 ( .A(n_34), .B(n_7), .Y(n_38) );
OAI221xp5_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_34), .B1(n_35), .B2(n_37), .C(n_38), .Y(n_39) );
BUFx6f_ASAP7_75t_L g40 ( .A(n_36), .Y(n_40) );
INVx2_ASAP7_75t_SL g41 ( .A(n_40), .Y(n_41) );
HB1xp67_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
AOI22xp33_ASAP7_75t_L g43 ( .A1(n_42), .A2(n_40), .B1(n_41), .B2(n_39), .Y(n_43) );
endmodule