module fake_jpeg_2838_n_711 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_711);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_711;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_566;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_3),
.B(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_11),
.B(n_17),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_66),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_10),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_67),
.Y(n_192)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_68),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_69),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_23),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_70),
.A2(n_38),
.B1(n_47),
.B2(n_39),
.Y(n_174)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_71),
.Y(n_229)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_23),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_77),
.Y(n_152)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_9),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_84),
.Y(n_214)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_87),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_9),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_99),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_11),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_44),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_107),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_11),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_19),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_108),
.B(n_114),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_19),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_29),
.B(n_19),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_119),
.B(n_121),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_29),
.B(n_18),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_25),
.Y(n_126)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_21),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_36),
.Y(n_128)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_36),
.Y(n_130)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_28),
.Y(n_131)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_28),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_78),
.A2(n_51),
.B1(n_35),
.B2(n_57),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_140),
.A2(n_160),
.B1(n_191),
.B2(n_220),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_75),
.B(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_150),
.B(n_184),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_37),
.B1(n_52),
.B2(n_34),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_151),
.B(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_99),
.A2(n_60),
.B1(n_47),
.B2(n_39),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_72),
.A2(n_44),
.B(n_52),
.C(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_161),
.B(n_174),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_91),
.A2(n_40),
.B1(n_27),
.B2(n_32),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_162),
.A2(n_164),
.B1(n_169),
.B2(n_82),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_93),
.A2(n_24),
.B1(n_40),
.B2(n_32),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_96),
.A2(n_24),
.B1(n_35),
.B2(n_60),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_72),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_176),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_88),
.B(n_41),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_182),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_38),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_88),
.A2(n_51),
.B1(n_35),
.B2(n_28),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_65),
.B(n_41),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_196),
.B(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_100),
.B(n_57),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_197),
.B(n_218),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_95),
.Y(n_208)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_213),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_62),
.B(n_57),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_62),
.B(n_57),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_63),
.A2(n_57),
.B1(n_28),
.B2(n_46),
.Y(n_220)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_71),
.Y(n_223)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_224),
.Y(n_310)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_83),
.Y(n_225)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_101),
.Y(n_226)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_104),
.B(n_12),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_126),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_152),
.A2(n_103),
.B1(n_97),
.B2(n_111),
.Y(n_231)
);

AOI22x1_ASAP7_75t_L g354 ( 
.A1(n_231),
.A2(n_294),
.B1(n_215),
.B2(n_228),
.Y(n_354)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g319 ( 
.A(n_232),
.Y(n_319)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_234),
.Y(n_336)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_235),
.Y(n_342)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_237),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_69),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_240),
.B(n_241),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_79),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_243),
.B(n_277),
.Y(n_351)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_246),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_248),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_162),
.A2(n_115),
.B1(n_116),
.B2(n_73),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_250),
.A2(n_264),
.B1(n_289),
.B2(n_212),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_251),
.B(n_263),
.Y(n_372)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_254),
.Y(n_355)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_136),
.Y(n_256)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_155),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g369 ( 
.A(n_259),
.Y(n_369)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_152),
.A2(n_44),
.B(n_126),
.C(n_46),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_262),
.B(n_151),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_190),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_158),
.Y(n_265)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_182),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_280),
.Y(n_315)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

CKINVDCx12_ASAP7_75t_R g332 ( 
.A(n_268),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_137),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_287),
.Y(n_312)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_167),
.A2(n_84),
.B1(n_44),
.B2(n_74),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_276),
.A2(n_278),
.B1(n_279),
.B2(n_286),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_153),
.B(n_209),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_144),
.A2(n_153),
.B1(n_209),
.B2(n_204),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_144),
.A2(n_80),
.B1(n_81),
.B2(n_131),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_135),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_139),
.Y(n_281)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_130),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_195),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_185),
.Y(n_283)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_283),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_167),
.B(n_128),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_284),
.B(n_288),
.Y(n_373)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_285),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_204),
.A2(n_124),
.B1(n_123),
.B2(n_25),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_166),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_142),
.B(n_18),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_164),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_290),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_169),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_291),
.A2(n_187),
.B1(n_165),
.B2(n_203),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_192),
.B(n_1),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_296),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_222),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_300),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_191),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_186),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_295),
.Y(n_371)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_216),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_186),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_297),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_201),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_298),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_143),
.B(n_14),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_159),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_306),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_201),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_294),
.Y(n_348)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_149),
.B(n_163),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_308),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_140),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_217),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_138),
.B(n_1),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_171),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_249),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_314),
.A2(n_329),
.B(n_356),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_157),
.B1(n_193),
.B2(n_183),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_316),
.A2(n_325),
.B1(n_354),
.B2(n_370),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_178),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_318),
.B(n_340),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_239),
.A2(n_151),
.B1(n_146),
.B2(n_175),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_327),
.A2(n_298),
.B1(n_297),
.B2(n_283),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_238),
.A2(n_299),
.B(n_262),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_333),
.B(n_237),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_242),
.B(n_145),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_346),
.Y(n_417)
);

AO22x1_ASAP7_75t_L g346 ( 
.A1(n_269),
.A2(n_194),
.B1(n_168),
.B2(n_222),
.Y(n_346)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_348),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_257),
.A2(n_228),
.B1(n_205),
.B2(n_229),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_231),
.A2(n_205),
.B1(n_229),
.B2(n_180),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_282),
.B(n_219),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_238),
.B(n_165),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_172),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_359),
.B(n_367),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_241),
.B(n_156),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_361),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_292),
.B(n_1),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_310),
.A2(n_211),
.B(n_3),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_363),
.A2(n_232),
.B(n_272),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_292),
.B(n_1),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_5),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_270),
.B(n_3),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_291),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_332),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_375),
.B(n_378),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_314),
.A2(n_245),
.B1(n_252),
.B2(n_295),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_376),
.A2(n_386),
.B1(n_398),
.B2(n_414),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_377),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_274),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_329),
.A2(n_268),
.B(n_271),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_380),
.A2(n_399),
.B(n_352),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_275),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_381),
.B(n_388),
.Y(n_441)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_354),
.A2(n_303),
.B1(n_261),
.B2(n_302),
.Y(n_386)
);

AND2x4_ASAP7_75t_SL g387 ( 
.A(n_358),
.B(n_233),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_230),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_272),
.B(n_247),
.C(n_258),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_389),
.A2(n_402),
.B(n_322),
.Y(n_442)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_344),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_401),
.Y(n_450)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_393),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_318),
.B(n_234),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_408),
.C(n_421),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_411),
.Y(n_443)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_337),
.B(n_271),
.Y(n_397)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_397),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_339),
.A2(n_309),
.B1(n_287),
.B2(n_265),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_363),
.A2(n_236),
.B(n_233),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_312),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_334),
.A2(n_255),
.B(n_235),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_403),
.A2(n_343),
.B1(n_349),
.B2(n_371),
.Y(n_426)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_406),
.B(n_366),
.Y(n_435)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_236),
.C(n_296),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_301),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_412),
.Y(n_451)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_415),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_354),
.A2(n_306),
.B1(n_273),
.B2(n_260),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_344),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_333),
.A2(n_266),
.B1(n_254),
.B2(n_259),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_416),
.A2(n_346),
.B1(n_316),
.B2(n_371),
.Y(n_459)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_319),
.Y(n_427)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_319),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_420),
.A2(n_319),
.B1(n_332),
.B2(n_362),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_290),
.C(n_256),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_322),
.B(n_253),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_424),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_253),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_375),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_425),
.B(n_437),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_426),
.A2(n_429),
.B1(n_461),
.B2(n_432),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

OAI22xp33_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_415),
.B1(n_382),
.B2(n_418),
.Y(n_429)
);

AO22x1_ASAP7_75t_L g432 ( 
.A1(n_414),
.A2(n_341),
.B1(n_337),
.B2(n_346),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_432),
.A2(n_387),
.B(n_416),
.C(n_398),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_379),
.B(n_337),
.C(n_324),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_448),
.C(n_452),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_411),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_391),
.B(n_394),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_442),
.B(n_387),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_315),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_401),
.B(n_395),
.C(n_393),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_391),
.B(n_321),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_453),
.B(n_463),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_355),
.C(n_323),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_460),
.C(n_462),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_457),
.A2(n_458),
.B(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_323),
.C(n_364),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_417),
.A2(n_396),
.B1(n_377),
.B2(n_418),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_352),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_388),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_386),
.A2(n_349),
.B1(n_343),
.B2(n_335),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_465),
.A2(n_417),
.B1(n_380),
.B2(n_409),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_405),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_466),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_423),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_468),
.B(n_475),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_470),
.A2(n_440),
.B1(n_432),
.B2(n_439),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_455),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_477),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_472),
.A2(n_481),
.B(n_486),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_449),
.A2(n_417),
.B1(n_385),
.B2(n_421),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_473),
.A2(n_483),
.B1(n_456),
.B2(n_444),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_455),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_389),
.C(n_397),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_482),
.C(n_493),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_450),
.Y(n_479)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_480),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_428),
.B(n_389),
.C(n_397),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_376),
.B1(n_387),
.B2(n_417),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_424),
.Y(n_484)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_484),
.Y(n_521)
);

INVx6_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_485),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_449),
.A2(n_402),
.B(n_420),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_434),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_487),
.B(n_489),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_434),
.B(n_423),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_441),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_450),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_490),
.A2(n_446),
.B(n_425),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_491),
.B(n_492),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_443),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_448),
.B(n_397),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_381),
.C(n_378),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_496),
.C(n_454),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_408),
.C(n_407),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_458),
.A2(n_402),
.B(n_400),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_497),
.A2(n_505),
.B(n_446),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_443),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_500),
.Y(n_544)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_447),
.Y(n_501)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_501),
.Y(n_528)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_447),
.Y(n_502)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_406),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_467),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_442),
.A2(n_440),
.B(n_464),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_462),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_506),
.B(n_509),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_511),
.A2(n_518),
.B1(n_529),
.B2(n_530),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_512),
.B(n_525),
.C(n_531),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_513),
.A2(n_517),
.B(n_540),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_469),
.B(n_464),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_514),
.B(n_516),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_439),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_472),
.A2(n_481),
.B(n_497),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_476),
.A2(n_456),
.B1(n_444),
.B2(n_465),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_522),
.B(n_524),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_523),
.A2(n_473),
.B1(n_470),
.B2(n_487),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_496),
.B(n_430),
.C(n_453),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_490),
.A2(n_486),
.B(n_505),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_527),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_503),
.A2(n_441),
.B1(n_430),
.B2(n_459),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_476),
.A2(n_426),
.B1(n_385),
.B2(n_400),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_435),
.C(n_451),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_451),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_532),
.B(n_542),
.Y(n_566)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_503),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_535),
.Y(n_573)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_494),
.Y(n_536)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_536),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_419),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_538),
.A2(n_390),
.B(n_384),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_490),
.A2(n_431),
.B(n_400),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_498),
.A2(n_410),
.B1(n_436),
.B2(n_438),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_471),
.B1(n_479),
.B2(n_489),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_493),
.B(n_413),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_483),
.A2(n_410),
.B(n_431),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_543),
.B(n_499),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_535),
.B(n_485),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_545),
.B(n_546),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_474),
.Y(n_546)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_508),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_548),
.A2(n_549),
.B1(n_555),
.B2(n_560),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_533),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_533),
.Y(n_550)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_550),
.Y(n_587)
);

OAI32xp33_ASAP7_75t_L g551 ( 
.A1(n_537),
.A2(n_484),
.A3(n_492),
.B1(n_500),
.B2(n_477),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_574),
.Y(n_583)
);

BUFx12_ASAP7_75t_L g554 ( 
.A(n_542),
.Y(n_554)
);

INVxp33_ASAP7_75t_SL g595 ( 
.A(n_554),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_557),
.A2(n_563),
.B1(n_571),
.B2(n_383),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_515),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_561),
.A2(n_528),
.B1(n_534),
.B2(n_520),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_530),
.A2(n_474),
.B1(n_495),
.B2(n_501),
.Y(n_562)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_537),
.A2(n_491),
.B1(n_480),
.B2(n_502),
.Y(n_563)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_565),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_567),
.B(n_570),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_506),
.B(n_504),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_516),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_519),
.Y(n_569)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_519),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_544),
.A2(n_491),
.B1(n_438),
.B2(n_436),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_544),
.B(n_491),
.Y(n_572)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_491),
.Y(n_574)
);

NAND5xp2_ASAP7_75t_L g575 ( 
.A(n_513),
.B(n_517),
.C(n_510),
.D(n_527),
.E(n_543),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_575),
.A2(n_518),
.B1(n_532),
.B2(n_531),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_521),
.B(n_526),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_577),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_521),
.B(n_412),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_507),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_509),
.C(n_512),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_580),
.B(n_591),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_581),
.A2(n_590),
.B1(n_600),
.B2(n_563),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_584),
.B(n_606),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_553),
.A2(n_510),
.B(n_524),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_585),
.A2(n_586),
.B(n_589),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_553),
.A2(n_540),
.B(n_511),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_588),
.B(n_601),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_552),
.A2(n_514),
.B(n_534),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_547),
.A2(n_536),
.B1(n_526),
.B2(n_528),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_507),
.C(n_520),
.Y(n_591)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_594),
.Y(n_609)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_597),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_550),
.A2(n_335),
.B1(n_338),
.B2(n_350),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_568),
.B(n_364),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_557),
.A2(n_419),
.B1(n_345),
.B2(n_365),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_603),
.A2(n_573),
.B1(n_569),
.B2(n_549),
.Y(n_614)
);

FAx1_ASAP7_75t_SL g604 ( 
.A(n_551),
.B(n_338),
.CI(n_352),
.CON(n_604),
.SN(n_604)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_579),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_556),
.B(n_347),
.C(n_328),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_605),
.B(n_608),
.C(n_566),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_556),
.B(n_347),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_578),
.B(n_328),
.C(n_362),
.Y(n_608)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_581),
.Y(n_610)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_610),
.Y(n_637)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_611),
.Y(n_643)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_598),
.Y(n_612)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_612),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_614),
.A2(n_621),
.B1(n_629),
.B2(n_597),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_615),
.B(n_617),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_616),
.B(n_625),
.Y(n_640)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_602),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_582),
.B(n_548),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_618),
.B(n_620),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_593),
.A2(n_552),
.B1(n_571),
.B2(n_573),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_587),
.A2(n_573),
.B1(n_575),
.B2(n_572),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_594),
.B(n_578),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_599),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_626),
.B(n_627),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_566),
.C(n_559),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_591),
.B(n_559),
.C(n_574),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_628),
.B(n_616),
.C(n_631),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_583),
.A2(n_607),
.B1(n_589),
.B2(n_588),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_606),
.B(n_576),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_630),
.B(n_631),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_605),
.B(n_554),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_585),
.A2(n_564),
.B(n_567),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_632),
.A2(n_586),
.B(n_592),
.Y(n_634)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_633),
.Y(n_645)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_613),
.A2(n_623),
.B(n_632),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_635),
.A2(n_621),
.B(n_630),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_636),
.B(n_644),
.Y(n_656)
);

MAJx2_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_595),
.C(n_584),
.Y(n_639)
);

XNOR2x1_ASAP7_75t_L g670 ( 
.A(n_639),
.B(n_652),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_641),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_625),
.B(n_580),
.C(n_601),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_624),
.B(n_592),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_647),
.B(n_317),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_609),
.B(n_603),
.C(n_596),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_648),
.B(n_649),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_609),
.B(n_600),
.C(n_554),
.Y(n_649)
);

MAJx2_ASAP7_75t_L g652 ( 
.A(n_629),
.B(n_604),
.C(n_570),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_627),
.B(n_622),
.C(n_624),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_653),
.B(n_336),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_SL g654 ( 
.A(n_622),
.B(n_623),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_SL g659 ( 
.A(n_654),
.B(n_619),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_643),
.A2(n_619),
.B1(n_633),
.B2(n_615),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_662),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_658),
.A2(n_649),
.B(n_647),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_659),
.B(n_660),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_636),
.B(n_614),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_651),
.B(n_604),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_661),
.B(n_664),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_646),
.A2(n_567),
.B(n_313),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g664 ( 
.A(n_651),
.B(n_336),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_665),
.B(n_667),
.Y(n_685)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_639),
.B(n_342),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_666),
.B(n_672),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_640),
.B(n_365),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_640),
.B(n_345),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_668),
.B(n_669),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_644),
.B(n_342),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_660),
.B(n_656),
.C(n_663),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_674),
.B(n_679),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_655),
.A2(n_637),
.B1(n_642),
.B2(n_641),
.Y(n_675)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_675),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_671),
.A2(n_638),
.B1(n_645),
.B2(n_648),
.Y(n_678)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_678),
.Y(n_693)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_670),
.B(n_653),
.C(n_645),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_681),
.A2(n_666),
.B(n_652),
.Y(n_687)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_659),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_683),
.B(n_661),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_670),
.B(n_650),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_684),
.A2(n_672),
.B(n_664),
.Y(n_688)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_686),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_687),
.B(n_692),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_688),
.A2(n_691),
.B(n_695),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_SL g691 ( 
.A1(n_680),
.A2(n_654),
.B(n_317),
.Y(n_691)
);

XNOR2xp5_ASAP7_75t_L g692 ( 
.A(n_674),
.B(n_374),
.Y(n_692)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_679),
.B(n_374),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_694),
.B(n_676),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_681),
.A2(n_313),
.B(n_369),
.Y(n_695)
);

MAJIxp5_ASAP7_75t_L g702 ( 
.A(n_696),
.B(n_686),
.C(n_690),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_689),
.B(n_676),
.Y(n_699)
);

AOI21xp33_ASAP7_75t_L g704 ( 
.A1(n_699),
.A2(n_701),
.B(n_697),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_693),
.A2(n_682),
.B(n_685),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_SL g705 ( 
.A1(n_702),
.A2(n_703),
.B(n_704),
.Y(n_705)
);

MAJIxp5_ASAP7_75t_L g703 ( 
.A(n_698),
.B(n_682),
.C(n_673),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_SL g706 ( 
.A1(n_704),
.A2(n_700),
.B(n_677),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_706),
.A2(n_248),
.B1(n_244),
.B2(n_285),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_707),
.B(n_705),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_SL g709 ( 
.A1(n_708),
.A2(n_369),
.B(n_330),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_SL g710 ( 
.A1(n_709),
.A2(n_369),
.B(n_7),
.C(n_8),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_SL g711 ( 
.A1(n_710),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_711)
);


endmodule