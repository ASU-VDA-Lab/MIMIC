module real_jpeg_10264_n_16 (n_5, n_4, n_8, n_0, n_12, n_325, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_325;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_1),
.A2(n_36),
.B1(n_49),
.B2(n_52),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_1),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_49),
.B1(n_52),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_3),
.A2(n_33),
.B1(n_49),
.B2(n_52),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_3),
.A2(n_33),
.B1(n_66),
.B2(n_67),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_5),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_5),
.A2(n_49),
.B1(n_52),
.B2(n_163),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_163),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_163),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_49),
.B1(n_52),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_172),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_172),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_172),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_13),
.A2(n_52),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_13),
.B(n_52),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_13),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_90),
.B1(n_93),
.B2(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_13),
.B(n_105),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_25),
.B(n_27),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_181),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_14),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_66),
.B1(n_67),
.B2(n_145),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_14),
.A2(n_49),
.B1(n_52),
.B2(n_145),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_145),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_15),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_15),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_106),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_86),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_21),
.A2(n_74),
.B1(n_75),
.B2(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_21),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_22),
.A2(n_23),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_23),
.B(n_60),
.C(n_73),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_29),
.B(n_32),
.C(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_24),
.A2(n_38),
.B1(n_264),
.B2(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_24),
.A2(n_38),
.B1(n_144),
.B2(n_273),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_45),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g206 ( 
.A(n_27),
.B(n_181),
.CON(n_206),
.SN(n_206)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_29),
.A2(n_32),
.B(n_181),
.C(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_35),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_37),
.A2(n_105),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_38),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_38),
.A2(n_144),
.B(n_146),
.Y(n_143)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_60),
.B1(n_61),
.B2(n_73),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_53),
.B(n_56),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_43),
.A2(n_59),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_43),
.A2(n_59),
.B1(n_224),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_43),
.A2(n_115),
.B(n_260),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_48),
.B1(n_54),
.B2(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_44),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_44),
.A2(n_48),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_44),
.A2(n_57),
.B(n_116),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_45),
.B(n_52),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_47),
.A2(n_49),
.B1(n_206),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_48),
.B(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_63),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_59),
.A2(n_78),
.B(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_59),
.B(n_181),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_61),
.B1(n_114),
.B2(n_119),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_70),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_62),
.A2(n_65),
.B1(n_97),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_62),
.A2(n_65),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_62),
.A2(n_65),
.B1(n_171),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_62),
.A2(n_65),
.B1(n_196),
.B2(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_62),
.A2(n_80),
.B(n_204),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_65),
.B(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_65),
.A2(n_82),
.B(n_141),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_66),
.B(n_69),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_66),
.B(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_67),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_71),
.A2(n_85),
.B(n_99),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_100),
.B(n_101),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_88),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_100),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_89),
.A2(n_96),
.B1(n_100),
.B2(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_94),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_90),
.A2(n_93),
.B1(n_162),
.B2(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_90),
.A2(n_139),
.B(n_165),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_90),
.A2(n_94),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_90),
.A2(n_93),
.B1(n_228),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_90),
.A2(n_214),
.B(n_250),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_91),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_91),
.A2(n_92),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_92),
.B(n_138),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_93),
.B(n_181),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_93),
.A2(n_137),
.B(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_96),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_103),
.B(n_105),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_121),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_120),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_152),
.B(n_323),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_149),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_125),
.B(n_149),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_133),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_315)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_133),
.A2(n_134),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.C(n_147),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_135),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_136),
.B(n_140),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI321xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_299),
.A3(n_311),
.B1(n_316),
.B2(n_322),
.C(n_325),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_266),
.C(n_295),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_240),
.B(n_265),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_217),
.B(n_239),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_199),
.B(n_216),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_190),
.B(n_198),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_178),
.B(n_189),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_166),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_173),
.B2(n_177),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_177),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_173),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_188),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_200),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.CI(n_197),
.CON(n_193),
.SN(n_193)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_210),
.B2(n_215),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_209),
.C(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_218),
.B(n_219),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_233),
.B2(n_234),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_236),
.C(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_232),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_222),
.Y(n_232)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_242),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_254),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_253),
.C(n_254),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_249),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_258),
.C(n_261),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_282),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_282),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_276),
.C(n_280),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_271),
.C(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_274),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_291),
.C(n_292),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_287),
.C(n_290),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_300),
.A2(n_317),
.B(n_321),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_301),
.B(n_302),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_308),
.C(n_310),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B(n_320),
.Y(n_317)
);


endmodule