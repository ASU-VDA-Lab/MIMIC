module fake_jpeg_104_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_18),
.Y(n_19)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_18),
.B(n_14),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_20),
.C(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_12),
.B1(n_7),
.B2(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_24),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_25),
.B(n_32),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B(n_26),
.Y(n_36)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_34),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_10),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_39),
.A3(n_10),
.B1(n_12),
.B2(n_7),
.C1(n_3),
.C2(n_2),
.Y(n_41)
);

OAI221xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_42)
);


endmodule