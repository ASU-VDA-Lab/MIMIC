module fake_aes_792_n_662 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_662);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_662;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_75), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_53), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_32), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_73), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_66), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_5), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_6), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_46), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_61), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_47), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_31), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_56), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_23), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_24), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_18), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_37), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_48), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_39), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_2), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_34), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_68), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_14), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_3), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_74), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_44), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_35), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_51), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_11), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_36), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_54), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_29), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_20), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_3), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_18), .B(n_26), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_43), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_63), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_42), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_33), .Y(n_123) );
NOR2xp67_ASAP7_75t_L g124 ( .A(n_97), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_103), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_95), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_77), .B(n_0), .Y(n_129) );
BUFx8_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_95), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_111), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_115), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_81), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_99), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_78), .B(n_1), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_88), .A2(n_76), .B(n_72), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_100), .B(n_1), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_99), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_81), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_109), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_82), .B(n_2), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_86), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_109), .B(n_4), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_118), .B(n_4), .Y(n_157) );
NOR2xp33_ASAP7_75t_R g158 ( .A(n_86), .B(n_27), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_110), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_110), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_79), .B(n_106), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_122), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_122), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_163), .B(n_92), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_163), .B(n_101), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_125), .B(n_80), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_125), .B(n_107), .Y(n_172) );
INVx8_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_148), .B(n_82), .Y(n_174) );
INVx8_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_124), .B(n_83), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_127), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_124), .B(n_83), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_143), .B(n_96), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
INVx4_ASAP7_75t_SL g182 ( .A(n_143), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_156), .B(n_92), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_133), .B(n_112), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_161), .B(n_90), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_133), .B(n_113), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
INVx6_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_157), .B(n_117), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_128), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_136), .B(n_108), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_136), .B(n_98), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_142), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_137), .B(n_102), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_131), .Y(n_206) );
AOI22x1_ASAP7_75t_L g207 ( .A1(n_137), .A2(n_121), .B1(n_96), .B2(n_114), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_141), .A2(n_105), .B1(n_104), .B2(n_121), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_141), .B(n_116), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_144), .B(n_120), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_132), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_134), .B(n_123), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_166), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_147), .A2(n_89), .B1(n_119), .B2(n_8), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_145), .B(n_52), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_135), .B(n_6), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_146), .B(n_55), .Y(n_221) );
AND2x4_ASAP7_75t_SL g222 ( .A(n_153), .B(n_7), .Y(n_222) );
NOR2x1p5_ASAP7_75t_L g223 ( .A(n_126), .B(n_7), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_212), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
INVx5_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_212), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_167), .B(n_149), .Y(n_229) );
NOR3xp33_ASAP7_75t_SL g230 ( .A(n_168), .B(n_129), .C(n_140), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_180), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_167), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_167), .A2(n_164), .B1(n_160), .B2(n_146), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_178), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_180), .A2(n_160), .B1(n_149), .B2(n_152), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_168), .B(n_152), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_214), .A2(n_142), .B(n_151), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_183), .B(n_169), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_206), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_176), .B(n_130), .Y(n_242) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_180), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_185), .B(n_158), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_173), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_185), .B(n_130), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_194), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_190), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_181), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_185), .B(n_130), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_204), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_211), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_187), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_204), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_183), .A2(n_159), .B1(n_9), .B2(n_10), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_183), .B(n_8), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_217), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_187), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_208), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_191), .B(n_159), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_177), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_191), .B(n_9), .Y(n_266) );
BUFx12f_ASAP7_75t_L g267 ( .A(n_216), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_208), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_191), .B(n_10), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_182), .B(n_11), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_177), .B(n_12), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_215), .B(n_38), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_188), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_209), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_210), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_177), .B(n_13), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_179), .A2(n_174), .B1(n_172), .B2(n_170), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_182), .B(n_14), .Y(n_280) );
NOR3xp33_ASAP7_75t_SL g281 ( .A(n_170), .B(n_15), .C(n_16), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_172), .B(n_15), .C(n_16), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_179), .B(n_17), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_187), .Y(n_284) );
AO22x1_ASAP7_75t_L g285 ( .A1(n_179), .A2(n_17), .B1(n_19), .B2(n_20), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_245), .B(n_173), .Y(n_286) );
AND2x6_ASAP7_75t_L g287 ( .A(n_271), .B(n_182), .Y(n_287) );
BUFx4f_ASAP7_75t_L g288 ( .A(n_271), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_228), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_275), .B(n_222), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_234), .B(n_173), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_245), .A2(n_175), .B1(n_218), .B2(n_197), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_275), .A2(n_198), .B(n_201), .C(n_221), .Y(n_293) );
INVx2_ASAP7_75t_SL g294 ( .A(n_271), .Y(n_294) );
AO22x1_ASAP7_75t_L g295 ( .A1(n_262), .A2(n_202), .B1(n_200), .B2(n_221), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_274), .B(n_222), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_229), .B(n_186), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_229), .B(n_213), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_255), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_243), .A2(n_175), .B1(n_198), .B2(n_201), .Y(n_300) );
AOI21x1_ASAP7_75t_SL g301 ( .A1(n_264), .A2(n_220), .B(n_202), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_228), .Y(n_302) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_227), .B(n_175), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_255), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_232), .B(n_223), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_236), .B(n_219), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_238), .B(n_219), .Y(n_308) );
INVx3_ASAP7_75t_SL g309 ( .A(n_253), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_238), .B(n_202), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_255), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_267), .Y(n_312) );
CKINVDCx8_ASAP7_75t_R g313 ( .A(n_231), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_224), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_268), .A2(n_200), .B1(n_193), .B2(n_205), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_269), .A2(n_205), .B(n_184), .C(n_193), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_243), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_255), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_233), .B(n_200), .Y(n_319) );
AOI21xp33_ASAP7_75t_SL g320 ( .A1(n_239), .A2(n_19), .B(n_21), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_247), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_225), .Y(n_322) );
BUFx12f_ASAP7_75t_L g323 ( .A(n_267), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_261), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_261), .Y(n_326) );
AND2x4_ASAP7_75t_SL g327 ( .A(n_259), .B(n_196), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_227), .B(n_196), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_261), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_259), .A2(n_184), .B1(n_192), .B2(n_189), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_227), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_270), .A2(n_203), .B1(n_192), .B2(n_189), .Y(n_332) );
AO32x2_ASAP7_75t_L g333 ( .A1(n_253), .A2(n_21), .A3(n_22), .B1(n_23), .B2(n_28), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_265), .B(n_22), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_248), .Y(n_335) );
CKINVDCx8_ASAP7_75t_R g336 ( .A(n_231), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_288), .B(n_270), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_288), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_288), .B(n_256), .Y(n_339) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_293), .A2(n_237), .B(n_263), .Y(n_340) );
OA21x2_ASAP7_75t_L g341 ( .A1(n_319), .A2(n_263), .B(n_281), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_295), .A2(n_284), .B(n_261), .Y(n_342) );
AO21x2_ASAP7_75t_L g343 ( .A1(n_320), .A2(n_258), .B(n_282), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_294), .A2(n_235), .B1(n_241), .B2(n_240), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_292), .A2(n_279), .B1(n_230), .B2(n_285), .C(n_265), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_323), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_294), .B(n_241), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_307), .A2(n_240), .B1(n_257), .B2(n_251), .Y(n_348) );
NOR2xp67_ASAP7_75t_L g349 ( .A(n_322), .B(n_280), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_321), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_287), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_321), .A2(n_266), .B1(n_283), .B2(n_272), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_310), .A2(n_265), .B1(n_280), .B2(n_242), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_295), .B(n_278), .C(n_261), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_310), .A2(n_244), .B1(n_260), .B2(n_252), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_310), .A2(n_246), .B1(n_284), .B2(n_254), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_290), .A2(n_284), .B1(n_273), .B2(n_277), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_335), .B(n_284), .Y(n_358) );
AOI221x1_ASAP7_75t_L g359 ( .A1(n_308), .A2(n_284), .B1(n_276), .B2(n_277), .C(n_171), .Y(n_359) );
INVx4_ASAP7_75t_L g360 ( .A(n_287), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_335), .A2(n_285), .B1(n_227), .B2(n_225), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_334), .B(n_225), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_323), .Y(n_363) );
INVx8_ASAP7_75t_L g364 ( .A(n_287), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_314), .B(n_250), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_290), .A2(n_276), .B1(n_250), .B2(n_226), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_298), .A2(n_226), .B1(n_249), .B2(n_225), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_287), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_345), .A2(n_296), .B1(n_300), .B2(n_334), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_337), .B(n_291), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_345), .A2(n_296), .B1(n_334), .B2(n_298), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_305), .B1(n_287), .B2(n_286), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_364), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_355), .A2(n_291), .B(n_297), .C(n_330), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_350), .B(n_314), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_365), .B(n_302), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_363), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_342), .A2(n_303), .B(n_311), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_364), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_346), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_341), .A2(n_287), .B1(n_327), .B2(n_309), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_303), .B1(n_309), .B2(n_327), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_364), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_354), .B(n_315), .C(n_332), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_365), .B(n_289), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_SL g387 ( .A1(n_367), .A2(n_324), .B(n_326), .C(n_329), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_341), .A2(n_289), .B1(n_302), .B2(n_306), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_312), .B1(n_317), .B2(n_306), .C(n_316), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_339), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_337), .B(n_326), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_340), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_348), .A2(n_336), .B1(n_313), .B2(n_325), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_370), .B(n_341), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_L g398 ( .A1(n_396), .A2(n_361), .B(n_352), .C(n_360), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_395), .A2(n_354), .B(n_342), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_371), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_371), .B(n_368), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_396), .A2(n_361), .B(n_362), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_373), .B(n_341), .C(n_359), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_391), .B(n_388), .C(n_382), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_372), .A2(n_353), .B1(n_366), .B2(n_357), .C(n_338), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_369), .A2(n_343), .B1(n_338), .B2(n_344), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_383), .B(n_349), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_371), .B(n_333), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_391), .A2(n_343), .B1(n_344), .B2(n_364), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_390), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_389), .B(n_343), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_392), .A2(n_343), .B1(n_364), .B2(n_362), .Y(n_415) );
NOR2xp33_ASAP7_75t_R g416 ( .A(n_381), .B(n_312), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_376), .Y(n_417) );
INVx3_ASAP7_75t_SL g418 ( .A(n_384), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_375), .B(n_359), .C(n_340), .Y(n_419) );
NAND2xp33_ASAP7_75t_SL g420 ( .A(n_374), .B(n_368), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_376), .B(n_333), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_392), .B(n_356), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_390), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_394), .B(n_349), .C(n_317), .D(n_333), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_377), .A2(n_362), .B1(n_360), .B2(n_368), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_378), .A2(n_362), .B1(n_336), .B2(n_313), .C(n_347), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_374), .B(n_368), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_414), .B(n_395), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_401), .B(n_333), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_414), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_411), .B(n_394), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_427), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_429), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_417), .B(n_333), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_427), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_412), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_416), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g443 ( .A1(n_428), .A2(n_393), .A3(n_385), .B(n_351), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_409), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_417), .B(n_393), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_413), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_402), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_429), .B(n_386), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_421), .B(n_386), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_411), .A2(n_385), .B1(n_364), .B2(n_351), .C1(n_380), .C2(n_360), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_387), .B1(n_362), .B2(n_380), .C(n_379), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_423), .B(n_340), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_425), .B(n_360), .C(n_328), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_410), .B(n_351), .C(n_324), .D(n_326), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_423), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_421), .B(n_340), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_400), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_400), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_397), .B(n_340), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_425), .B(n_329), .C(n_324), .Y(n_462) );
AOI21xp33_ASAP7_75t_L g463 ( .A1(n_419), .A2(n_322), .B(n_299), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_420), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_408), .A2(n_347), .B(n_329), .C(n_299), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_400), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_402), .B(n_374), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_422), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_402), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_430), .B(n_374), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_407), .B(n_318), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_399), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_418), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_418), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_399), .Y(n_476) );
OAI31xp33_ASAP7_75t_SL g477 ( .A1(n_426), .A2(n_318), .A3(n_311), .B(n_304), .Y(n_477) );
NAND2xp33_ASAP7_75t_R g478 ( .A(n_471), .B(n_430), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_433), .B(n_405), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
CKINVDCx8_ASAP7_75t_R g482 ( .A(n_464), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_442), .B(n_418), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_434), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_433), .B(n_405), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
NAND2xp33_ASAP7_75t_L g489 ( .A(n_474), .B(n_399), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_475), .B(n_430), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_468), .B(n_415), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_445), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g495 ( .A1(n_446), .A2(n_430), .A3(n_398), .B1(n_304), .B2(n_403), .B3(n_404), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_457), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_458), .B(n_404), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_446), .B(n_424), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_431), .B(n_424), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_458), .B(n_424), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_440), .B(n_424), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_454), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_450), .B(n_424), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_440), .B(n_399), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_435), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_441), .Y(n_509) );
AND2x2_ASAP7_75t_SL g510 ( .A(n_477), .B(n_399), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_444), .B(n_30), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_450), .B(n_322), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_444), .B(n_40), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_456), .B(n_331), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_461), .B(n_45), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_49), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_469), .B(n_50), .Y(n_518) );
AND2x4_ASAP7_75t_SL g519 ( .A(n_471), .B(n_325), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_449), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_467), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_469), .B(n_58), .Y(n_523) );
AND2x2_ASAP7_75t_SL g524 ( .A(n_455), .B(n_325), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_448), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_467), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_438), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_438), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_432), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_435), .B(n_322), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_432), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_470), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_521), .B(n_460), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_520), .B(n_470), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_510), .A2(n_465), .B(n_452), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_481), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_487), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_483), .B(n_462), .C(n_463), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_500), .B(n_460), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_500), .B(n_459), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_479), .A2(n_459), .B1(n_466), .B2(n_472), .C(n_443), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_503), .B(n_466), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
NAND4xp25_ASAP7_75t_L g549 ( .A(n_480), .B(n_451), .C(n_453), .D(n_471), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_492), .A2(n_473), .B1(n_476), .B2(n_453), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_490), .Y(n_553) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_515), .A2(n_473), .B(n_476), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_482), .A2(n_347), .B1(n_322), .B2(n_325), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_503), .B(n_59), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_524), .A2(n_331), .B1(n_325), .B2(n_301), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_527), .B(n_64), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
AOI21xp33_ASAP7_75t_L g560 ( .A1(n_480), .A2(n_65), .B(n_69), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_527), .B(n_70), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_508), .B(n_71), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_493), .Y(n_563) );
OAI31xp33_ASAP7_75t_L g564 ( .A1(n_486), .A2(n_227), .A3(n_249), .B(n_225), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_482), .A2(n_249), .B1(n_189), .B2(n_192), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_524), .A2(n_249), .B(n_189), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_519), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_509), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_489), .A2(n_249), .B(n_192), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g570 ( .A1(n_516), .A2(n_171), .B(n_203), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_528), .B(n_171), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_486), .B(n_171), .C(n_203), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_495), .A2(n_203), .B(n_491), .C(n_525), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_525), .B(n_514), .Y(n_574) );
AOI211x1_ASAP7_75t_L g575 ( .A1(n_528), .A2(n_530), .B(n_512), .C(n_501), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_529), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_529), .B(n_531), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_493), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_531), .B(n_507), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_494), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_573), .B(n_497), .C(n_511), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_554), .A2(n_519), .B(n_517), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_543), .B(n_497), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_575), .B(n_532), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_577), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_533), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_543), .B(n_504), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_567), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_555), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_577), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_576), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_535), .A2(n_517), .B(n_516), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_579), .B(n_504), .Y(n_594) );
AOI322xp5_ASAP7_75t_L g595 ( .A1(n_576), .A2(n_513), .A3(n_511), .B1(n_514), .B2(n_506), .C1(n_499), .C2(n_498), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_537), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_534), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_549), .A2(n_499), .B1(n_494), .B2(n_496), .C(n_498), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_537), .Y(n_599) );
NOR3xp33_ASAP7_75t_SL g600 ( .A(n_545), .B(n_478), .C(n_496), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_536), .Y(n_601) );
NOR3xp33_ASAP7_75t_SL g602 ( .A(n_565), .B(n_505), .C(n_522), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_544), .B(n_505), .Y(n_603) );
OAI211xp5_ASAP7_75t_L g604 ( .A1(n_551), .A2(n_502), .B(n_523), .C(n_518), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_551), .A2(n_502), .B(n_518), .C(n_523), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_551), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_536), .Y(n_607) );
XNOR2xp5_ASAP7_75t_L g608 ( .A(n_544), .B(n_522), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_574), .B(n_509), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_546), .B(n_538), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_539), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_546), .B(n_538), .Y(n_612) );
NOR3xp33_ASAP7_75t_L g613 ( .A(n_598), .B(n_560), .C(n_562), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_600), .A2(n_592), .B1(n_581), .B2(n_584), .C(n_589), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_601), .Y(n_615) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_609), .B(n_572), .Y(n_616) );
AOI221x1_ASAP7_75t_L g617 ( .A1(n_582), .A2(n_542), .B1(n_566), .B2(n_569), .C(n_556), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_588), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_588), .Y(n_619) );
BUFx3_ASAP7_75t_L g620 ( .A(n_583), .Y(n_620) );
AOI21xp33_ASAP7_75t_R g621 ( .A1(n_597), .A2(n_580), .B(n_563), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_607), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_609), .A2(n_570), .B(n_556), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_589), .B(n_552), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_602), .A2(n_553), .B(n_550), .Y(n_625) );
AO22x2_ASAP7_75t_L g626 ( .A1(n_606), .A2(n_541), .B1(n_547), .B2(n_548), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_604), .A2(n_561), .B1(n_558), .B2(n_547), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_611), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_606), .A2(n_561), .B1(n_558), .B2(n_548), .Y(n_629) );
INVx5_ASAP7_75t_L g630 ( .A(n_586), .Y(n_630) );
NOR4xp25_ASAP7_75t_L g631 ( .A(n_586), .B(n_580), .C(n_563), .D(n_578), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_618), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_614), .A2(n_605), .B(n_608), .C(n_583), .Y(n_633) );
NOR2x1_ASAP7_75t_R g634 ( .A(n_618), .B(n_591), .Y(n_634) );
AOI211x1_ASAP7_75t_SL g635 ( .A1(n_624), .A2(n_603), .B(n_587), .C(n_599), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_630), .B(n_612), .Y(n_636) );
NOR2xp33_ASAP7_75t_R g637 ( .A(n_619), .B(n_585), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_625), .A2(n_593), .B(n_590), .C(n_564), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_630), .Y(n_639) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_616), .B(n_599), .Y(n_640) );
NOR2xp33_ASAP7_75t_R g641 ( .A(n_620), .B(n_630), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_617), .B(n_595), .C(n_557), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_631), .A2(n_594), .B1(n_610), .B2(n_596), .C(n_540), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_626), .B(n_571), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g645 ( .A1(n_625), .A2(n_571), .B(n_559), .C(n_568), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_627), .Y(n_646) );
OAI222xp33_ASAP7_75t_L g647 ( .A1(n_629), .A2(n_559), .B1(n_568), .B2(n_623), .C1(n_621), .C2(n_615), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_626), .B(n_622), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_628), .A2(n_614), .B1(n_630), .B2(n_589), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_613), .A2(n_625), .B(n_631), .Y(n_650) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_647), .B(n_642), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g652 ( .A(n_650), .B(n_633), .C(n_635), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_649), .A2(n_646), .B1(n_632), .B2(n_643), .C1(n_648), .C2(n_639), .Y(n_653) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_633), .A2(n_638), .B(n_640), .C(n_645), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_651), .B(n_636), .Y(n_655) );
NAND4xp75_ASAP7_75t_L g656 ( .A(n_652), .B(n_641), .C(n_634), .D(n_637), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_654), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_657), .Y(n_658) );
BUFx2_ASAP7_75t_L g659 ( .A(n_655), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_659), .Y(n_660) );
AOI22xp5_ASAP7_75t_SL g661 ( .A1(n_660), .A2(n_658), .B1(n_656), .B2(n_655), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_653), .B(n_644), .Y(n_662) );
endmodule