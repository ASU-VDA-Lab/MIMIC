module fake_jpeg_18405_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_2),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_10),
.B(n_1),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_7),
.B(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_10),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_8),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_21),
.C(n_12),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_23),
.B(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_8),
.B1(n_0),
.B2(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_27),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_4),
.B(n_9),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_9),
.C(n_11),
.Y(n_35)
);

OAI211xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_9),
.C(n_11),
.Y(n_37)
);


endmodule