module fake_jpeg_3593_n_119 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_26),
.Y(n_27)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_38),
.B(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_25),
.B1(n_26),
.B2(n_14),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_13),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_58),
.B1(n_41),
.B2(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_15),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_30),
.A2(n_14),
.B1(n_25),
.B2(n_1),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_67),
.B1(n_60),
.B2(n_62),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_2),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_78),
.C(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_86),
.Y(n_87)
);

OAI22x1_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_44),
.B1(n_43),
.B2(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_67),
.B1(n_53),
.B2(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_54),
.C(n_70),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_80),
.C(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_63),
.B(n_71),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_76),
.B(n_81),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_77),
.B(n_80),
.C(n_76),
.D(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_94),
.C(n_87),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_108),
.C(n_109),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_92),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_100),
.Y(n_112)
);

AOI211xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_98),
.B(n_105),
.C(n_106),
.Y(n_113)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_72),
.B(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_114),
.B1(n_56),
.B2(n_11),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_10),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_10),
.Y(n_119)
);


endmodule