module fake_netlist_5_2149_n_1038 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1038);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1038;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_443;
wire n_293;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_679;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_985;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_144),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_90),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_6),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_5),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_74),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_131),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_146),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_139),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_37),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_16),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_150),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_8),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_44),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_161),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_38),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_87),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_54),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_21),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_205),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_133),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_46),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_121),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_171),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_31),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_142),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_111),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_65),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_27),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_13),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_36),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_30),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_93),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_62),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_22),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_42),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_98),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_14),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_47),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_211),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_221),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_55),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_154),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_9),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_180),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_89),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_64),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_1),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_40),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_203),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_100),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_109),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_12),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_129),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_99),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_155),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_200),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_189),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_175),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_72),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_102),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_132),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_33),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_183),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_149),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_124),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_78),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_170),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_192),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_230),
.Y(n_320)
);

BUFx6f_ASAP7_75t_SL g321 ( 
.A(n_244),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_254),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_230),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_224),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_226),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_228),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_232),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_242),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_233),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_234),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_227),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_262),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_242),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_251),
.B(n_0),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_250),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_239),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_227),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_262),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_250),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_243),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_248),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_241),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_288),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_269),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_270),
.B(n_1),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_249),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_252),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_240),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_255),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_241),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_260),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_257),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_261),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_263),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_251),
.B(n_260),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_253),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_225),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_264),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_253),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_333),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_326),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_327),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_328),
.B(n_331),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_332),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_342),
.Y(n_391)
);

OA21x2_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_256),
.B(n_247),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_346),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_347),
.B(n_235),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_355),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_258),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_321),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_343),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_361),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_366),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_268),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_344),
.B(n_244),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_353),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_340),
.A2(n_277),
.B(n_275),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_281),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_374),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_321),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_338),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_338),
.B(n_282),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_343),
.B(n_282),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_348),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_368),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_414),
.A2(n_323),
.B1(n_329),
.B2(n_296),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_236),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_278),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_313),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_229),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_398),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_274),
.C(n_259),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_315),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_291),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_427),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_237),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_291),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_382),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

AND2x2_ASAP7_75t_SL g471 ( 
.A(n_419),
.B(n_295),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_400),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_432),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_400),
.B(n_300),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_407),
.B(n_246),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_265),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_380),
.B(n_308),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_309),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_379),
.B(n_272),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_424),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_428),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

AND3x2_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_318),
.C(n_310),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_385),
.B(n_273),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_389),
.B(n_231),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_380),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_419),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_395),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_SL g497 ( 
.A(n_383),
.B(n_279),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_419),
.B(n_283),
.Y(n_498)
);

NOR2x1p5_ASAP7_75t_L g499 ( 
.A(n_424),
.B(n_286),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_390),
.A2(n_271),
.B1(n_292),
.B2(n_245),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_383),
.Y(n_501)
);

INVx6_ASAP7_75t_L g502 ( 
.A(n_393),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_386),
.B(n_284),
.Y(n_503)
);

AO22x2_ASAP7_75t_L g504 ( 
.A1(n_390),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_386),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_450),
.B(n_419),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_448),
.B(n_388),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_448),
.B(n_388),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_443),
.A2(n_405),
.B(n_426),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_449),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_465),
.B(n_391),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_391),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_473),
.B(n_397),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_466),
.B(n_397),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_466),
.B(n_399),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_399),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_439),
.B(n_401),
.Y(n_522)
);

NAND2x1_ASAP7_75t_L g523 ( 
.A(n_439),
.B(n_426),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_445),
.B(n_401),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_471),
.A2(n_312),
.B1(n_293),
.B2(n_299),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_472),
.B(n_479),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_474),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_SL g529 ( 
.A(n_478),
.B(n_411),
.C(n_406),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_498),
.A2(n_289),
.B(n_285),
.Y(n_530)
);

A2O1A1Ixp33_ASAP7_75t_L g531 ( 
.A1(n_472),
.A2(n_474),
.B(n_484),
.C(n_471),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_484),
.A2(n_297),
.B(n_294),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_479),
.B(n_406),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_479),
.A2(n_411),
.B1(n_422),
.B2(n_304),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_479),
.B(n_422),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_474),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_SL g539 ( 
.A(n_497),
.B(n_306),
.C(n_425),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_479),
.B(n_302),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_454),
.B(n_461),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_461),
.B(n_303),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_464),
.B(n_305),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_463),
.B(n_348),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_477),
.B(n_307),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_438),
.B(n_402),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_486),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_464),
.B(n_311),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_495),
.A2(n_488),
.B1(n_478),
.B2(n_503),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_455),
.B(n_231),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_506),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_495),
.A2(n_362),
.B1(n_371),
.B2(n_375),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_492),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_488),
.A2(n_316),
.B(n_314),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_444),
.B(n_425),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_362),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_492),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_437),
.Y(n_560)
);

O2A1O1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_455),
.A2(n_371),
.B(n_375),
.C(n_320),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_503),
.B(n_244),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_489),
.B(n_266),
.Y(n_563)
);

AND2x6_ASAP7_75t_SL g564 ( 
.A(n_491),
.B(n_320),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_457),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_485),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_440),
.B(n_507),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_467),
.B(n_324),
.C(n_377),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_483),
.B(n_497),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_462),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_463),
.A2(n_324),
.B1(n_404),
.B2(n_429),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_467),
.A2(n_266),
.B1(n_106),
.B2(n_107),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_43),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_507),
.B(n_266),
.Y(n_576)
);

AND3x2_ASAP7_75t_L g577 ( 
.A(n_504),
.B(n_2),
.C(n_4),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_508),
.B(n_45),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_508),
.B(n_50),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_501),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_493),
.B(n_5),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_440),
.B(n_51),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_496),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_502),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_446),
.B(n_52),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_502),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_480),
.A2(n_113),
.B1(n_222),
.B2(n_220),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_504),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_451),
.B(n_7),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_447),
.B(n_53),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_490),
.A2(n_57),
.B(n_56),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_459),
.B(n_58),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_502),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_536),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_511),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_518),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_566),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_589),
.B(n_501),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_591),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_584),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_514),
.B(n_558),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_510),
.B(n_482),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_566),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_519),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_554),
.B(n_499),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_512),
.B(n_491),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_536),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_555),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_542),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_441),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_590),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_559),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_591),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_528),
.B(n_548),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_550),
.A2(n_460),
.B1(n_469),
.B2(n_494),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_534),
.B(n_460),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_541),
.B(n_441),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_585),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_560),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_551),
.B(n_469),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_562),
.A2(n_475),
.B1(n_494),
.B2(n_500),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_587),
.B(n_504),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_475),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_552),
.B(n_487),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_560),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_562),
.B(n_522),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_581),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_435),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_509),
.A2(n_452),
.B(n_437),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_520),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_533),
.A2(n_535),
.B1(n_520),
.B2(n_529),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_538),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_575),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_553),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_577),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_565),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_578),
.B(n_500),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_570),
.B(n_435),
.Y(n_642)
);

O2A1O1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_531),
.A2(n_582),
.B(n_589),
.C(n_529),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_569),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_567),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_583),
.B(n_436),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_527),
.A2(n_500),
.B1(n_437),
.B2(n_452),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_574),
.B(n_487),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_564),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_573),
.B(n_516),
.Y(n_650)
);

NOR3xp33_ASAP7_75t_SL g651 ( 
.A(n_572),
.B(n_482),
.C(n_9),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_583),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_521),
.Y(n_653)
);

NAND2x1_ASAP7_75t_L g654 ( 
.A(n_579),
.B(n_437),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_517),
.B(n_458),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_526),
.B(n_436),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_513),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_609),
.B(n_526),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_633),
.A2(n_544),
.B(n_543),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_607),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

AOI221xp5_ASAP7_75t_L g664 ( 
.A1(n_643),
.A2(n_561),
.B1(n_568),
.B2(n_545),
.C(n_572),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_654),
.A2(n_580),
.B(n_586),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_646),
.A2(n_658),
.B(n_629),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_623),
.A2(n_549),
.B(n_556),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_659),
.A2(n_593),
.B(n_592),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_596),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_659),
.A2(n_523),
.B(n_540),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_620),
.A2(n_530),
.B(n_532),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_600),
.B(n_539),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_618),
.A2(n_588),
.B(n_576),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_645),
.A2(n_547),
.B(n_563),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_600),
.A2(n_453),
.B(n_452),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_599),
.A2(n_563),
.B(n_539),
.C(n_557),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_606),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_626),
.A2(n_622),
.B(n_613),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_628),
.A2(n_453),
.B(n_452),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_628),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_652),
.B(n_524),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_657),
.A2(n_453),
.B(n_546),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_655),
.B(n_482),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_652),
.A2(n_453),
.B1(n_481),
.B2(n_524),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_611),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_652),
.A2(n_481),
.B1(n_118),
.B2(n_119),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_631),
.A2(n_481),
.B(n_60),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_621),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_598),
.A2(n_481),
.B(n_117),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_600),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_651),
.B(n_604),
.C(n_653),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_619),
.A2(n_120),
.B(n_219),
.Y(n_693)
);

INVx3_ASAP7_75t_SL g694 ( 
.A(n_615),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_598),
.A2(n_116),
.B(n_218),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_616),
.B(n_11),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_636),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_616),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_616),
.A2(n_122),
.B(n_217),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_635),
.B(n_59),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_642),
.B(n_597),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_605),
.A2(n_115),
.B(n_213),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_640),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_601),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_605),
.A2(n_112),
.B(n_212),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_602),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_603),
.B(n_14),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_632),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_650),
.B(n_61),
.Y(n_709)
);

AOI21x1_ASAP7_75t_L g710 ( 
.A1(n_638),
.A2(n_125),
.B(n_210),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_644),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_647),
.A2(n_123),
.B(n_209),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_612),
.A2(n_110),
.B(n_208),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_637),
.A2(n_108),
.B(n_207),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_610),
.Y(n_715)
);

AOI21x1_ASAP7_75t_SL g716 ( 
.A1(n_648),
.A2(n_17),
.B(n_18),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_656),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_694),
.Y(n_718)
);

CKINVDCx11_ASAP7_75t_R g719 ( 
.A(n_694),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_663),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_L g721 ( 
.A1(n_660),
.A2(n_608),
.B1(n_614),
.B2(n_630),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_670),
.A2(n_624),
.B(n_595),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_663),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_669),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_669),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_677),
.B(n_634),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_708),
.A2(n_634),
.B1(n_632),
.B2(n_639),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_670),
.A2(n_650),
.B(n_656),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_661),
.A2(n_639),
.A3(n_650),
.B(n_625),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_717),
.B(n_625),
.Y(n_730)
);

AOI22x1_ASAP7_75t_L g731 ( 
.A1(n_666),
.A2(n_678),
.B1(n_667),
.B2(n_693),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_662),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_704),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_717),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_683),
.A2(n_650),
.B(n_648),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_686),
.B(n_649),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_706),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_697),
.Y(n_738)
);

CKINVDCx16_ASAP7_75t_R g739 ( 
.A(n_684),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_673),
.A2(n_617),
.B(n_627),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_683),
.A2(n_627),
.B(n_617),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_697),
.Y(n_742)
);

OAI21x1_ASAP7_75t_SL g743 ( 
.A1(n_710),
.A2(n_641),
.B(n_127),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_708),
.A2(n_641),
.B1(n_649),
.B2(n_621),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_676),
.A2(n_18),
.A3(n_19),
.B(n_20),
.Y(n_745)
);

AO21x2_ASAP7_75t_L g746 ( 
.A1(n_700),
.A2(n_126),
.B(n_206),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_690),
.A2(n_105),
.B(n_204),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_698),
.B(n_63),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_703),
.B(n_66),
.Y(n_749)
);

OA21x2_ASAP7_75t_L g750 ( 
.A1(n_668),
.A2(n_19),
.B(n_20),
.Y(n_750)
);

OAI21x1_ASAP7_75t_L g751 ( 
.A1(n_690),
.A2(n_134),
.B(n_201),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_703),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_686),
.Y(n_753)
);

OAI21x1_ASAP7_75t_L g754 ( 
.A1(n_665),
.A2(n_130),
.B(n_199),
.Y(n_754)
);

AO21x2_ASAP7_75t_L g755 ( 
.A1(n_700),
.A2(n_104),
.B(n_198),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_711),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_711),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_715),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_715),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_675),
.B(n_67),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_707),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_692),
.A2(n_701),
.B1(n_664),
.B2(n_696),
.Y(n_762)
);

OA21x2_ASAP7_75t_L g763 ( 
.A1(n_668),
.A2(n_712),
.B(n_713),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_682),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_679),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_676),
.B(n_21),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_672),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_665),
.A2(n_135),
.B(n_194),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_679),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_681),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_770)
);

OAI222xp33_ASAP7_75t_L g771 ( 
.A1(n_691),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C1(n_26),
.C2(n_27),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_730),
.B(n_698),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_761),
.B(n_707),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_766),
.A2(n_708),
.B1(n_682),
.B2(n_672),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_766),
.A2(n_709),
.B(n_672),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_759),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_730),
.B(n_698),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_744),
.A2(n_687),
.B1(n_685),
.B2(n_681),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_764),
.A2(n_709),
.B1(n_712),
.B2(n_674),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_759),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_739),
.B(n_689),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_733),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_762),
.A2(n_699),
.B1(n_705),
.B2(n_714),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_767),
.B(n_713),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_767),
.B(n_695),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_733),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_758),
.B(n_680),
.Y(n_787)
);

AO31x2_ASAP7_75t_L g788 ( 
.A1(n_720),
.A2(n_716),
.A3(n_671),
.B(n_688),
.Y(n_788)
);

AO31x2_ASAP7_75t_L g789 ( 
.A1(n_720),
.A2(n_671),
.A3(n_702),
.B(n_695),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_721),
.A2(n_702),
.B1(n_28),
.B2(n_29),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_727),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_737),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_739),
.B(n_34),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_732),
.B(n_34),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_731),
.A2(n_143),
.B(n_193),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_737),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_760),
.B(n_68),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_731),
.A2(n_223),
.B(n_141),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_718),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_719),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_753),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

AO22x1_ASAP7_75t_L g803 ( 
.A1(n_764),
.A2(n_753),
.B1(n_726),
.B2(n_770),
.Y(n_803)
);

CKINVDCx8_ASAP7_75t_R g804 ( 
.A(n_748),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_748),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_740),
.A2(n_191),
.B(n_140),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_734),
.B(n_756),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_746),
.A2(n_755),
.B(n_743),
.Y(n_808)
);

AND2x6_ASAP7_75t_L g809 ( 
.A(n_748),
.B(n_138),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_748),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_736),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_746),
.A2(n_35),
.B1(n_39),
.B2(n_69),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_756),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_757),
.B(n_39),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_757),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_734),
.B(n_70),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_742),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_742),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_724),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_749),
.B(n_71),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_765),
.B(n_73),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_L g822 ( 
.A(n_765),
.B(n_75),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_724),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_738),
.B(n_76),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_749),
.B(n_77),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_725),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_738),
.B(n_79),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_752),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_769),
.Y(n_830)
);

AOI221xp5_ASAP7_75t_L g831 ( 
.A1(n_811),
.A2(n_771),
.B1(n_743),
.B2(n_755),
.C(n_746),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_775),
.A2(n_755),
.B1(n_760),
.B2(n_741),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_830),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_775),
.A2(n_760),
.B1(n_741),
.B2(n_769),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_SL g835 ( 
.A1(n_774),
.A2(n_814),
.B1(n_778),
.B2(n_809),
.Y(n_835)
);

OAI33xp33_ASAP7_75t_L g836 ( 
.A1(n_792),
.A2(n_723),
.A3(n_752),
.B1(n_745),
.B2(n_729),
.B3(n_750),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_745),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_774),
.A2(n_760),
.B1(n_723),
.B2(n_735),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_782),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_806),
.A2(n_747),
.B(n_751),
.C(n_768),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_772),
.B(n_745),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_786),
.B(n_745),
.Y(n_842)
);

OAI321xp33_ASAP7_75t_L g843 ( 
.A1(n_792),
.A2(n_745),
.A3(n_729),
.B1(n_750),
.B2(n_722),
.C(n_735),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_797),
.B(n_728),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_791),
.A2(n_750),
.B1(n_722),
.B2(n_763),
.Y(n_845)
);

AOI221xp5_ASAP7_75t_L g846 ( 
.A1(n_773),
.A2(n_729),
.B1(n_750),
.B2(n_728),
.C(n_754),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_783),
.A2(n_751),
.B(n_747),
.C(n_754),
.Y(n_847)
);

AOI221xp5_ASAP7_75t_L g848 ( 
.A1(n_812),
.A2(n_729),
.B1(n_768),
.B2(n_763),
.C(n_84),
.Y(n_848)
);

AO21x2_ASAP7_75t_L g849 ( 
.A1(n_808),
.A2(n_763),
.B(n_729),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_L g850 ( 
.A1(n_797),
.A2(n_763),
.B1(n_81),
.B2(n_83),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_772),
.B(n_80),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_777),
.B(n_85),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_797),
.A2(n_190),
.B1(n_88),
.B2(n_91),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_809),
.A2(n_86),
.B1(n_92),
.B2(n_94),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_804),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_788),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_800),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_778),
.A2(n_101),
.B1(n_103),
.B2(n_136),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_809),
.A2(n_137),
.B1(n_145),
.B2(n_147),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_777),
.B(n_148),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_793),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_799),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_803),
.B(n_156),
.Y(n_863)
);

AOI221xp5_ASAP7_75t_L g864 ( 
.A1(n_790),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.C(n_160),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_809),
.A2(n_822),
.B1(n_810),
.B2(n_784),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_794),
.A2(n_188),
.B1(n_163),
.B2(n_164),
.Y(n_866)
);

OAI221xp5_ASAP7_75t_L g867 ( 
.A1(n_779),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.C(n_169),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_820),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_819),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_781),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_805),
.B(n_181),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_816),
.B(n_184),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_824),
.B(n_185),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_801),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_796),
.Y(n_875)
);

BUFx4f_ASAP7_75t_L g876 ( 
.A(n_844),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_844),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_856),
.B(n_789),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_839),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_843),
.A2(n_808),
.B(n_798),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_849),
.B(n_841),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_844),
.B(n_789),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_849),
.B(n_788),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_842),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_837),
.B(n_788),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_835),
.A2(n_795),
.B1(n_826),
.B2(n_821),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_875),
.B(n_815),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_869),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_871),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_846),
.B(n_776),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_838),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_862),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_873),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_853),
.A2(n_802),
.B1(n_799),
.B2(n_813),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_871),
.Y(n_895)
);

NOR2x1_ASAP7_75t_L g896 ( 
.A(n_850),
.B(n_780),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_832),
.B(n_845),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_833),
.Y(n_898)
);

NOR2x1_ASAP7_75t_SL g899 ( 
.A(n_863),
.B(n_785),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_845),
.B(n_817),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_847),
.B(n_818),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_840),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_834),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_860),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_848),
.B(n_829),
.Y(n_905)
);

BUFx12f_ASAP7_75t_L g906 ( 
.A(n_857),
.Y(n_906)
);

INVxp67_ASAP7_75t_SL g907 ( 
.A(n_836),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_831),
.B(n_823),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_865),
.B(n_823),
.Y(n_909)
);

OAI31xp33_ASAP7_75t_L g910 ( 
.A1(n_894),
.A2(n_850),
.A3(n_861),
.B(n_855),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_882),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_879),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_882),
.Y(n_913)
);

NOR2x1_ASAP7_75t_SL g914 ( 
.A(n_877),
.B(n_802),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_881),
.B(n_853),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_902),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_881),
.B(n_858),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_902),
.B(n_866),
.C(n_864),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_891),
.A2(n_867),
.B1(n_855),
.B2(n_861),
.Y(n_919)
);

AOI221xp5_ASAP7_75t_L g920 ( 
.A1(n_907),
.A2(n_866),
.B1(n_870),
.B2(n_859),
.C(n_854),
.Y(n_920)
);

AOI221xp5_ASAP7_75t_L g921 ( 
.A1(n_907),
.A2(n_868),
.B1(n_872),
.B2(n_852),
.C(n_851),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_890),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_891),
.A2(n_821),
.B1(n_874),
.B2(n_828),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_897),
.A2(n_903),
.B1(n_886),
.B2(n_909),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_886),
.B(n_825),
.C(n_787),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_879),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_888),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

OAI221xp5_ASAP7_75t_L g930 ( 
.A1(n_903),
.A2(n_186),
.B1(n_827),
.B2(n_894),
.C(n_896),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_912),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_913),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_911),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_929),
.B(n_881),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_911),
.B(n_882),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_922),
.B(n_885),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_916),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_913),
.B(n_876),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_913),
.B(n_877),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_912),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_910),
.B(n_896),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_913),
.B(n_882),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_918),
.A2(n_897),
.B1(n_876),
.B2(n_909),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_915),
.B(n_882),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_928),
.Y(n_945)
);

NAND4xp25_ASAP7_75t_L g946 ( 
.A(n_941),
.B(n_910),
.C(n_918),
.D(n_919),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_931),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_933),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_941),
.B(n_906),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_944),
.B(n_898),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_936),
.B(n_915),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_936),
.B(n_926),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_944),
.B(n_898),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_950),
.B(n_935),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_948),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_947),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_951),
.B(n_937),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_953),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_952),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_898),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_949),
.Y(n_961)
);

OAI22xp33_ASAP7_75t_L g962 ( 
.A1(n_958),
.A2(n_946),
.B1(n_930),
.B2(n_925),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_956),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_959),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_961),
.A2(n_957),
.B(n_937),
.C(n_920),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_964),
.Y(n_967)
);

AOI221xp5_ASAP7_75t_L g968 ( 
.A1(n_965),
.A2(n_957),
.B1(n_955),
.B2(n_924),
.C(n_943),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_962),
.A2(n_963),
.B(n_925),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_967),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_969),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_966),
.B(n_958),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_968),
.B(n_906),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_969),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_SL g975 ( 
.A1(n_972),
.A2(n_954),
.B(n_935),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_970),
.B(n_934),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_SL g977 ( 
.A1(n_971),
.A2(n_899),
.B1(n_917),
.B2(n_914),
.Y(n_977)
);

OAI211xp5_ASAP7_75t_L g978 ( 
.A1(n_973),
.A2(n_974),
.B(n_921),
.C(n_917),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_970),
.Y(n_979)
);

INVxp33_ASAP7_75t_L g980 ( 
.A(n_972),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_971),
.B(n_934),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_970),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_980),
.B(n_933),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_979),
.A2(n_938),
.B(n_932),
.Y(n_984)
);

AOI211xp5_ASAP7_75t_L g985 ( 
.A1(n_978),
.A2(n_897),
.B(n_939),
.C(n_933),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_SL g986 ( 
.A(n_977),
.B(n_938),
.C(n_923),
.Y(n_986)
);

AOI21xp33_ASAP7_75t_L g987 ( 
.A1(n_982),
.A2(n_906),
.B(n_893),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_975),
.B(n_940),
.Y(n_988)
);

O2A1O1Ixp5_ASAP7_75t_SL g989 ( 
.A1(n_981),
.A2(n_932),
.B(n_940),
.C(n_931),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_R g990 ( 
.A(n_976),
.B(n_932),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_983),
.B(n_892),
.Y(n_991)
);

OAI221xp5_ASAP7_75t_L g992 ( 
.A1(n_985),
.A2(n_938),
.B1(n_876),
.B2(n_932),
.C(n_877),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_987),
.B(n_942),
.Y(n_993)
);

AOI33xp33_ASAP7_75t_L g994 ( 
.A1(n_990),
.A2(n_939),
.A3(n_942),
.B1(n_905),
.B2(n_893),
.B3(n_901),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_988),
.B(n_899),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_986),
.Y(n_996)
);

OAI211xp5_ASAP7_75t_L g997 ( 
.A1(n_984),
.A2(n_989),
.B(n_877),
.C(n_908),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_R g998 ( 
.A(n_983),
.B(n_892),
.Y(n_998)
);

NAND2x1_ASAP7_75t_L g999 ( 
.A(n_983),
.B(n_939),
.Y(n_999)
);

AOI211xp5_ASAP7_75t_L g1000 ( 
.A1(n_996),
.A2(n_939),
.B(n_892),
.C(n_908),
.Y(n_1000)
);

NOR2x1_ASAP7_75t_L g1001 ( 
.A(n_999),
.B(n_945),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_992),
.A2(n_876),
.B1(n_877),
.B2(n_893),
.C(n_904),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_993),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_995),
.B(n_914),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_991),
.B(n_945),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_997),
.B(n_927),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1005),
.A2(n_876),
.B1(n_892),
.B2(n_890),
.Y(n_1009)
);

NAND5xp2_ASAP7_75t_L g1010 ( 
.A(n_1000),
.B(n_905),
.C(n_885),
.D(n_900),
.E(n_883),
.Y(n_1010)
);

AND4x1_ASAP7_75t_L g1011 ( 
.A(n_1001),
.B(n_905),
.C(n_900),
.D(n_884),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_1003),
.A2(n_892),
.B1(n_904),
.B2(n_889),
.Y(n_1012)
);

NOR3x1_ASAP7_75t_SL g1013 ( 
.A(n_1004),
.B(n_892),
.C(n_904),
.Y(n_1013)
);

AOI32xp33_ASAP7_75t_L g1014 ( 
.A1(n_1007),
.A2(n_889),
.A3(n_909),
.B1(n_904),
.B2(n_901),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1008),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1006),
.Y(n_1016)
);

INVxp67_ASAP7_75t_SL g1017 ( 
.A(n_1002),
.Y(n_1017)
);

CKINVDCx16_ASAP7_75t_R g1018 ( 
.A(n_1016),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_1015),
.Y(n_1019)
);

NAND2x1_ASAP7_75t_L g1020 ( 
.A(n_1013),
.B(n_892),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_1017),
.B(n_904),
.C(n_889),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_1011),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_L g1023 ( 
.A(n_1020),
.B(n_1012),
.Y(n_1023)
);

OAI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_1021),
.A2(n_1009),
.B1(n_1014),
.B2(n_1010),
.C(n_889),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1018),
.B(n_1022),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1019),
.Y(n_1026)
);

NAND4xp25_ASAP7_75t_L g1027 ( 
.A(n_1025),
.B(n_889),
.C(n_895),
.D(n_909),
.Y(n_1027)
);

OAI211xp5_ASAP7_75t_L g1028 ( 
.A1(n_1026),
.A2(n_887),
.B(n_880),
.C(n_926),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_1027),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_1030),
.A2(n_1023),
.B(n_1024),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1029),
.B(n_888),
.Y(n_1032)
);

AOI222xp33_ASAP7_75t_L g1033 ( 
.A1(n_1032),
.A2(n_909),
.B1(n_927),
.B2(n_901),
.C1(n_895),
.C2(n_887),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_1031),
.A2(n_895),
.B1(n_880),
.B2(n_901),
.Y(n_1034)
);

AOI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_1031),
.A2(n_888),
.B(n_928),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_1035),
.A2(n_901),
.B1(n_880),
.B2(n_900),
.Y(n_1036)
);

AOI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_1036),
.A2(n_1034),
.B1(n_1033),
.B2(n_928),
.C(n_883),
.Y(n_1037)
);

AOI211xp5_ASAP7_75t_L g1038 ( 
.A1(n_1037),
.A2(n_883),
.B(n_885),
.C(n_878),
.Y(n_1038)
);


endmodule