module fake_jpeg_29782_n_366 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_366);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_366;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_16),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_59),
.Y(n_90)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_27),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_15),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_24),
.B1(n_34),
.B2(n_33),
.Y(n_115)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_94),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_41),
.B1(n_21),
.B2(n_28),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_83),
.A2(n_100),
.B1(n_101),
.B2(n_121),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_24),
.B1(n_38),
.B2(n_35),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_33),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_46),
.A2(n_41),
.B1(n_21),
.B2(n_28),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_41),
.B1(n_21),
.B2(n_28),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_142)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_29),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_25),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_35),
.B1(n_26),
.B2(n_34),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_80),
.B1(n_99),
.B2(n_77),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_4),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_7),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_55),
.A2(n_28),
.B1(n_21),
.B2(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_30),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_0),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_152),
.B1(n_162),
.B2(n_80),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_26),
.B(n_10),
.C(n_15),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_149),
.C(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_8),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_127),
.B(n_139),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_79),
.B(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_86),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_137),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_143),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_147),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_141),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_150),
.B1(n_128),
.B2(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_145),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_10),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_10),
.B(n_11),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_155),
.B1(n_105),
.B2(n_119),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_4),
.B1(n_5),
.B2(n_99),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_109),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_159),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_120),
.Y(n_159)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_5),
.A3(n_92),
.B1(n_86),
.B2(n_77),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_82),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_78),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_108),
.B(n_92),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_165),
.B(n_188),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_173),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_170),
.A2(n_171),
.B(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_119),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_189),
.B1(n_196),
.B2(n_197),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_95),
.B1(n_104),
.B2(n_137),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_176),
.A2(n_201),
.B1(n_141),
.B2(n_165),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_135),
.Y(n_178)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_178),
.A2(n_170),
.B1(n_169),
.B2(n_183),
.Y(n_223)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_95),
.A3(n_139),
.B1(n_132),
.B2(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_133),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_135),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_142),
.B(n_162),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_194),
.B(n_188),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_143),
.B(n_138),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_126),
.C(n_129),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_177),
.C(n_187),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_136),
.B1(n_154),
.B2(n_153),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_146),
.B1(n_152),
.B2(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_127),
.B(n_124),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_198),
.B(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_151),
.B1(n_148),
.B2(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_157),
.B1(n_141),
.B2(n_164),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_219),
.B(n_223),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_207),
.A2(n_209),
.B1(n_221),
.B2(n_225),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_171),
.B(n_198),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_210),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_226),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_192),
.B1(n_185),
.B2(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_227),
.B1(n_230),
.B2(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_224),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_173),
.A2(n_201),
.B1(n_193),
.B2(n_181),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_176),
.A2(n_199),
.B1(n_196),
.B2(n_194),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_166),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_174),
.B1(n_178),
.B2(n_170),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_231),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_235),
.B(n_205),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_200),
.B1(n_184),
.B2(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_172),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_236),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_202),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_179),
.A2(n_167),
.B1(n_173),
.B2(n_201),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_251),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_250),
.B(n_257),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_216),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_225),
.B1(n_236),
.B2(n_209),
.Y(n_268)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_219),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_270),
.B1(n_275),
.B2(n_287),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_218),
.C(n_206),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_274),
.C(n_281),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_217),
.B1(n_227),
.B2(n_229),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_207),
.B1(n_219),
.B2(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_231),
.C(n_207),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_258),
.B1(n_259),
.B2(n_264),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_280),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_241),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_265),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_243),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_259),
.B1(n_244),
.B2(n_250),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_289),
.B(n_305),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_251),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_295),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_240),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_296),
.A2(n_275),
.B(n_270),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_240),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_303),
.Y(n_307)
);

OAI31xp33_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_244),
.A3(n_249),
.B(n_257),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_279),
.B(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_239),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_300),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_245),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_272),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_267),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_282),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_274),
.C(n_271),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_316),
.C(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_317),
.B(n_293),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_268),
.B1(n_271),
.B2(n_267),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_295),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_282),
.B1(n_283),
.B2(n_266),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_249),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_283),
.B(n_242),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_277),
.B1(n_242),
.B2(n_246),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_277),
.B1(n_252),
.B2(n_248),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_241),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_SL g339 ( 
.A1(n_327),
.A2(n_315),
.B(n_314),
.C(n_297),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_330),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_303),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_298),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_246),
.B1(n_248),
.B2(n_262),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_304),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_316),
.B(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_327),
.B1(n_322),
.B2(n_307),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_340),
.B(n_325),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_328),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_308),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_307),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_347),
.B(n_348),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_345),
.A2(n_329),
.B(n_335),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_349),
.A2(n_345),
.B(n_339),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_352),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_330),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_329),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_351),
.A2(n_342),
.B(n_338),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_354),
.B(n_357),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_359),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_358),
.B(n_349),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_360),
.Y(n_363)
);

OAI21xp33_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_355),
.B(n_254),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_363),
.C(n_361),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_344),
.Y(n_366)
);


endmodule