module fake_jpeg_22356_n_85 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_0),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_45),
.C(n_37),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_36),
.C(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_58),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_57),
.B(n_44),
.C(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_43),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_1),
.Y(n_58)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_59),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_6),
.C(n_7),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_65),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_13),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_76),
.B1(n_74),
.B2(n_73),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_71),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_31),
.Y(n_85)
);


endmodule