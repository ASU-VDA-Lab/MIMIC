module real_jpeg_19901_n_17 (n_8, n_0, n_2, n_338, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_338;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_0),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_0),
.A2(n_70),
.B1(n_71),
.B2(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_105),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_105),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_1),
.A2(n_39),
.B1(n_70),
.B2(n_71),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_1),
.A2(n_39),
.B1(n_47),
.B2(n_49),
.Y(n_284)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_3),
.A2(n_70),
.B1(n_71),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_3),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_47),
.B1(n_49),
.B2(n_122),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_122),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_4),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_5),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_5),
.A2(n_47),
.B1(n_49),
.B2(n_63),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_63),
.Y(n_277)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_6),
.B(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_6),
.A2(n_145),
.B(n_171),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_7),
.A2(n_29),
.B1(n_70),
.B2(n_71),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_7),
.A2(n_29),
.B1(n_47),
.B2(n_49),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_9),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_70),
.B1(n_71),
.B2(n_84),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_47),
.B1(n_49),
.B2(n_84),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_84),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_49),
.B(n_66),
.C(n_102),
.D(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_10),
.B(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_10),
.B(n_46),
.Y(n_113)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_123),
.B(n_125),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_10),
.A2(n_36),
.B(n_43),
.C(n_161),
.D(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_10),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_40),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_35),
.B(n_37),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_142),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_12),
.A2(n_47),
.B1(n_49),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_12),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_70),
.B1(n_71),
.B2(n_117),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_117),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_117),
.Y(n_230)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_53),
.B1(n_54),
.B2(n_75),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_27),
.A2(n_32),
.B(n_142),
.C(n_203),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_30),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_30),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_31),
.A2(n_34),
.B1(n_62),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_31),
.A2(n_34),
.B1(n_230),
.B2(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_31),
.A2(n_221),
.B(n_261),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_34),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_34),
.A2(n_83),
.B(n_231),
.Y(n_303)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_40),
.B(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_43),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_43),
.A2(n_46),
.B1(n_258),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_43),
.A2(n_46),
.B1(n_89),
.B2(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_45),
.Y(n_169)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_47),
.B(n_48),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_49),
.A2(n_161),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_64),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_57),
.A2(n_59),
.B1(n_181),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_57),
.A2(n_216),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_59),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_59),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_59),
.A2(n_182),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_64),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_65),
.A2(n_73),
.B1(n_116),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_65),
.A2(n_159),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_65),
.A2(n_73),
.B1(n_213),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_65),
.A2(n_73),
.B1(n_243),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_65),
.A2(n_73),
.B1(n_252),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_66),
.A2(n_69),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_71),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_70),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_71),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_73),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_73),
.A2(n_118),
.B(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_74),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.C(n_85),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_82),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_82),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_85),
.B(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_319),
.A3(n_329),
.B1(n_334),
.B2(n_335),
.C(n_337),
.Y(n_92)
);

AOI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_269),
.A3(n_307),
.B1(n_313),
.B2(n_318),
.C(n_338),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_224),
.C(n_265),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_196),
.B(n_223),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_175),
.B(n_195),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_153),
.B(n_174),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_128),
.B(n_152),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_100),
.B(n_110),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_138),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B(n_125),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_123),
.A2(n_124),
.B1(n_172),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_123),
.A2(n_136),
.B1(n_186),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_123),
.A2(n_206),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_123),
.A2(n_136),
.B1(n_241),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_123),
.A2(n_124),
.B(n_250),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_132),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_142),
.Y(n_149)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_139),
.B(n_151),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_137),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_146),
.B(n_150),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_143),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_166),
.B2(n_173),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_165),
.C(n_173),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_177),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_191),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_192),
.C(n_193),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_190),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_187),
.C(n_188),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_198),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_210),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_209),
.C(n_210),
.Y(n_266)
);

AOI22x1_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_205),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_225),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_245),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_226),
.B(n_245),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.C(n_244),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_263),
.B2(n_264),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_253),
.C(n_264),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_251),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_259),
.C(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_267),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_287),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_270),
.B(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.C(n_286),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_271),
.A2(n_272),
.B1(n_280),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_282),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_299),
.B(n_303),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_283),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_305),
.B2(n_306),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_298),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_298),
.C(n_306),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_295),
.B(n_296),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_295),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_296),
.A2(n_321),
.B1(n_325),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_301),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.C(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);


endmodule