module fake_jpeg_29559_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVxp67_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NOR3xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_3),
.C(n_4),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_17),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_19),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_1),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_12),
.B1(n_6),
.B2(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_20),
.B1(n_16),
.B2(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_28),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_17),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_23),
.Y(n_29)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_14),
.B1(n_15),
.B2(n_21),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_21),
.C(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

AOI31xp33_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_19),
.A3(n_9),
.B(n_28),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_30),
.B(n_15),
.Y(n_36)
);


endmodule