module real_aes_17725_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_1840;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_1749;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1842;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_0), .A2(n_281), .B1(n_847), .B2(n_848), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_0), .A2(n_176), .B1(n_773), .B2(n_891), .Y(n_897) );
XNOR2xp5_ASAP7_75t_L g903 ( .A(n_1), .B(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g979 ( .A(n_2), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1853 ( .A1(n_3), .A2(n_57), .B1(n_576), .B2(n_750), .Y(n_1853) );
INVxp67_ASAP7_75t_SL g1869 ( .A(n_3), .Y(n_1869) );
INVx1_ASAP7_75t_L g1323 ( .A(n_4), .Y(n_1323) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_5), .A2(n_269), .B1(n_675), .B2(n_679), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_5), .A2(n_356), .B1(n_714), .B2(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g436 ( .A(n_6), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_6), .B(n_397), .Y(n_502) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_6), .B(n_401), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_6), .B(n_263), .Y(n_1755) );
INVx1_ASAP7_75t_L g868 ( .A(n_7), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_7), .A2(n_199), .B1(n_732), .B2(n_879), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_8), .Y(n_1179) );
INVx1_ASAP7_75t_L g504 ( .A(n_9), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_10), .A2(n_267), .B1(n_679), .B2(n_1287), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_10), .A2(n_206), .B1(n_1075), .B2(n_1083), .Y(n_1303) );
OAI22xp33_ASAP7_75t_SL g1202 ( .A1(n_11), .A2(n_363), .B1(n_743), .B2(n_1105), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1213 ( .A1(n_11), .A2(n_190), .B1(n_481), .B2(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1277 ( .A(n_12), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_12), .A2(n_267), .B1(n_1083), .B2(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g988 ( .A(n_13), .Y(n_988) );
INVx1_ASAP7_75t_L g874 ( .A(n_14), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_15), .Y(n_613) );
INVx1_ASAP7_75t_L g1837 ( .A(n_16), .Y(n_1837) );
INVx1_ASAP7_75t_L g1362 ( .A(n_17), .Y(n_1362) );
OAI221xp5_ASAP7_75t_L g1369 ( .A1(n_17), .A2(n_317), .B1(n_733), .B2(n_790), .C(n_1370), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_18), .A2(n_115), .B1(n_847), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g889 ( .A(n_18), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g1224 ( .A(n_19), .Y(n_1224) );
XOR2x2_ASAP7_75t_L g722 ( .A(n_20), .B(n_723), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_21), .A2(n_335), .B1(n_425), .B2(n_427), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_21), .A2(n_335), .B1(n_443), .B2(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g447 ( .A(n_22), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g1555 ( .A1(n_23), .A2(n_24), .B1(n_1526), .B2(n_1534), .Y(n_1555) );
OAI22xp33_ASAP7_75t_SL g1413 ( .A1(n_25), .A2(n_280), .B1(n_481), .B2(n_1214), .Y(n_1413) );
OAI22xp33_ASAP7_75t_L g1421 ( .A1(n_25), .A2(n_280), .B1(n_743), .B2(n_1138), .Y(n_1421) );
INVx1_ASAP7_75t_L g1120 ( .A(n_26), .Y(n_1120) );
INVx1_ASAP7_75t_L g1742 ( .A(n_27), .Y(n_1742) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_28), .A2(n_188), .B1(n_1078), .B2(n_1080), .Y(n_1077) );
AOI22xp33_ASAP7_75t_SL g1098 ( .A1(n_28), .A2(n_139), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_29), .A2(n_296), .B1(n_1376), .B2(n_1378), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_29), .A2(n_162), .B1(n_771), .B2(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1115 ( .A(n_30), .Y(n_1115) );
OAI211xp5_ASAP7_75t_L g1139 ( .A1(n_31), .A2(n_953), .B(n_1140), .C(n_1144), .Y(n_1139) );
INVx1_ASAP7_75t_L g1153 ( .A(n_31), .Y(n_1153) );
INVx1_ASAP7_75t_L g1429 ( .A(n_32), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g1334 ( .A1(n_33), .A2(n_84), .B1(n_444), .B2(n_1214), .C(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1346 ( .A(n_33), .Y(n_1346) );
HB1xp67_ASAP7_75t_L g1511 ( .A(n_34), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_34), .B(n_1509), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1594 ( .A1(n_35), .A2(n_202), .B1(n_1534), .B2(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g915 ( .A(n_36), .Y(n_915) );
OAI22xp33_ASAP7_75t_SL g424 ( .A1(n_37), .A2(n_177), .B1(n_425), .B2(n_427), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_37), .A2(n_177), .B1(n_443), .B2(n_452), .Y(n_442) );
OAI222xp33_ASAP7_75t_L g1064 ( .A1(n_38), .A2(n_211), .B1(n_362), .B2(n_664), .C1(n_1065), .C2(n_1066), .Y(n_1064) );
OAI222xp33_ASAP7_75t_L g1107 ( .A1(n_38), .A2(n_211), .B1(n_362), .B2(n_518), .C1(n_576), .C2(n_750), .Y(n_1107) );
OAI211xp5_ASAP7_75t_SL g1737 ( .A1(n_39), .A2(n_1738), .B(n_1741), .C(n_1747), .Y(n_1737) );
OAI22xp5_ASAP7_75t_L g1805 ( .A1(n_39), .A2(n_290), .B1(n_1806), .B2(n_1810), .Y(n_1805) );
CKINVDCx5p33_ASAP7_75t_R g1477 ( .A(n_40), .Y(n_1477) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_41), .A2(n_276), .B1(n_679), .B2(n_761), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_41), .A2(n_161), .B1(n_770), .B2(n_771), .Y(n_775) );
INVx1_ASAP7_75t_L g1022 ( .A(n_42), .Y(n_1022) );
INVxp67_ASAP7_75t_SL g1852 ( .A(n_43), .Y(n_1852) );
OAI22xp5_ASAP7_75t_L g1870 ( .A1(n_43), .A2(n_57), .B1(n_664), .B2(n_1065), .Y(n_1870) );
OAI221xp5_ASAP7_75t_L g1756 ( .A1(n_44), .A2(n_120), .B1(n_1757), .B2(n_1761), .C(n_1765), .Y(n_1756) );
OAI22xp33_ASAP7_75t_L g1789 ( .A1(n_44), .A2(n_120), .B1(n_1790), .B2(n_1792), .Y(n_1789) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_45), .A2(n_309), .B1(n_657), .B2(n_658), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_45), .A2(n_309), .B1(n_444), .B2(n_454), .Y(n_662) );
XNOR2x1_ASAP7_75t_L g1391 ( .A(n_46), .B(n_1392), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1608 ( .A1(n_46), .A2(n_220), .B1(n_1526), .B2(n_1531), .Y(n_1608) );
AOI22xp33_ASAP7_75t_SL g1768 ( .A1(n_47), .A2(n_272), .B1(n_1100), .B2(n_1381), .Y(n_1768) );
AOI22xp33_ASAP7_75t_L g1784 ( .A1(n_47), .A2(n_368), .B1(n_714), .B2(n_1083), .Y(n_1784) );
AOI22xp5_ASAP7_75t_L g1541 ( .A1(n_48), .A2(n_354), .B1(n_1534), .B2(n_1542), .Y(n_1541) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_49), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_50), .Y(n_1275) );
INVx1_ASAP7_75t_L g919 ( .A(n_51), .Y(n_919) );
INVx1_ASAP7_75t_L g828 ( .A(n_52), .Y(n_828) );
INVx1_ASAP7_75t_L g1326 ( .A(n_53), .Y(n_1326) );
AOI22xp5_ASAP7_75t_L g1609 ( .A1(n_54), .A2(n_331), .B1(n_1534), .B2(n_1595), .Y(n_1609) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_55), .A2(n_273), .B1(n_682), .B2(n_685), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_55), .A2(n_89), .B1(n_710), .B2(n_712), .Y(n_709) );
XNOR2xp5_ASAP7_75t_L g949 ( .A(n_56), .B(n_950), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_56), .A2(n_129), .B1(n_1526), .B2(n_1531), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_58), .B(n_473), .Y(n_1336) );
INVxp67_ASAP7_75t_SL g1343 ( .A(n_58), .Y(n_1343) );
OAI211xp5_ASAP7_75t_L g1196 ( .A1(n_59), .A2(n_1197), .B(n_1198), .C(n_1199), .Y(n_1196) );
INVx1_ASAP7_75t_L g1212 ( .A(n_59), .Y(n_1212) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_60), .A2(n_244), .B1(n_444), .B2(n_582), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_60), .A2(n_244), .B1(n_426), .B2(n_802), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g1169 ( .A(n_61), .Y(n_1169) );
INVx1_ASAP7_75t_L g1855 ( .A(n_62), .Y(n_1855) );
INVx1_ASAP7_75t_L g825 ( .A(n_63), .Y(n_825) );
OAI222xp33_ASAP7_75t_L g1264 ( .A1(n_64), .A2(n_193), .B1(n_654), .B2(n_744), .C1(n_1265), .C2(n_1266), .Y(n_1264) );
OAI222xp33_ASAP7_75t_L g1293 ( .A1(n_64), .A2(n_193), .B1(n_232), .B2(n_732), .C1(n_1294), .C2(n_1295), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_65), .A2(n_126), .B1(n_657), .B2(n_658), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_65), .A2(n_126), .B1(n_444), .B2(n_454), .Y(n_1371) );
OAI22xp33_ASAP7_75t_L g1038 ( .A1(n_66), .A2(n_321), .B1(n_389), .B2(n_398), .Y(n_1038) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_66), .A2(n_321), .B1(n_591), .B2(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1143 ( .A(n_67), .Y(n_1143) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_67), .A2(n_631), .B(n_968), .C(n_1151), .Y(n_1150) );
OAI22xp33_ASAP7_75t_L g1339 ( .A1(n_68), .A2(n_195), .B1(n_481), .B2(n_1063), .Y(n_1339) );
INVxp67_ASAP7_75t_SL g1345 ( .A(n_68), .Y(n_1345) );
CKINVDCx5p33_ASAP7_75t_R g1234 ( .A(n_69), .Y(n_1234) );
INVx1_ASAP7_75t_L g1856 ( .A(n_70), .Y(n_1856) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_71), .Y(n_1442) );
INVx1_ASAP7_75t_L g1406 ( .A(n_72), .Y(n_1406) );
INVx1_ASAP7_75t_L g1848 ( .A(n_73), .Y(n_1848) );
INVx1_ASAP7_75t_L g844 ( .A(n_74), .Y(n_844) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_75), .A2(n_645), .B(n_646), .C(n_650), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_75), .A2(n_213), .B1(n_587), .B2(n_664), .C(n_665), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g1767 ( .A1(n_76), .A2(n_766), .B(n_1284), .Y(n_1767) );
INVx1_ASAP7_75t_L g1780 ( .A(n_76), .Y(n_1780) );
XNOR2xp5_ASAP7_75t_L g1351 ( .A(n_77), .B(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g958 ( .A(n_78), .Y(n_958) );
OAI211xp5_ASAP7_75t_L g967 ( .A1(n_78), .A2(n_631), .B(n_968), .C(n_969), .Y(n_967) );
INVx1_ASAP7_75t_L g1325 ( .A(n_79), .Y(n_1325) );
INVx1_ASAP7_75t_L g537 ( .A(n_80), .Y(n_537) );
INVx1_ASAP7_75t_L g913 ( .A(n_81), .Y(n_913) );
OAI22xp33_ASAP7_75t_L g1419 ( .A1(n_82), .A2(n_113), .B1(n_444), .B2(n_454), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_82), .A2(n_113), .B1(n_657), .B2(n_658), .Y(n_1425) );
XNOR2xp5_ASAP7_75t_L g1466 ( .A(n_83), .B(n_1467), .Y(n_1466) );
AOI22xp5_ASAP7_75t_L g1549 ( .A1(n_83), .A2(n_367), .B1(n_1526), .B2(n_1531), .Y(n_1549) );
OAI22xp33_ASAP7_75t_L g1348 ( .A1(n_84), .A2(n_195), .B1(n_743), .B2(n_1138), .Y(n_1348) );
INVx1_ASAP7_75t_L g1122 ( .A(n_85), .Y(n_1122) );
INVx1_ASAP7_75t_L g1457 ( .A(n_86), .Y(n_1457) );
OAI211xp5_ASAP7_75t_L g1462 ( .A1(n_86), .A2(n_466), .B(n_546), .C(n_1463), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1244 ( .A1(n_87), .A2(n_284), .B1(n_658), .B2(n_743), .Y(n_1244) );
OAI22xp5_ASAP7_75t_SL g1252 ( .A1(n_87), .A2(n_135), .B1(n_454), .B2(n_481), .Y(n_1252) );
INVx1_ASAP7_75t_L g1338 ( .A(n_88), .Y(n_1338) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_89), .A2(n_369), .B1(n_679), .B2(n_690), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g1247 ( .A(n_90), .Y(n_1247) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_91), .Y(n_1222) );
OAI22xp33_ASAP7_75t_L g1137 ( .A1(n_92), .A2(n_168), .B1(n_389), .B2(n_1138), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_92), .A2(n_168), .B1(n_975), .B2(n_1149), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_93), .Y(n_1167) );
OAI211xp5_ASAP7_75t_L g787 ( .A1(n_94), .A2(n_466), .B(n_788), .C(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g800 ( .A(n_94), .Y(n_800) );
AOI22xp5_ASAP7_75t_SL g1550 ( .A1(n_95), .A2(n_229), .B1(n_1534), .B2(n_1542), .Y(n_1550) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_96), .A2(n_256), .B1(n_1096), .B2(n_1376), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_96), .A2(n_173), .B1(n_714), .B2(n_1076), .Y(n_1386) );
XOR2xp5_ASAP7_75t_L g1161 ( .A(n_97), .B(n_1162), .Y(n_1161) );
XNOR2x2_ASAP7_75t_SL g783 ( .A(n_98), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g916 ( .A(n_99), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g1480 ( .A(n_100), .Y(n_1480) );
INVx1_ASAP7_75t_L g1838 ( .A(n_101), .Y(n_1838) );
AOI22xp33_ASAP7_75t_L g1866 ( .A1(n_101), .A2(n_307), .B1(n_675), .B2(n_1862), .Y(n_1866) );
CKINVDCx5p33_ASAP7_75t_R g1231 ( .A(n_102), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_103), .A2(n_147), .B1(n_398), .B2(n_743), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_103), .A2(n_133), .B1(n_443), .B2(n_481), .Y(n_938) );
INVx1_ASAP7_75t_L g909 ( .A(n_104), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_105), .A2(n_233), .B1(n_732), .B2(n_733), .Y(n_731) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_105), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_106), .A2(n_304), .B1(n_679), .B2(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_106), .A2(n_271), .B1(n_773), .B2(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g921 ( .A(n_107), .Y(n_921) );
INVx1_ASAP7_75t_L g1026 ( .A(n_108), .Y(n_1026) );
OAI211xp5_ASAP7_75t_L g1454 ( .A1(n_109), .A2(n_604), .B(n_1198), .C(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1464 ( .A(n_109), .Y(n_1464) );
INVx1_ASAP7_75t_L g1509 ( .A(n_110), .Y(n_1509) );
INVx1_ASAP7_75t_L g1844 ( .A(n_111), .Y(n_1844) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_112), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_112), .A2(n_233), .B1(n_576), .B2(n_750), .Y(n_749) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_114), .A2(n_312), .B1(n_398), .B2(n_426), .Y(n_1459) );
OAI22xp33_ASAP7_75t_L g1465 ( .A1(n_114), .A2(n_165), .B1(n_444), .B2(n_454), .Y(n_1465) );
INVxp67_ASAP7_75t_SL g896 ( .A(n_115), .Y(n_896) );
XNOR2xp5_ASAP7_75t_L g1826 ( .A(n_116), .B(n_1827), .Y(n_1826) );
XOR2xp5_ASAP7_75t_L g1257 ( .A(n_117), .B(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g982 ( .A(n_118), .Y(n_982) );
INVx1_ASAP7_75t_L g1399 ( .A(n_119), .Y(n_1399) );
INVx1_ASAP7_75t_L g1396 ( .A(n_121), .Y(n_1396) );
AOI22xp5_ASAP7_75t_L g1546 ( .A1(n_122), .A2(n_342), .B1(n_1531), .B2(n_1542), .Y(n_1546) );
INVx1_ASAP7_75t_L g419 ( .A(n_123), .Y(n_419) );
INVx1_ASAP7_75t_L g869 ( .A(n_124), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_125), .Y(n_931) );
INVx1_ASAP7_75t_L g1015 ( .A(n_127), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1752 ( .A1(n_128), .A2(n_246), .B1(n_1099), .B2(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1783 ( .A(n_128), .Y(n_1783) );
INVx1_ASAP7_75t_L g1835 ( .A(n_130), .Y(n_1835) );
INVx1_ASAP7_75t_L g511 ( .A(n_131), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_132), .A2(n_266), .B1(n_884), .B2(n_1063), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_132), .A2(n_266), .B1(n_934), .B2(n_1105), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_133), .A2(n_227), .B1(n_802), .B2(n_934), .Y(n_933) );
OAI22xp33_ASAP7_75t_SL g1249 ( .A1(n_134), .A2(n_135), .B1(n_657), .B2(n_1138), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_134), .A2(n_137), .B1(n_1210), .B2(n_1211), .Y(n_1255) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_136), .Y(n_608) );
INVx1_ASAP7_75t_L g1248 ( .A(n_137), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_138), .A2(n_361), .B1(n_481), .B2(n_795), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g803 ( .A1(n_138), .A2(n_361), .B1(n_398), .B2(n_743), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_139), .A2(n_305), .B1(n_712), .B2(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g827 ( .A(n_140), .Y(n_827) );
INVx1_ASAP7_75t_L g1355 ( .A(n_141), .Y(n_1355) );
INVx1_ASAP7_75t_L g1418 ( .A(n_142), .Y(n_1418) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_142), .A2(n_853), .B(n_1198), .C(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g845 ( .A(n_143), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g1417 ( .A(n_144), .Y(n_1417) );
INVx1_ASAP7_75t_L g1117 ( .A(n_145), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_146), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_147), .A2(n_227), .B1(n_591), .B2(n_944), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g1478 ( .A(n_148), .Y(n_1478) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_149), .A2(n_196), .B1(n_398), .B2(n_657), .Y(n_1493) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_149), .A2(n_187), .B1(n_444), .B2(n_454), .Y(n_1499) );
CKINVDCx5p33_ASAP7_75t_R g1227 ( .A(n_150), .Y(n_1227) );
CKINVDCx5p33_ASAP7_75t_R g1471 ( .A(n_151), .Y(n_1471) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_152), .A2(n_405), .B(n_410), .C(n_415), .Y(n_404) );
INVx1_ASAP7_75t_L g475 ( .A(n_152), .Y(n_475) );
INVx1_ASAP7_75t_L g423 ( .A(n_153), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g458 ( .A1(n_153), .A2(n_459), .B(n_466), .C(n_470), .Y(n_458) );
INVx1_ASAP7_75t_L g822 ( .A(n_154), .Y(n_822) );
INVx1_ASAP7_75t_L g1124 ( .A(n_155), .Y(n_1124) );
INVx1_ASAP7_75t_L g506 ( .A(n_156), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g1171 ( .A(n_157), .Y(n_1171) );
OAI211xp5_ASAP7_75t_L g1033 ( .A1(n_158), .A2(n_407), .B(n_410), .C(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1046 ( .A(n_158), .Y(n_1046) );
INVx1_ASAP7_75t_L g911 ( .A(n_159), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_160), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_161), .A2(n_348), .B1(n_756), .B2(n_759), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g1380 ( .A1(n_162), .A2(n_216), .B1(n_858), .B2(n_1381), .Y(n_1380) );
AOI221xp5_ASAP7_75t_L g1748 ( .A1(n_163), .A2(n_368), .B1(n_1749), .B2(n_1750), .C(n_1751), .Y(n_1748) );
AOI22xp33_ASAP7_75t_L g1788 ( .A1(n_163), .A2(n_272), .B1(n_714), .B2(n_877), .Y(n_1788) );
INVx1_ASAP7_75t_L g1035 ( .A(n_164), .Y(n_1035) );
OAI22xp33_ASAP7_75t_L g1458 ( .A1(n_165), .A2(n_287), .B1(n_743), .B2(n_864), .Y(n_1458) );
INVx1_ASAP7_75t_L g1491 ( .A(n_166), .Y(n_1491) );
OAI211xp5_ASAP7_75t_L g1496 ( .A1(n_166), .A2(n_466), .B(n_546), .C(n_1497), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g1434 ( .A(n_167), .Y(n_1434) );
INVx1_ASAP7_75t_L g1322 ( .A(n_169), .Y(n_1322) );
INVx1_ASAP7_75t_L g957 ( .A(n_170), .Y(n_957) );
INVx1_ASAP7_75t_L g1357 ( .A(n_171), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_172), .A2(n_303), .B1(n_425), .B2(n_427), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_172), .A2(n_303), .B1(n_443), .B2(n_452), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_173), .A2(n_277), .B1(n_1099), .B2(n_1100), .Y(n_1374) );
OAI211xp5_ASAP7_75t_L g1488 ( .A1(n_174), .A2(n_604), .B(n_1198), .C(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1498 ( .A(n_174), .Y(n_1498) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_175), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_175), .A2(n_281), .B1(n_891), .B2(n_892), .Y(n_890) );
INVxp67_ASAP7_75t_SL g854 ( .A(n_176), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_178), .Y(n_1176) );
XNOR2xp5_ASAP7_75t_L g840 ( .A(n_179), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1591 ( .A(n_179), .Y(n_1591) );
CKINVDCx5p33_ASAP7_75t_R g1361 ( .A(n_180), .Y(n_1361) );
AOI22xp5_ASAP7_75t_SL g1561 ( .A1(n_181), .A2(n_191), .B1(n_1534), .B2(n_1542), .Y(n_1561) );
INVx1_ASAP7_75t_L g536 ( .A(n_182), .Y(n_536) );
INVx1_ASAP7_75t_L g1025 ( .A(n_183), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_184), .A2(n_264), .B1(n_934), .B2(n_961), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_184), .A2(n_264), .B1(n_965), .B2(n_966), .Y(n_964) );
OAI22xp33_ASAP7_75t_L g1492 ( .A1(n_185), .A2(n_187), .B1(n_743), .B2(n_864), .Y(n_1492) );
OAI22xp33_ASAP7_75t_L g1495 ( .A1(n_185), .A2(n_196), .B1(n_481), .B2(n_1214), .Y(n_1495) );
INVx1_ASAP7_75t_L g992 ( .A(n_186), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_188), .A2(n_305), .B1(n_1092), .B2(n_1096), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g1414 ( .A1(n_189), .A2(n_466), .B(n_1415), .C(n_1416), .Y(n_1414) );
INVx1_ASAP7_75t_L g1424 ( .A(n_189), .Y(n_1424) );
OAI22xp33_ASAP7_75t_SL g1203 ( .A1(n_190), .A2(n_324), .B1(n_398), .B2(n_426), .Y(n_1203) );
INVx1_ASAP7_75t_L g1011 ( .A(n_192), .Y(n_1011) );
INVx2_ASAP7_75t_L g1529 ( .A(n_194), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_194), .B(n_1530), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_194), .B(n_318), .Y(n_1537) );
AOI22xp5_ASAP7_75t_SL g1554 ( .A1(n_197), .A2(n_274), .B1(n_1531), .B2(n_1536), .Y(n_1554) );
XNOR2xp5_ASAP7_75t_L g1734 ( .A(n_197), .B(n_1735), .Y(n_1734) );
AOI22xp33_ASAP7_75t_L g1821 ( .A1(n_197), .A2(n_1822), .B1(n_1825), .B2(n_1873), .Y(n_1821) );
CKINVDCx5p33_ASAP7_75t_R g1475 ( .A(n_198), .Y(n_1475) );
INVx1_ASAP7_75t_L g871 ( .A(n_199), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_200), .Y(n_1230) );
INVx1_ASAP7_75t_L g987 ( .A(n_201), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g1533 ( .A1(n_203), .A2(n_339), .B1(n_1534), .B2(n_1536), .Y(n_1533) );
INVx1_ASAP7_75t_L g642 ( .A(n_204), .Y(n_642) );
INVx1_ASAP7_75t_L g932 ( .A(n_205), .Y(n_932) );
OAI211xp5_ASAP7_75t_L g939 ( .A1(n_205), .A2(n_466), .B(n_940), .C(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g1280 ( .A(n_206), .Y(n_1280) );
XOR2xp5_ASAP7_75t_L g1310 ( .A(n_207), .B(n_1311), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1540 ( .A1(n_207), .A2(n_278), .B1(n_1526), .B2(n_1531), .Y(n_1540) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_208), .A2(n_350), .B1(n_1072), .B2(n_1082), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_208), .A2(n_255), .B1(n_1092), .B2(n_1096), .Y(n_1097) );
XNOR2x2_ASAP7_75t_L g1109 ( .A(n_209), .B(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1316 ( .A(n_210), .Y(n_1316) );
CKINVDCx5p33_ASAP7_75t_R g1440 ( .A(n_212), .Y(n_1440) );
INVx1_ASAP7_75t_L g655 ( .A(n_213), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_214), .A2(n_271), .B1(n_759), .B2(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_214), .A2(n_304), .B1(n_714), .B2(n_773), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g1547 ( .A1(n_215), .A2(n_295), .B1(n_1526), .B2(n_1534), .Y(n_1547) );
AOI22xp33_ASAP7_75t_SL g1388 ( .A1(n_216), .A2(n_296), .B1(n_771), .B2(n_815), .Y(n_1388) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_217), .Y(n_574) );
OAI211xp5_ASAP7_75t_L g1260 ( .A1(n_218), .A2(n_1261), .B(n_1262), .C(n_1270), .Y(n_1260) );
INVx1_ASAP7_75t_L g1298 ( .A(n_218), .Y(n_1298) );
INVx1_ASAP7_75t_L g1017 ( .A(n_219), .Y(n_1017) );
INVx1_ASAP7_75t_L g1319 ( .A(n_221), .Y(n_1319) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_222), .A2(n_306), .B1(n_389), .B2(n_398), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_222), .A2(n_306), .B1(n_479), .B2(n_482), .Y(n_478) );
INVx2_ASAP7_75t_L g491 ( .A(n_223), .Y(n_491) );
INVx1_ASAP7_75t_L g565 ( .A(n_223), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g1801 ( .A(n_223), .B(n_447), .Y(n_1801) );
CKINVDCx5p33_ASAP7_75t_R g1435 ( .A(n_224), .Y(n_1435) );
INVx1_ASAP7_75t_L g1804 ( .A(n_225), .Y(n_1804) );
INVx1_ASAP7_75t_L g809 ( .A(n_226), .Y(n_809) );
INVx1_ASAP7_75t_L g1403 ( .A(n_228), .Y(n_1403) );
XOR2xp5_ASAP7_75t_L g1055 ( .A(n_230), .B(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1269 ( .A(n_231), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_231), .A2(n_262), .B1(n_444), .B2(n_454), .Y(n_1296) );
INVx1_ASAP7_75t_L g1263 ( .A(n_232), .Y(n_1263) );
BUFx3_ASAP7_75t_L g449 ( .A(n_234), .Y(n_449) );
INVx1_ASAP7_75t_L g1397 ( .A(n_235), .Y(n_1397) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_236), .Y(n_1445) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_237), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_238), .Y(n_1481) );
XOR2xp5_ASAP7_75t_L g1006 ( .A(n_239), .B(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_240), .A2(n_255), .B1(n_1072), .B2(n_1076), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_240), .A2(n_350), .B1(n_761), .B2(n_1090), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g1525 ( .A1(n_241), .A2(n_292), .B1(n_1526), .B2(n_1531), .Y(n_1525) );
INVx1_ASAP7_75t_L g1840 ( .A(n_242), .Y(n_1840) );
INVx1_ASAP7_75t_L g577 ( .A(n_243), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g584 ( .A1(n_243), .A2(n_466), .B(n_585), .C(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g1274 ( .A(n_245), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_245), .B(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1787 ( .A(n_246), .Y(n_1787) );
INVx1_ASAP7_75t_L g727 ( .A(n_247), .Y(n_727) );
INVx1_ASAP7_75t_L g1012 ( .A(n_248), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1474 ( .A(n_249), .Y(n_1474) );
CKINVDCx5p33_ASAP7_75t_R g1437 ( .A(n_250), .Y(n_1437) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_251), .A2(n_338), .B1(n_389), .B2(n_398), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_251), .A2(n_338), .B1(n_591), .B2(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g517 ( .A(n_252), .Y(n_517) );
INVx1_ASAP7_75t_L g652 ( .A(n_253), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_254), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g1389 ( .A1(n_256), .A2(n_277), .B1(n_714), .B2(n_773), .C(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1843 ( .A(n_257), .Y(n_1843) );
AOI22xp33_ASAP7_75t_L g1860 ( .A1(n_257), .A2(n_319), .B1(n_1861), .B2(n_1862), .Y(n_1860) );
INVx1_ASAP7_75t_L g1402 ( .A(n_258), .Y(n_1402) );
INVx1_ASAP7_75t_L g1745 ( .A(n_259), .Y(n_1745) );
INVx1_ASAP7_75t_L g985 ( .A(n_260), .Y(n_985) );
XOR2xp5_ASAP7_75t_L g1217 ( .A(n_261), .B(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1271 ( .A(n_262), .Y(n_1271) );
BUFx3_ASAP7_75t_L g397 ( .A(n_263), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_263), .Y(n_401) );
INVx1_ASAP7_75t_L g1141 ( .A(n_265), .Y(n_1141) );
INVx1_ASAP7_75t_L g1315 ( .A(n_268), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_269), .A2(n_316), .B1(n_696), .B2(n_700), .Y(n_695) );
INVx1_ASAP7_75t_L g792 ( .A(n_270), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_273), .A2(n_369), .B1(n_703), .B2(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g1127 ( .A(n_275), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_276), .A2(n_348), .B1(n_770), .B2(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g1060 ( .A(n_279), .Y(n_1060) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_282), .Y(n_1174) );
INVx1_ASAP7_75t_L g873 ( .A(n_283), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_284), .B(n_444), .Y(n_1251) );
INVx1_ASAP7_75t_L g808 ( .A(n_285), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g1233 ( .A(n_286), .Y(n_1233) );
OAI22xp33_ASAP7_75t_L g1461 ( .A1(n_287), .A2(n_312), .B1(n_481), .B2(n_1214), .Y(n_1461) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_288), .Y(n_1177) );
INVx1_ASAP7_75t_L g793 ( .A(n_289), .Y(n_793) );
OAI211xp5_ASAP7_75t_L g797 ( .A1(n_289), .A2(n_571), .B(n_798), .C(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g726 ( .A(n_291), .Y(n_726) );
XOR2x2_ASAP7_75t_L g385 ( .A(n_293), .B(n_386), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g1472 ( .A(n_294), .Y(n_1472) );
INVx1_ASAP7_75t_L g451 ( .A(n_297), .Y(n_451) );
INVx1_ASAP7_75t_L g457 ( .A(n_297), .Y(n_457) );
INVx1_ASAP7_75t_L g1126 ( .A(n_298), .Y(n_1126) );
INVx1_ASAP7_75t_L g1119 ( .A(n_299), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_300), .A2(n_358), .B1(n_934), .B2(n_1146), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_300), .A2(n_358), .B1(n_443), .B2(n_582), .Y(n_1154) );
INVx1_ASAP7_75t_L g817 ( .A(n_301), .Y(n_817) );
INVx1_ASAP7_75t_L g862 ( .A(n_302), .Y(n_862) );
INVx1_ASAP7_75t_L g1841 ( .A(n_307), .Y(n_1841) );
INVx1_ASAP7_75t_L g1200 ( .A(n_308), .Y(n_1200) );
OAI211xp5_ASAP7_75t_SL g1206 ( .A1(n_308), .A2(n_968), .B(n_1065), .C(n_1207), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_310), .A2(n_311), .B1(n_389), .B2(n_398), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_310), .A2(n_311), .B1(n_479), .B2(n_591), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g1766 ( .A(n_313), .Y(n_1766) );
INVx1_ASAP7_75t_L g813 ( .A(n_314), .Y(n_813) );
INVx1_ASAP7_75t_L g1318 ( .A(n_315), .Y(n_1318) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_316), .A2(n_356), .B1(n_682), .B2(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g1364 ( .A(n_317), .Y(n_1364) );
INVx1_ASAP7_75t_L g1530 ( .A(n_318), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_318), .B(n_1529), .Y(n_1535) );
INVx1_ASAP7_75t_L g1832 ( .A(n_319), .Y(n_1832) );
INVx1_ASAP7_75t_L g736 ( .A(n_320), .Y(n_736) );
INVx1_ASAP7_75t_L g1405 ( .A(n_322), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1438 ( .A(n_323), .Y(n_1438) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_324), .A2(n_363), .B1(n_444), .B2(n_454), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_325), .Y(n_595) );
INVx1_ASAP7_75t_L g1059 ( .A(n_326), .Y(n_1059) );
INVx1_ASAP7_75t_L g1847 ( .A(n_327), .Y(n_1847) );
CKINVDCx5p33_ASAP7_75t_R g1490 ( .A(n_328), .Y(n_1490) );
INVx1_ASAP7_75t_L g1593 ( .A(n_329), .Y(n_1593) );
CKINVDCx5p33_ASAP7_75t_R g1282 ( .A(n_330), .Y(n_1282) );
OAI211xp5_ASAP7_75t_SL g1245 ( .A1(n_332), .A2(n_1197), .B(n_1198), .C(n_1246), .Y(n_1245) );
OAI211xp5_ASAP7_75t_SL g1253 ( .A1(n_332), .A2(n_879), .B(n_968), .C(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1400 ( .A(n_333), .Y(n_1400) );
INVx1_ASAP7_75t_L g1337 ( .A(n_334), .Y(n_1337) );
OAI211xp5_ASAP7_75t_L g570 ( .A1(n_336), .A2(n_407), .B(n_571), .C(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g589 ( .A(n_336), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g928 ( .A1(n_337), .A2(n_571), .B(n_929), .C(n_930), .Y(n_928) );
INVx1_ASAP7_75t_L g942 ( .A(n_337), .Y(n_942) );
INVx1_ASAP7_75t_L g865 ( .A(n_340), .Y(n_865) );
INVx1_ASAP7_75t_L g1036 ( .A(n_341), .Y(n_1036) );
OAI211xp5_ASAP7_75t_L g1044 ( .A1(n_341), .A2(n_460), .B(n_466), .C(n_1045), .Y(n_1044) );
OAI211xp5_ASAP7_75t_SL g952 ( .A1(n_343), .A2(n_571), .B(n_953), .C(n_955), .Y(n_952) );
INVx1_ASAP7_75t_L g972 ( .A(n_343), .Y(n_972) );
INVx1_ASAP7_75t_L g980 ( .A(n_344), .Y(n_980) );
INVx1_ASAP7_75t_L g640 ( .A(n_345), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_346), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_347), .Y(n_597) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
INVx1_ASAP7_75t_L g523 ( .A(n_351), .Y(n_523) );
INVx1_ASAP7_75t_L g1021 ( .A(n_352), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_353), .Y(n_601) );
OA22x2_ASAP7_75t_L g636 ( .A1(n_355), .A2(n_637), .B1(n_720), .B2(n_721), .Y(n_636) );
INVxp67_ASAP7_75t_SL g721 ( .A(n_355), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_357), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1201 ( .A(n_359), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_360), .Y(n_1226) );
XOR2x2_ASAP7_75t_L g567 ( .A(n_364), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g440 ( .A(n_365), .Y(n_440) );
INVx2_ASAP7_75t_L g501 ( .A(n_365), .Y(n_501) );
INVx1_ASAP7_75t_L g564 ( .A(n_365), .Y(n_564) );
INVx1_ASAP7_75t_L g908 ( .A(n_366), .Y(n_908) );
INVx1_ASAP7_75t_L g738 ( .A(n_370), .Y(n_738) );
INVx1_ASAP7_75t_L g526 ( .A(n_371), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g1283 ( .A1(n_372), .A2(n_766), .B(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1301 ( .A(n_372), .Y(n_1301) );
CKINVDCx5p33_ASAP7_75t_R g1446 ( .A(n_373), .Y(n_1446) );
CKINVDCx5p33_ASAP7_75t_R g1267 ( .A(n_374), .Y(n_1267) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_1503), .B(n_1515), .Y(n_375) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_1049), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B1(n_946), .B2(n_1048), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
XNOR2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_633), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_567), .B2(n_632), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_441), .C(n_495), .Y(n_386) );
OAI31xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_404), .A3(n_424), .B(n_433), .Y(n_387) );
INVx3_ASAP7_75t_L g641 ( .A(n_389), .Y(n_641) );
OR2x6_ASAP7_75t_L g389 ( .A(n_390), .B(n_395), .Y(n_389) );
OR2x6_ASAP7_75t_L g426 ( .A(n_390), .B(n_400), .Y(n_426) );
BUFx4f_ASAP7_75t_L g505 ( .A(n_390), .Y(n_505) );
OR2x2_ASAP7_75t_L g657 ( .A(n_390), .B(n_400), .Y(n_657) );
INVx1_ASAP7_75t_L g1193 ( .A(n_390), .Y(n_1193) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx4f_ASAP7_75t_L g535 ( .A(n_391), .Y(n_535) );
INVx3_ASAP7_75t_L g744 ( .A(n_391), .Y(n_744) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g402 ( .A(n_393), .B(n_403), .Y(n_402) );
NAND2x1_ASAP7_75t_L g409 ( .A(n_393), .B(n_394), .Y(n_409) );
AND2x2_ASAP7_75t_L g414 ( .A(n_393), .B(n_394), .Y(n_414) );
INVx1_ASAP7_75t_L g422 ( .A(n_393), .Y(n_422) );
INVx2_ASAP7_75t_L g432 ( .A(n_393), .Y(n_432) );
INVx2_ASAP7_75t_L g516 ( .A(n_393), .Y(n_516) );
INVx2_ASAP7_75t_L g403 ( .A(n_394), .Y(n_403) );
BUFx2_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_394), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g515 ( .A(n_394), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g678 ( .A(n_394), .Y(n_678) );
AND2x2_ASAP7_75t_L g680 ( .A(n_394), .B(n_432), .Y(n_680) );
OR2x6_ASAP7_75t_L g743 ( .A(n_395), .B(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g1266 ( .A1(n_395), .A2(n_1267), .B1(n_1268), .B2(n_1269), .Y(n_1266) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g412 ( .A(n_396), .Y(n_412) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_396), .B(n_436), .Y(n_1285) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g417 ( .A(n_397), .Y(n_417) );
AND2x4_ASAP7_75t_L g420 ( .A(n_397), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g529 ( .A(n_397), .B(n_436), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_399), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_399), .A2(n_726), .B1(n_727), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g872 ( .A1(n_399), .A2(n_641), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_399), .A2(n_641), .B1(n_1059), .B2(n_1060), .Y(n_1102) );
INVx4_ASAP7_75t_L g1138 ( .A(n_399), .Y(n_1138) );
INVx3_ASAP7_75t_SL g1261 ( .A(n_399), .Y(n_1261) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_399), .A2(n_1355), .B1(n_1356), .B2(n_1357), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1846 ( .A1(n_399), .A2(n_641), .B1(n_1847), .B2(n_1848), .Y(n_1846) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_402), .Y(n_684) );
BUFx3_ASAP7_75t_L g758 ( .A(n_402), .Y(n_758) );
INVx2_ASAP7_75t_L g1095 ( .A(n_402), .Y(n_1095) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_407), .A2(n_813), .B1(n_822), .B2(n_835), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_407), .A2(n_809), .B1(n_828), .B2(n_835), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g1859 ( .A1(n_407), .A2(n_983), .B1(n_1837), .B2(n_1840), .C(n_1860), .Y(n_1859) );
OAI221xp5_ASAP7_75t_L g1863 ( .A1(n_407), .A2(n_1835), .B1(n_1844), .B2(n_1864), .C(n_1866), .Y(n_1863) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g519 ( .A(n_408), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_408), .A2(n_851), .B1(n_987), .B2(n_988), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_408), .A2(n_983), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
BUFx2_ASAP7_75t_SL g1123 ( .A(n_408), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1451 ( .A1(n_408), .A2(n_835), .B1(n_1435), .B2(n_1446), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g1473 ( .A1(n_408), .A2(n_1450), .B1(n_1474), .B2(n_1475), .Y(n_1473) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_409), .Y(n_525) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g571 ( .A(n_411), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g1103 ( .A(n_411), .B(n_1104), .C(n_1107), .Y(n_1103) );
INVx1_ASAP7_75t_L g1144 ( .A(n_411), .Y(n_1144) );
AOI211xp5_ASAP7_75t_L g1849 ( .A1(n_411), .A2(n_1850), .B(n_1852), .C(n_1853), .Y(n_1849) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AND2x2_ASAP7_75t_L g647 ( .A(n_412), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g651 ( .A(n_412), .B(n_418), .Y(n_651) );
OR2x2_ASAP7_75t_L g658 ( .A(n_412), .B(n_430), .Y(n_658) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_413), .Y(n_685) );
BUFx3_ASAP7_75t_L g687 ( .A(n_413), .Y(n_687) );
BUFx3_ASAP7_75t_L g759 ( .A(n_413), .Y(n_759) );
BUFx3_ASAP7_75t_L g1749 ( .A(n_413), .Y(n_1749) );
AND2x6_ASAP7_75t_L g1754 ( .A(n_413), .B(n_1755), .Y(n_1754) );
AND2x4_ASAP7_75t_SL g1760 ( .A(n_413), .B(n_1740), .Y(n_1760) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g649 ( .A(n_414), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B1(n_420), .B2(n_423), .Y(n_415) );
INVx1_ASAP7_75t_L g750 ( .A(n_416), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_416), .A2(n_653), .B1(n_931), .B2(n_932), .Y(n_930) );
BUFx3_ASAP7_75t_L g956 ( .A(n_416), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_416), .A2(n_653), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g1246 ( .A1(n_416), .A2(n_959), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g429 ( .A(n_417), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g573 ( .A(n_417), .B(n_418), .Y(n_573) );
AND2x2_ASAP7_75t_L g752 ( .A(n_417), .B(n_676), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g1262 ( .A1(n_417), .A2(n_687), .B(n_1263), .C(n_1264), .Y(n_1262) );
INVx1_ASAP7_75t_L g1268 ( .A(n_417), .Y(n_1268) );
INVx1_ASAP7_75t_L g1763 ( .A(n_418), .Y(n_1763) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_419), .A2(n_471), .B1(n_475), .B2(n_476), .Y(n_470) );
INVx2_ASAP7_75t_L g576 ( .A(n_420), .Y(n_576) );
INVx2_ASAP7_75t_L g654 ( .A(n_420), .Y(n_654) );
BUFx3_ASAP7_75t_L g959 ( .A(n_420), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_420), .A2(n_651), .B1(n_1361), .B2(n_1362), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1809 ( .A(n_421), .B(n_1755), .Y(n_1809) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g934 ( .A(n_426), .Y(n_934) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_428), .A2(n_736), .B1(n_738), .B2(n_752), .Y(n_751) );
INVxp67_ASAP7_75t_SL g802 ( .A(n_428), .Y(n_802) );
INVx2_ASAP7_75t_L g1146 ( .A(n_428), .Y(n_1146) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g864 ( .A(n_429), .Y(n_864) );
INVx1_ASAP7_75t_L g1106 ( .A(n_429), .Y(n_1106) );
INVx8_ASAP7_75t_L g509 ( .A(n_430), .Y(n_509) );
BUFx2_ASAP7_75t_L g833 ( .A(n_430), .Y(n_833) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI31xp33_ASAP7_75t_L g569 ( .A1(n_433), .A2(n_570), .A3(n_578), .B(n_579), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_433), .A2(n_724), .B1(n_739), .B2(n_740), .C(n_753), .Y(n_723) );
OAI31xp33_ASAP7_75t_L g796 ( .A1(n_433), .A2(n_797), .A3(n_801), .B(n_803), .Y(n_796) );
BUFx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g659 ( .A(n_434), .Y(n_659) );
BUFx2_ASAP7_75t_L g936 ( .A(n_434), .Y(n_936) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_434), .Y(n_1039) );
OAI31xp33_ASAP7_75t_L g1243 ( .A1(n_434), .A2(n_1244), .A3(n_1245), .B(n_1249), .Y(n_1243) );
OAI21xp5_ASAP7_75t_L g1340 ( .A1(n_434), .A2(n_1341), .B(n_1348), .Y(n_1340) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
AOI21xp5_ASAP7_75t_SL g1259 ( .A1(n_435), .A2(n_1260), .B(n_1272), .Y(n_1259) );
INVx1_ASAP7_75t_L g1514 ( .A(n_435), .Y(n_1514) );
NOR2xp33_ASAP7_75t_L g1820 ( .A(n_435), .B(n_1506), .Y(n_1820) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g1808 ( .A(n_438), .B(n_1809), .Y(n_1808) );
INVxp67_ASAP7_75t_L g1812 ( .A(n_438), .Y(n_1812) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g494 ( .A(n_439), .Y(n_494) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI31xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_458), .A3(n_478), .B(n_488), .Y(n_441) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g737 ( .A(n_444), .Y(n_737) );
BUFx2_ASAP7_75t_L g884 ( .A(n_444), .Y(n_884) );
BUFx2_ASAP7_75t_L g965 ( .A(n_444), .Y(n_965) );
OR2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .Y(n_444) );
AND2x4_ASAP7_75t_L g483 ( .A(n_445), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_445), .B(n_484), .Y(n_1215) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g454 ( .A(n_446), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g467 ( .A(n_446), .B(n_468), .Y(n_467) );
OR2x4_ASAP7_75t_L g481 ( .A(n_446), .B(n_448), .Y(n_481) );
NAND3x1_ASAP7_75t_L g562 ( .A(n_446), .B(n_563), .C(n_565), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g719 ( .A(n_446), .B(n_565), .Y(n_719) );
AND2x4_ASAP7_75t_L g1775 ( .A(n_446), .B(n_1776), .Y(n_1775) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g473 ( .A(n_447), .Y(n_473) );
NAND2xp33_ASAP7_75t_SL g541 ( .A(n_447), .B(n_491), .Y(n_541) );
INVx2_ASAP7_75t_L g545 ( .A(n_448), .Y(n_545) );
BUFx3_ASAP7_75t_L g619 ( .A(n_448), .Y(n_619) );
BUFx3_ASAP7_75t_L g998 ( .A(n_448), .Y(n_998) );
BUFx4f_ASAP7_75t_L g1168 ( .A(n_448), .Y(n_1168) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_449), .B(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_449), .Y(n_465) );
AND2x4_ASAP7_75t_L g468 ( .A(n_449), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
INVx1_ASAP7_75t_L g699 ( .A(n_450), .Y(n_699) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_453), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g583 ( .A(n_454), .Y(n_583) );
INVx2_ASAP7_75t_L g885 ( .A(n_454), .Y(n_885) );
BUFx3_ASAP7_75t_L g944 ( .A(n_454), .Y(n_944) );
INVx1_ASAP7_75t_L g554 ( .A(n_455), .Y(n_554) );
BUFx3_ASAP7_75t_L g888 ( .A(n_455), .Y(n_888) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g559 ( .A(n_456), .Y(n_559) );
INVx1_ASAP7_75t_L g464 ( .A(n_457), .Y(n_464) );
INVx2_ASAP7_75t_L g469 ( .A(n_457), .Y(n_469) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_460), .A2(n_506), .B1(n_526), .B2(n_543), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_460), .A2(n_617), .B1(n_908), .B2(n_915), .Y(n_923) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g631 ( .A(n_461), .Y(n_631) );
INVx1_ASAP7_75t_L g940 ( .A(n_461), .Y(n_940) );
INVx1_ASAP7_75t_L g1066 ( .A(n_461), .Y(n_1066) );
INVx2_ASAP7_75t_L g1294 ( .A(n_461), .Y(n_1294) );
INVx4_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_462), .Y(n_587) );
INVx3_ASAP7_75t_L g621 ( .A(n_462), .Y(n_621) );
OR2x2_ASAP7_75t_L g1807 ( .A(n_462), .B(n_1800), .Y(n_1807) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g548 ( .A(n_463), .Y(n_548) );
BUFx3_ASAP7_75t_L g790 ( .A(n_463), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
BUFx2_ASAP7_75t_L g477 ( .A(n_464), .Y(n_477) );
BUFx2_ASAP7_75t_L g474 ( .A(n_465), .Y(n_474) );
AND2x4_ASAP7_75t_L g707 ( .A(n_465), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g1211 ( .A(n_465), .Y(n_1211) );
CKINVDCx8_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_467), .B(n_662), .C(n_663), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g728 ( .A1(n_467), .A2(n_729), .B(n_730), .C(n_731), .Y(n_728) );
AOI211xp5_ASAP7_75t_L g876 ( .A1(n_467), .A2(n_869), .B(n_877), .C(n_878), .Y(n_876) );
CKINVDCx8_ASAP7_75t_R g968 ( .A(n_467), .Y(n_968) );
NOR3xp33_ASAP7_75t_L g1061 ( .A(n_467), .B(n_1062), .C(n_1064), .Y(n_1061) );
NOR3xp33_ASAP7_75t_L g1292 ( .A(n_467), .B(n_1293), .C(n_1296), .Y(n_1292) );
NOR3xp33_ASAP7_75t_L g1368 ( .A(n_467), .B(n_1369), .C(n_1371), .Y(n_1368) );
AOI211xp5_ASAP7_75t_L g1868 ( .A1(n_467), .A2(n_773), .B(n_1869), .C(n_1870), .Y(n_1868) );
INVx2_ASAP7_75t_L g701 ( .A(n_468), .Y(n_701) );
BUFx2_ASAP7_75t_L g716 ( .A(n_468), .Y(n_716) );
BUFx2_ASAP7_75t_L g730 ( .A(n_468), .Y(n_730) );
BUFx3_ASAP7_75t_L g773 ( .A(n_468), .Y(n_773) );
BUFx2_ASAP7_75t_L g892 ( .A(n_468), .Y(n_892) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_468), .Y(n_1083) );
INVx1_ASAP7_75t_L g708 ( .A(n_469), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_471), .A2(n_476), .B1(n_574), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_471), .A2(n_476), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_471), .A2(n_476), .B1(n_931), .B2(n_942), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_471), .A2(n_476), .B1(n_1035), .B2(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1065 ( .A(n_471), .Y(n_1065) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
AND2x4_ASAP7_75t_L g476 ( .A(n_472), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g666 ( .A(n_472), .B(n_474), .Y(n_666) );
AND2x2_ASAP7_75t_L g734 ( .A(n_472), .B(n_477), .Y(n_734) );
AND2x2_ASAP7_75t_L g971 ( .A(n_472), .B(n_474), .Y(n_971) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND3x4_ASAP7_75t_L g693 ( .A(n_473), .B(n_491), .C(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_473), .B(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g664 ( .A(n_476), .Y(n_664) );
BUFx6f_ASAP7_75t_L g973 ( .A(n_476), .Y(n_973) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g1297 ( .A1(n_480), .A2(n_1215), .B1(n_1267), .B2(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g668 ( .A(n_481), .Y(n_668) );
INVx2_ASAP7_75t_SL g881 ( .A(n_481), .Y(n_881) );
INVx1_ASAP7_75t_L g1043 ( .A(n_481), .Y(n_1043) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g591 ( .A(n_483), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_483), .A2(n_640), .B1(n_642), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_483), .A2(n_668), .B1(n_726), .B2(n_727), .Y(n_725) );
INVx2_ASAP7_75t_L g795 ( .A(n_483), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_483), .A2(n_873), .B1(n_874), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_483), .A2(n_668), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
INVx1_ASAP7_75t_L g1149 ( .A(n_483), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1871 ( .A1(n_483), .A2(n_668), .B1(n_1847), .B2(n_1848), .Y(n_1871) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_484), .Y(n_624) );
INVx2_ASAP7_75t_L g626 ( .A(n_484), .Y(n_626) );
INVx2_ASAP7_75t_L g704 ( .A(n_484), .Y(n_704) );
INVx1_ASAP7_75t_L g711 ( .A(n_484), .Y(n_711) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_484), .Y(n_770) );
INVx2_ASAP7_75t_L g894 ( .A(n_484), .Y(n_894) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
INVx2_ASAP7_75t_L g816 ( .A(n_485), .Y(n_816) );
BUFx8_ASAP7_75t_L g821 ( .A(n_485), .Y(n_821) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AND2x4_ASAP7_75t_L g698 ( .A(n_487), .B(n_699), .Y(n_698) );
OAI31xp33_ASAP7_75t_L g580 ( .A1(n_488), .A2(n_581), .A3(n_584), .B(n_590), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g937 ( .A1(n_488), .A2(n_938), .A3(n_939), .B(n_943), .Y(n_937) );
OAI31xp33_ASAP7_75t_L g1040 ( .A1(n_488), .A2(n_1041), .A3(n_1044), .B(n_1047), .Y(n_1040) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
AND2x2_ASAP7_75t_L g670 ( .A(n_489), .B(n_492), .Y(n_670) );
AND2x2_ASAP7_75t_SL g739 ( .A(n_489), .B(n_492), .Y(n_739) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_489), .B(n_492), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_489), .B(n_492), .Y(n_1216) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g1776 ( .A(n_491), .Y(n_1776) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g531 ( .A(n_494), .Y(n_531) );
OR2x2_ASAP7_75t_L g540 ( .A(n_494), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_494), .B(n_529), .Y(n_688) );
OR2x2_ASAP7_75t_L g1800 ( .A(n_494), .B(n_1801), .Y(n_1800) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_538), .Y(n_495) );
OAI33xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_503), .A3(n_510), .B1(n_520), .B2(n_527), .B3(n_532), .Y(n_496) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_497), .A2(n_843), .B1(n_850), .B2(n_859), .Y(n_842) );
OAI33xp33_ASAP7_75t_L g1027 ( .A1(n_497), .A2(n_989), .A3(n_1028), .B1(n_1029), .B2(n_1030), .B3(n_1031), .Y(n_1027) );
INVx1_ASAP7_75t_L g1088 ( .A(n_497), .Y(n_1088) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI33xp33_ASAP7_75t_L g1235 ( .A1(n_498), .A2(n_1194), .A3(n_1236), .B1(n_1240), .B2(n_1241), .B3(n_1242), .Y(n_1235) );
OAI33xp33_ASAP7_75t_L g1469 ( .A1(n_498), .A2(n_839), .A3(n_1470), .B1(n_1473), .B2(n_1476), .B3(n_1479), .Y(n_1469) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g599 ( .A(n_499), .Y(n_599) );
INVx4_ASAP7_75t_L g673 ( .A(n_499), .Y(n_673) );
INVx2_ASAP7_75t_L g1113 ( .A(n_499), .Y(n_1113) );
INVx2_ASAP7_75t_L g1183 ( .A(n_499), .Y(n_1183) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
OR2x6_ASAP7_75t_L g718 ( .A(n_500), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_500), .B(n_719), .Y(n_1181) );
INVx1_ASAP7_75t_L g1289 ( .A(n_500), .Y(n_1289) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g694 ( .A(n_501), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_503) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_504), .A2(n_523), .B1(n_543), .B2(n_546), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g1028 ( .A1(n_505), .A2(n_507), .B1(n_1011), .B2(n_1025), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1273 ( .A1(n_505), .A2(n_507), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_507), .A2(n_533), .B1(n_536), .B2(n_537), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_507), .A2(n_533), .B1(n_1017), .B2(n_1022), .Y(n_1031) );
INVx5_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx6_ASAP7_75t_L g598 ( .A(n_508), .Y(n_598) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g838 ( .A(n_509), .Y(n_838) );
INVx2_ASAP7_75t_L g920 ( .A(n_509), .Y(n_920) );
INVx1_ASAP7_75t_L g994 ( .A(n_509), .Y(n_994) );
INVx4_ASAP7_75t_L g1186 ( .A(n_509), .Y(n_1186) );
INVx2_ASAP7_75t_L g1239 ( .A(n_509), .Y(n_1239) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_517), .B2(n_518), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_511), .A2(n_536), .B1(n_550), .B2(n_552), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g1029 ( .A1(n_512), .A2(n_604), .B1(n_1015), .B2(n_1021), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_512), .A2(n_524), .B1(n_1012), .B2(n_1026), .Y(n_1030) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g851 ( .A(n_513), .Y(n_851) );
INVx2_ASAP7_75t_L g912 ( .A(n_513), .Y(n_912) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx3_ASAP7_75t_L g522 ( .A(n_515), .Y(n_522) );
INVx1_ASAP7_75t_L g603 ( .A(n_515), .Y(n_603) );
BUFx2_ASAP7_75t_L g835 ( .A(n_515), .Y(n_835) );
INVx2_ASAP7_75t_L g984 ( .A(n_515), .Y(n_984) );
AND2x2_ASAP7_75t_L g677 ( .A(n_516), .B(n_678), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_517), .A2(n_537), .B1(n_556), .B2(n_557), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_518), .A2(n_602), .B1(n_915), .B2(n_916), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_518), .A2(n_982), .B1(n_983), .B2(n_985), .Y(n_981) );
INVx5_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_523), .B1(n_524), .B2(n_526), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_522), .A2(n_929), .B1(n_1224), .B2(n_1234), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_522), .A2(n_1197), .B1(n_1318), .B2(n_1322), .Y(n_1329) );
INVx2_ASAP7_75t_L g1865 ( .A(n_522), .Y(n_1865) );
OAI211xp5_ASAP7_75t_SL g1281 ( .A1(n_524), .A2(n_1282), .B(n_1283), .C(n_1286), .Y(n_1281) );
OAI211xp5_ASAP7_75t_L g1765 ( .A1(n_524), .A2(n_1766), .B(n_1767), .C(n_1768), .Y(n_1765) );
BUFx4f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g605 ( .A(n_525), .Y(n_605) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
BUFx4f_ASAP7_75t_L g798 ( .A(n_525), .Y(n_798) );
BUFx6f_ASAP7_75t_L g853 ( .A(n_525), .Y(n_853) );
BUFx4f_ASAP7_75t_L g1197 ( .A(n_525), .Y(n_1197) );
OAI33xp33_ASAP7_75t_L g593 ( .A1(n_527), .A2(n_594), .A3(n_599), .B1(n_600), .B2(n_607), .B3(n_611), .Y(n_593) );
OAI33xp33_ASAP7_75t_L g906 ( .A1(n_527), .A2(n_673), .A3(n_907), .B1(n_910), .B2(n_914), .B3(n_917), .Y(n_906) );
OAI22xp5_ASAP7_75t_SL g1858 ( .A1(n_527), .A2(n_1183), .B1(n_1859), .B2(n_1863), .Y(n_1858) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_528), .B(n_765), .C(n_767), .Y(n_764) );
INVx2_ASAP7_75t_L g989 ( .A(n_528), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g1087 ( .A1(n_528), .A2(n_1088), .A3(n_1089), .B1(n_1091), .B2(n_1097), .B3(n_1098), .Y(n_1087) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_529), .B(n_530), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_529), .A2(n_645), .B1(n_1277), .B2(n_1278), .C(n_1280), .Y(n_1276) );
INVx4_ASAP7_75t_L g1751 ( .A(n_529), .Y(n_1751) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g596 ( .A(n_534), .Y(n_596) );
INVx2_ASAP7_75t_L g991 ( .A(n_534), .Y(n_991) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g1116 ( .A(n_535), .Y(n_1116) );
INVx4_ASAP7_75t_L g1185 ( .A(n_535), .Y(n_1185) );
OAI33xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_542), .A3(n_549), .B1(n_555), .B2(n_560), .B3(n_566), .Y(n_538) );
OAI33xp33_ASAP7_75t_L g1009 ( .A1(n_539), .A2(n_1010), .A3(n_1014), .B1(n_1018), .B2(n_1023), .B3(n_1024), .Y(n_1009) );
OAI33xp33_ASAP7_75t_L g1128 ( .A1(n_539), .A2(n_1129), .A3(n_1132), .B1(n_1133), .B2(n_1134), .B3(n_1135), .Y(n_1128) );
BUFx4f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx8_ASAP7_75t_L g615 ( .A(n_540), .Y(n_615) );
BUFx2_ASAP7_75t_L g806 ( .A(n_540), .Y(n_806) );
BUFx4f_ASAP7_75t_L g1165 ( .A(n_540), .Y(n_1165) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_543), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_543), .A2(n_1011), .B1(n_1012), .B2(n_1013), .Y(n_1010) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_543), .A2(n_631), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
BUFx4f_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g826 ( .A1(n_544), .A2(n_790), .B1(n_827), .B2(n_828), .Y(n_826) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g1444 ( .A(n_545), .Y(n_1444) );
OAI22xp33_ASAP7_75t_L g1135 ( .A1(n_546), .A2(n_1117), .B1(n_1124), .B2(n_1130), .Y(n_1135) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g811 ( .A(n_548), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_550), .A2(n_888), .B1(n_1120), .B2(n_1127), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_550), .A2(n_895), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_550), .A2(n_1173), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1485 ( .A1(n_550), .A2(n_818), .B1(n_1475), .B2(n_1481), .Y(n_1485) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx5_ASAP7_75t_L g556 ( .A(n_551), .Y(n_556) );
INVx3_ASAP7_75t_L g1016 ( .A(n_551), .Y(n_1016) );
INVx2_ASAP7_75t_SL g1385 ( .A(n_551), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_552), .A2(n_601), .B1(n_612), .B2(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_552), .A2(n_606), .B1(n_613), .B2(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_SL g1014 ( .A1(n_552), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
OAI21xp33_ASAP7_75t_L g1782 ( .A1(n_552), .A2(n_1783), .B(n_1784), .Y(n_1782) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1173 ( .A(n_554), .Y(n_1173) );
INVx8_ASAP7_75t_L g1020 ( .A(n_556), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_556), .A2(n_557), .B1(n_1119), .B2(n_1126), .Y(n_1132) );
OAI22xp33_ASAP7_75t_SL g925 ( .A1(n_557), .A2(n_626), .B1(n_913), .B2(n_921), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_557), .A2(n_1019), .B1(n_1021), .B2(n_1022), .Y(n_1018) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_557), .A2(n_1275), .B1(n_1282), .B2(n_1307), .C(n_1308), .Y(n_1306) );
OAI221xp5_ASAP7_75t_L g1785 ( .A1(n_557), .A2(n_1766), .B1(n_1786), .B2(n_1787), .C(n_1788), .Y(n_1785) );
CKINVDCx8_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g818 ( .A(n_558), .Y(n_818) );
INVx3_ASAP7_75t_L g895 ( .A(n_558), .Y(n_895) );
INVx3_ASAP7_75t_L g1228 ( .A(n_558), .Y(n_1228) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g824 ( .A(n_559), .Y(n_824) );
OAI33xp33_ASAP7_75t_L g996 ( .A1(n_560), .A2(n_615), .A3(n_997), .B1(n_1000), .B2(n_1002), .B3(n_1003), .Y(n_996) );
INVx1_ASAP7_75t_L g1086 ( .A(n_560), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_560), .A2(n_806), .B1(n_1300), .B2(n_1306), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1777 ( .A1(n_560), .A2(n_1778), .B1(n_1782), .B2(n_1785), .Y(n_1777) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g627 ( .A(n_561), .Y(n_627) );
INVx2_ASAP7_75t_L g1134 ( .A(n_561), .Y(n_1134) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g777 ( .A(n_562), .Y(n_777) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g1774 ( .A(n_564), .Y(n_1774) );
INVx1_ASAP7_75t_L g632 ( .A(n_567), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g568 ( .A(n_569), .B(n_580), .C(n_592), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_577), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_573), .A2(n_575), .B1(n_792), .B2(n_800), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_573), .A2(n_653), .B1(n_1200), .B2(n_1201), .Y(n_1199) );
AOI222xp33_ASAP7_75t_L g1342 ( .A1(n_573), .A2(n_687), .B1(n_959), .B2(n_1337), .C1(n_1338), .C2(n_1343), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_573), .A2(n_653), .B1(n_1417), .B2(n_1424), .Y(n_1423) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g1142 ( .A(n_576), .Y(n_1142) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g1166 ( .A1(n_587), .A2(n_1167), .B1(n_1168), .B2(n_1169), .Y(n_1166) );
OAI22xp33_ASAP7_75t_L g1324 ( .A1(n_587), .A2(n_1168), .B1(n_1325), .B2(n_1326), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1483 ( .A1(n_587), .A2(n_1444), .B1(n_1471), .B2(n_1477), .Y(n_1483) );
OAI22xp33_ASAP7_75t_L g1831 ( .A1(n_587), .A2(n_1832), .B1(n_1833), .B2(n_1835), .Y(n_1831) );
NOR2xp33_ASAP7_75t_SL g592 ( .A(n_593), .B(n_614), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_595), .A2(n_608), .B1(n_617), .B2(n_620), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_596), .A2(n_598), .B1(n_612), .B2(n_613), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g907 ( .A1(n_596), .A2(n_838), .B1(n_908), .B2(n_909), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_597), .A2(n_609), .B1(n_629), .B2(n_631), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_598), .A2(n_918), .B1(n_979), .B2(n_980), .Y(n_978) );
OAI22xp5_ASAP7_75t_SL g1114 ( .A1(n_598), .A2(n_1115), .B1(n_1116), .B2(n_1117), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_598), .A2(n_918), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_606), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_602), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_602), .A2(n_798), .B1(n_844), .B2(n_845), .C(n_846), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_602), .A2(n_853), .B1(n_1316), .B2(n_1326), .Y(n_1330) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g1188 ( .A(n_603), .Y(n_1188) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g645 ( .A(n_605), .Y(n_645) );
INVx2_ASAP7_75t_L g929 ( .A(n_605), .Y(n_929) );
INVx2_ASAP7_75t_L g1189 ( .A(n_605), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_610), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
INVx1_ASAP7_75t_L g954 ( .A(n_610), .Y(n_954) );
OAI33xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .A3(n_622), .B1(n_625), .B2(n_627), .B3(n_628), .Y(n_614) );
OAI33xp33_ASAP7_75t_L g922 ( .A1(n_615), .A2(n_627), .A3(n_923), .B1(n_924), .B2(n_925), .B3(n_926), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g1781 ( .A(n_615), .Y(n_1781) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_617), .A2(n_620), .B1(n_909), .B2(n_916), .Y(n_926) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g630 ( .A(n_619), .Y(n_630) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_619), .Y(n_1131) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g1223 ( .A(n_621), .Y(n_1223) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g1001 ( .A(n_624), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_629), .A2(n_631), .B1(n_980), .B2(n_988), .Y(n_1003) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_901), .B1(n_902), .B2(n_945), .Y(n_633) );
INVx1_ASAP7_75t_L g945 ( .A(n_634), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_781), .B1(n_782), .B2(n_900), .Y(n_634) );
INVx1_ASAP7_75t_L g900 ( .A(n_635), .Y(n_900) );
XNOR2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_722), .Y(n_635) );
INVx1_ASAP7_75t_L g720 ( .A(n_637), .Y(n_720) );
NAND4xp75_ASAP7_75t_L g637 ( .A(n_638), .B(n_660), .C(n_671), .D(n_692), .Y(n_637) );
AO21x1_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_643), .B(n_659), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_641), .B(n_1514), .Y(n_1513) );
AND2x4_ASAP7_75t_SL g1819 ( .A(n_641), .B(n_1820), .Y(n_1819) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_656), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g866 ( .A(n_646), .B(n_867), .C(n_870), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g1359 ( .A(n_646), .B(n_1360), .C(n_1363), .Y(n_1359) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI211xp5_ASAP7_75t_L g745 ( .A1(n_647), .A2(n_746), .B(n_748), .C(n_749), .Y(n_745) );
INVx2_ASAP7_75t_L g1198 ( .A(n_647), .Y(n_1198) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g747 ( .A(n_649), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_655), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_651), .A2(n_653), .B1(n_868), .B2(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g1265 ( .A(n_651), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_651), .A2(n_653), .B1(n_1456), .B2(n_1457), .Y(n_1455) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_651), .A2(n_959), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_652), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g1347 ( .A(n_658), .Y(n_1347) );
AOI21xp33_ASAP7_75t_L g860 ( .A1(n_659), .A2(n_861), .B(n_872), .Y(n_860) );
AO21x1_ASAP7_75t_L g1101 ( .A1(n_659), .A2(n_1102), .B(n_1103), .Y(n_1101) );
AO21x1_ASAP7_75t_L g1353 ( .A1(n_659), .A2(n_1354), .B(n_1358), .Y(n_1353) );
AOI31xp33_ASAP7_75t_SL g1845 ( .A1(n_659), .A2(n_1846), .A3(n_1849), .B(n_1854), .Y(n_1845) );
AO21x1_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_667), .B(n_669), .Y(n_660) );
INVx1_ASAP7_75t_L g732 ( .A(n_666), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g1254 ( .A1(n_666), .A2(n_1208), .B1(n_1247), .B2(n_1255), .Y(n_1254) );
AOI222xp33_ASAP7_75t_L g1335 ( .A1(n_666), .A2(n_734), .B1(n_892), .B2(n_1336), .C1(n_1337), .C2(n_1338), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_666), .B(n_1361), .Y(n_1370) );
AOI22xp33_ASAP7_75t_SL g1416 ( .A1(n_666), .A2(n_734), .B1(n_1417), .B2(n_1418), .Y(n_1416) );
AOI22xp33_ASAP7_75t_SL g1463 ( .A1(n_666), .A2(n_734), .B1(n_1456), .B2(n_1464), .Y(n_1463) );
AOI22xp33_ASAP7_75t_SL g1497 ( .A1(n_666), .A2(n_734), .B1(n_1490), .B2(n_1498), .Y(n_1497) );
AOI22xp5_ASAP7_75t_L g1367 ( .A1(n_668), .A2(n_1215), .B1(n_1355), .B2(n_1357), .Y(n_1367) );
AOI31xp33_ASAP7_75t_L g875 ( .A1(n_669), .A2(n_876), .A3(n_880), .B(n_882), .Y(n_875) );
AO21x1_ASAP7_75t_L g1366 ( .A1(n_669), .A2(n_1367), .B(n_1368), .Y(n_1366) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI31xp33_ASAP7_75t_L g785 ( .A1(n_670), .A2(n_786), .A3(n_787), .B(n_794), .Y(n_785) );
AOI33xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .A3(n_681), .B1(n_686), .B2(n_688), .B3(n_689), .Y(n_671) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_672), .Y(n_763) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
OAI33xp33_ASAP7_75t_L g829 ( .A1(n_673), .A2(n_830), .A3(n_834), .B1(n_836), .B2(n_837), .B3(n_839), .Y(n_829) );
OAI33xp33_ASAP7_75t_L g977 ( .A1(n_673), .A2(n_978), .A3(n_981), .B1(n_986), .B2(n_989), .B3(n_990), .Y(n_977) );
INVx2_ASAP7_75t_SL g1373 ( .A(n_673), .Y(n_1373) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g691 ( .A(n_676), .Y(n_691) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g762 ( .A(n_677), .Y(n_762) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_677), .B(n_1740), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1803 ( .A(n_677), .B(n_1755), .Y(n_1803) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_679), .Y(n_1090) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g849 ( .A(n_680), .Y(n_849) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_680), .Y(n_858) );
BUFx3_ASAP7_75t_L g1753 ( .A(n_680), .Y(n_1753) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_684), .Y(n_766) );
INVx2_ASAP7_75t_L g1377 ( .A(n_684), .Y(n_1377) );
AND2x4_ASAP7_75t_L g1746 ( .A(n_684), .B(n_1740), .Y(n_1746) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_685), .B(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g1851 ( .A(n_685), .Y(n_1851) );
INVx2_ASAP7_75t_L g839 ( .A(n_688), .Y(n_839) );
INVx2_ASAP7_75t_L g1194 ( .A(n_688), .Y(n_1194) );
AOI33xp33_ASAP7_75t_L g1372 ( .A1(n_688), .A2(n_1373), .A3(n_1374), .B1(n_1375), .B2(n_1379), .B3(n_1380), .Y(n_1372) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
AOI33xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .A3(n_702), .B1(n_709), .B2(n_713), .B3(n_717), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_693), .B(n_769), .C(n_772), .Y(n_768) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_693), .Y(n_1070) );
INVx1_ASAP7_75t_L g1390 ( .A(n_693), .Y(n_1390) );
INVx1_ASAP7_75t_L g1770 ( .A(n_694), .Y(n_1770) );
BUFx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g780 ( .A(n_697), .Y(n_780) );
BUFx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx8_ASAP7_75t_L g715 ( .A(n_698), .Y(n_715) );
BUFx3_ASAP7_75t_L g1075 ( .A(n_698), .Y(n_1075) );
NAND2x1p5_ASAP7_75t_L g1811 ( .A(n_698), .B(n_1775), .Y(n_1811) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g877 ( .A(n_701), .Y(n_877) );
INVx2_ASAP7_75t_L g1076 ( .A(n_701), .Y(n_1076) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_704), .A2(n_844), .B1(n_888), .B2(n_889), .C(n_890), .Y(n_887) );
INVx2_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g712 ( .A(n_706), .Y(n_712) );
INVx1_ASAP7_75t_L g1080 ( .A(n_706), .Y(n_1080) );
INVx5_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
BUFx12f_ASAP7_75t_L g771 ( .A(n_707), .Y(n_771) );
BUFx2_ASAP7_75t_L g1305 ( .A(n_707), .Y(n_1305) );
INVx1_ASAP7_75t_L g1209 ( .A(n_708), .Y(n_1209) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx8_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g891 ( .A(n_715), .Y(n_891) );
INVx2_ASAP7_75t_L g1309 ( .A(n_715), .Y(n_1309) );
INVx2_ASAP7_75t_L g1815 ( .A(n_715), .Y(n_1815) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g805 ( .A1(n_718), .A2(n_806), .A3(n_807), .B1(n_812), .B2(n_819), .B3(n_826), .Y(n_805) );
OAI33xp33_ASAP7_75t_L g1313 ( .A1(n_718), .A2(n_806), .A3(n_1314), .B1(n_1317), .B2(n_1320), .B3(n_1324), .Y(n_1313) );
INVx1_ASAP7_75t_L g1387 ( .A(n_718), .Y(n_1387) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .C(n_735), .Y(n_724) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g879 ( .A(n_734), .Y(n_879) );
AOI32xp33_ASAP7_75t_L g1207 ( .A1(n_734), .A2(n_1201), .A3(n_1208), .B1(n_1210), .B2(n_1212), .Y(n_1207) );
INVxp67_ASAP7_75t_L g1295 ( .A(n_734), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1872 ( .A1(n_737), .A2(n_885), .B1(n_1855), .B2(n_1856), .Y(n_1872) );
OAI31xp33_ASAP7_75t_L g963 ( .A1(n_739), .A2(n_964), .A3(n_967), .B(n_974), .Y(n_963) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_739), .Y(n_1155) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_739), .A2(n_1291), .B(n_1299), .Y(n_1290) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .C(n_751), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g1356 ( .A(n_743), .Y(n_1356) );
INVx2_ASAP7_75t_SL g832 ( .A(n_744), .Y(n_832) );
BUFx3_ASAP7_75t_L g918 ( .A(n_744), .Y(n_918) );
BUFx3_ASAP7_75t_L g1237 ( .A(n_744), .Y(n_1237) );
BUFx6f_ASAP7_75t_L g1332 ( .A(n_744), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_746), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g1096 ( .A(n_747), .Y(n_1096) );
INVx2_ASAP7_75t_L g1378 ( .A(n_747), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g861 ( .A1(n_752), .A2(n_862), .B1(n_863), .B2(n_865), .C(n_866), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_752), .A2(n_1345), .B1(n_1346), .B2(n_1347), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g1854 ( .A1(n_752), .A2(n_1855), .B1(n_1856), .B2(n_1857), .Y(n_1854) );
NAND4xp25_ASAP7_75t_L g753 ( .A(n_754), .B(n_764), .C(n_768), .D(n_774), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_760), .C(n_763), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g847 ( .A(n_762), .Y(n_847) );
INVx2_ASAP7_75t_SL g1099 ( .A(n_762), .Y(n_1099) );
INVx2_ASAP7_75t_L g1287 ( .A(n_762), .Y(n_1287) );
INVx1_ASAP7_75t_L g1381 ( .A(n_762), .Y(n_1381) );
INVx2_ASAP7_75t_L g1861 ( .A(n_762), .Y(n_1861) );
INVx2_ASAP7_75t_SL g1302 ( .A(n_770), .Y(n_1302) );
INVx2_ASAP7_75t_L g1786 ( .A(n_770), .Y(n_1786) );
NAND3xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .C(n_778), .Y(n_774) );
INVx1_ASAP7_75t_L g1023 ( .A(n_776), .Y(n_1023) );
BUFx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
BUFx2_ASAP7_75t_L g899 ( .A(n_777), .Y(n_899) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_840), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_796), .C(n_804), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_788), .A2(n_1115), .B1(n_1122), .B2(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_790), .Y(n_999) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_790), .A2(n_1168), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_790), .A2(n_1168), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_790), .A2(n_1168), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
BUFx6f_ASAP7_75t_L g1415 ( .A(n_790), .Y(n_1415) );
OAI22xp33_ASAP7_75t_L g1443 ( .A1(n_790), .A2(n_1444), .B1(n_1445), .B2(n_1446), .Y(n_1443) );
OAI22xp33_ASAP7_75t_L g1486 ( .A1(n_790), .A2(n_1444), .B1(n_1472), .B2(n_1478), .Y(n_1486) );
OAI22xp5_ASAP7_75t_L g1240 ( .A1(n_798), .A2(n_1188), .B1(n_1226), .B2(n_1230), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1409 ( .A1(n_798), .A2(n_835), .B1(n_1396), .B2(n_1405), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_829), .Y(n_804) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_806), .A2(n_887), .B1(n_893), .B2(n_898), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_808), .A2(n_827), .B1(n_831), .B2(n_833), .Y(n_830) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
INVxp67_ASAP7_75t_SL g1013 ( .A(n_811), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .B1(n_817), .B2(n_818), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_814), .A2(n_888), .B1(n_911), .B2(n_919), .Y(n_924) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g1441 ( .A(n_815), .Y(n_1441) );
INVx3_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_816), .Y(n_1079) );
INVx1_ASAP7_75t_L g1085 ( .A(n_816), .Y(n_1085) );
BUFx2_ASAP7_75t_L g1307 ( .A(n_816), .Y(n_1307) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_817), .A2(n_825), .B1(n_831), .B2(n_838), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_818), .A2(n_1321), .B1(n_1322), .B2(n_1323), .Y(n_1320) );
OAI22xp5_ASAP7_75t_L g1836 ( .A1(n_818), .A2(n_1385), .B1(n_1837), .B2(n_1838), .Y(n_1836) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_822), .B1(n_823), .B2(n_825), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g1839 ( .A1(n_820), .A2(n_823), .B1(n_1840), .B2(n_1841), .Y(n_1839) );
INVx2_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_SL g1172 ( .A(n_821), .Y(n_1172) );
INVx3_ASAP7_75t_L g1321 ( .A(n_821), .Y(n_1321) );
INVx3_ASAP7_75t_L g1779 ( .A(n_821), .Y(n_1779) );
AND2x4_ASAP7_75t_L g1817 ( .A(n_821), .B(n_1816), .Y(n_1817) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_823), .A2(n_1016), .B1(n_1176), .B2(n_1177), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_823), .A2(n_1307), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OR2x2_ASAP7_75t_L g1799 ( .A(n_824), .B(n_1800), .Y(n_1799) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_838), .A2(n_1185), .B1(n_1471), .B2(n_1472), .Y(n_1470) );
OAI33xp33_ASAP7_75t_L g1447 ( .A1(n_839), .A2(n_1183), .A3(n_1448), .B1(n_1449), .B2(n_1451), .B3(n_1452), .Y(n_1447) );
NOR4xp25_ASAP7_75t_L g841 ( .A(n_842), .B(n_860), .C(n_875), .D(n_886), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g893 ( .A1(n_845), .A2(n_894), .B1(n_895), .B2(n_896), .C(n_897), .Y(n_893) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_848), .B(n_1740), .Y(n_1739) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g1100 ( .A(n_849), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_853), .B2(n_854), .C(n_855), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_851), .A2(n_1122), .B1(n_1123), .B2(n_1124), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1476 ( .A1(n_853), .A2(n_1450), .B1(n_1477), .B2(n_1478), .Y(n_1476) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx2_ASAP7_75t_L g1862 ( .A(n_858), .Y(n_1862) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_862), .A2(n_865), .B1(n_883), .B2(n_885), .Y(n_882) );
INVx2_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_864), .Y(n_961) );
INVx2_ASAP7_75t_L g975 ( .A(n_881), .Y(n_975) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g966 ( .A(n_885), .Y(n_966) );
INVx2_ASAP7_75t_L g1063 ( .A(n_885), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_888), .A2(n_982), .B1(n_992), .B2(n_1001), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_888), .A2(n_894), .B1(n_985), .B2(n_995), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_894), .A2(n_1226), .B1(n_1227), .B2(n_1228), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1436 ( .A1(n_894), .A2(n_1228), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
OAI22xp5_ASAP7_75t_L g1484 ( .A1(n_894), .A2(n_1228), .B1(n_1474), .B2(n_1480), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_895), .A2(n_1016), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NAND3xp33_ASAP7_75t_L g904 ( .A(n_905), .B(n_927), .C(n_937), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_922), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_917) );
OAI31xp33_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_933), .A3(n_935), .B(n_936), .Y(n_927) );
OAI31xp33_ASAP7_75t_L g951 ( .A1(n_936), .A2(n_952), .A3(n_960), .B(n_962), .Y(n_951) );
OAI31xp33_ASAP7_75t_L g1195 ( .A1(n_936), .A2(n_1196), .A3(n_1202), .B(n_1203), .Y(n_1195) );
OAI31xp33_ASAP7_75t_SL g1420 ( .A1(n_936), .A2(n_1421), .A3(n_1422), .B(n_1425), .Y(n_1420) );
OAI31xp33_ASAP7_75t_L g1453 ( .A1(n_936), .A2(n_1454), .A3(n_1458), .B(n_1459), .Y(n_1453) );
OAI31xp33_ASAP7_75t_L g1487 ( .A1(n_936), .A2(n_1488), .A3(n_1492), .B(n_1493), .Y(n_1487) );
INVx1_ASAP7_75t_L g1048 ( .A(n_946), .Y(n_1048) );
XNOR2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_1004), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g950 ( .A(n_951), .B(n_963), .C(n_976), .Y(n_950) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_957), .B1(n_958), .B2(n_959), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_956), .A2(n_1141), .B1(n_1142), .B2(n_1143), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_957), .A2(n_970), .B1(n_972), .B2(n_973), .Y(n_969) );
BUFx3_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
BUFx3_ASAP7_75t_L g1152 ( .A(n_971), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_973), .A2(n_1141), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
NOR2xp33_ASAP7_75t_SL g976 ( .A(n_977), .B(n_996), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g997 ( .A1(n_979), .A2(n_987), .B1(n_998), .B2(n_999), .Y(n_997) );
INVx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
BUFx2_ASAP7_75t_L g1279 ( .A(n_984), .Y(n_1279) );
INVx2_ASAP7_75t_L g1450 ( .A(n_984), .Y(n_1450) );
OAI33xp33_ASAP7_75t_L g1112 ( .A1(n_989), .A2(n_1113), .A3(n_1114), .B1(n_1118), .B2(n_1121), .B3(n_1125), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B1(n_993), .B2(n_995), .Y(n_990) );
BUFx3_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI22xp33_ASAP7_75t_L g1408 ( .A1(n_994), .A2(n_1185), .B1(n_1399), .B2(n_1402), .Y(n_1408) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1032), .C(n_1040), .Y(n_1007) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1027), .Y(n_1008) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g1829 ( .A1(n_1023), .A2(n_1830), .A3(n_1831), .B1(n_1836), .B2(n_1839), .B3(n_1842), .Y(n_1829) );
OAI31xp33_ASAP7_75t_SL g1032 ( .A1(n_1033), .A2(n_1037), .A3(n_1038), .B(n_1039), .Y(n_1032) );
OAI31xp33_ASAP7_75t_L g1136 ( .A1(n_1039), .A2(n_1137), .A3(n_1139), .B(n_1145), .Y(n_1136) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1158), .B1(n_1501), .B2(n_1502), .Y(n_1050) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1051), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1108), .B1(n_1109), .B2(n_1156), .Y(n_1051) );
INVxp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1055), .Y(n_1157) );
NAND4xp25_ASAP7_75t_SL g1056 ( .A(n_1057), .B(n_1069), .C(n_1087), .D(n_1101), .Y(n_1056) );
AO21x1_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1061), .B(n_1067), .Y(n_1057) );
AOI31xp33_ASAP7_75t_L g1867 ( .A1(n_1067), .A2(n_1868), .A3(n_1871), .B(n_1872), .Y(n_1867) );
CKINVDCx14_ASAP7_75t_R g1067 ( .A(n_1068), .Y(n_1067) );
AOI33xp33_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1071), .A3(n_1077), .B1(n_1081), .B2(n_1084), .B3(n_1086), .Y(n_1069) );
BUFx2_ASAP7_75t_SL g1072 ( .A(n_1073), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1772 ( .A(n_1083), .B(n_1773), .Y(n_1772) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_L g1857 ( .A(n_1105), .Y(n_1857) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
NAND2xp5_ASAP7_75t_SL g1270 ( .A(n_1106), .B(n_1271), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1108 ( .A(n_1109), .Y(n_1108) );
NAND3xp33_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1136), .C(n_1147), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1128), .Y(n_1111) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
OAI31xp33_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1150), .A3(n_1154), .B(n_1155), .Y(n_1147) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1158), .Y(n_1502) );
XOR2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1349), .Y(n_1158) );
XNOR2xp5_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1256), .Y(n_1159) );
XNOR2xp5_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1217), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1195), .C(n_1204), .Y(n_1162) );
NOR2xp33_ASAP7_75t_SL g1163 ( .A(n_1164), .B(n_1182), .Y(n_1163) );
OAI33xp33_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1166), .A3(n_1170), .B1(n_1175), .B2(n_1178), .B3(n_1181), .Y(n_1164) );
OAI33xp33_ASAP7_75t_L g1220 ( .A1(n_1165), .A2(n_1181), .A3(n_1221), .B1(n_1225), .B2(n_1229), .B3(n_1232), .Y(n_1220) );
OAI33xp33_ASAP7_75t_L g1394 ( .A1(n_1165), .A2(n_1181), .A3(n_1395), .B1(n_1398), .B2(n_1401), .B3(n_1404), .Y(n_1394) );
OAI33xp33_ASAP7_75t_L g1432 ( .A1(n_1165), .A2(n_1181), .A3(n_1433), .B1(n_1436), .B2(n_1439), .B3(n_1443), .Y(n_1432) );
OAI33xp33_ASAP7_75t_L g1482 ( .A1(n_1165), .A2(n_1181), .A3(n_1483), .B1(n_1484), .B2(n_1485), .B3(n_1486), .Y(n_1482) );
BUFx3_ASAP7_75t_L g1830 ( .A(n_1165), .Y(n_1830) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_1167), .A2(n_1179), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1168), .A2(n_1222), .B1(n_1223), .B2(n_1224), .Y(n_1221) );
OAI22xp33_ASAP7_75t_L g1314 ( .A1(n_1168), .A2(n_1294), .B1(n_1315), .B2(n_1316), .Y(n_1314) );
OAI22xp5_ASAP7_75t_SL g1398 ( .A1(n_1168), .A2(n_1223), .B1(n_1399), .B2(n_1400), .Y(n_1398) );
OAI22xp5_ASAP7_75t_L g1433 ( .A1(n_1168), .A2(n_1223), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1169), .A2(n_1180), .B1(n_1188), .B2(n_1189), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1171), .A2(n_1176), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1439 ( .A1(n_1173), .A2(n_1440), .B1(n_1441), .B2(n_1442), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_1174), .A2(n_1177), .B1(n_1186), .B2(n_1192), .Y(n_1191) );
OAI33xp33_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1184), .A3(n_1187), .B1(n_1190), .B2(n_1191), .B3(n_1194), .Y(n_1182) );
OAI33xp33_ASAP7_75t_L g1327 ( .A1(n_1183), .A2(n_1194), .A3(n_1328), .B1(n_1329), .B2(n_1330), .B3(n_1331), .Y(n_1327) );
OAI33xp33_ASAP7_75t_L g1407 ( .A1(n_1183), .A2(n_1194), .A3(n_1408), .B1(n_1409), .B2(n_1410), .B3(n_1411), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_1185), .A2(n_1186), .B1(n_1397), .B2(n_1406), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_1185), .A2(n_1238), .B1(n_1434), .B2(n_1445), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_1185), .A2(n_1186), .B1(n_1438), .B2(n_1442), .Y(n_1452) );
OAI22xp5_ASAP7_75t_L g1479 ( .A1(n_1185), .A2(n_1238), .B1(n_1480), .B2(n_1481), .Y(n_1479) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_1186), .A2(n_1227), .B1(n_1231), .B2(n_1237), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_1186), .A2(n_1237), .B1(n_1315), .B2(n_1325), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g1410 ( .A1(n_1188), .A2(n_1189), .B1(n_1400), .B2(n_1403), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g1449 ( .A1(n_1189), .A2(n_1437), .B1(n_1440), .B2(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
NAND3xp33_ASAP7_75t_SL g1341 ( .A(n_1198), .B(n_1342), .C(n_1344), .Y(n_1341) );
OAI31xp33_ASAP7_75t_SL g1204 ( .A1(n_1205), .A2(n_1206), .A3(n_1213), .B(n_1216), .Y(n_1204) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1209), .Y(n_1795) );
AND2x4_ASAP7_75t_SL g1791 ( .A(n_1210), .B(n_1773), .Y(n_1791) );
INVx3_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
OAI31xp33_ASAP7_75t_SL g1250 ( .A1(n_1216), .A2(n_1251), .A3(n_1252), .B(n_1253), .Y(n_1250) );
OAI21xp5_ASAP7_75t_L g1333 ( .A1(n_1216), .A2(n_1334), .B(n_1339), .Y(n_1333) );
OAI31xp33_ASAP7_75t_L g1412 ( .A1(n_1216), .A2(n_1413), .A3(n_1414), .B(n_1419), .Y(n_1412) );
OAI31xp33_ASAP7_75t_SL g1460 ( .A1(n_1216), .A2(n_1461), .A3(n_1462), .B(n_1465), .Y(n_1460) );
OAI31xp33_ASAP7_75t_SL g1494 ( .A1(n_1216), .A2(n_1495), .A3(n_1496), .B(n_1499), .Y(n_1494) );
NAND3xp33_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1243), .C(n_1250), .Y(n_1218) );
NOR2xp33_ASAP7_75t_SL g1219 ( .A(n_1220), .B(n_1235), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1222), .A2(n_1233), .B1(n_1237), .B2(n_1238), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_1238), .A2(n_1319), .B1(n_1323), .B2(n_1332), .Y(n_1331) );
BUFx6f_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
XOR2xp5_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1310), .Y(n_1256) );
OAI21xp5_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1288), .B(n_1290), .Y(n_1258) );
OAI21xp5_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1276), .B(n_1281), .Y(n_1272) );
INVx4_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
BUFx2_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_SL g1291 ( .A(n_1292), .B(n_1297), .Y(n_1291) );
OAI211xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B(n_1303), .C(n_1304), .Y(n_1300) );
NAND3xp33_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1333), .C(n_1340), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1327), .Y(n_1312) );
AOI22xp5_ASAP7_75t_L g1349 ( .A1(n_1350), .A2(n_1426), .B1(n_1427), .B2(n_1500), .Y(n_1349) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1350), .Y(n_1500) );
XNOR2x1_ASAP7_75t_SL g1350 ( .A(n_1351), .B(n_1391), .Y(n_1350) );
NAND4xp75_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1366), .C(n_1372), .D(n_1382), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1365), .Y(n_1358) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_L g1750 ( .A(n_1377), .Y(n_1750) );
AOI32xp33_ASAP7_75t_L g1382 ( .A1(n_1383), .A2(n_1386), .A3(n_1387), .B1(n_1388), .B2(n_1389), .Y(n_1382) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
AND3x1_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1412), .C(n_1420), .Y(n_1392) );
NOR2xp33_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1407), .Y(n_1393) );
OAI22xp33_ASAP7_75t_L g1842 ( .A1(n_1415), .A2(n_1444), .B1(n_1843), .B2(n_1844), .Y(n_1842) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
XNOR2x1_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1466), .Y(n_1427) );
XNOR2xp5_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1430), .Y(n_1428) );
AND3x1_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1453), .C(n_1460), .Y(n_1430) );
NOR2xp33_ASAP7_75t_SL g1431 ( .A(n_1432), .B(n_1447), .Y(n_1431) );
INVx2_ASAP7_75t_SL g1834 ( .A(n_1444), .Y(n_1834) );
AND3x1_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1487), .C(n_1494), .Y(n_1467) );
NOR2xp33_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1482), .Y(n_1468) );
BUFx3_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx3_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1512), .Y(n_1505) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
NOR2xp33_ASAP7_75t_L g1507 ( .A(n_1508), .B(n_1510), .Y(n_1507) );
NOR2xp33_ASAP7_75t_L g1824 ( .A(n_1508), .B(n_1511), .Y(n_1824) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1508), .Y(n_1877) );
HB1xp67_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
NOR2xp33_ASAP7_75t_L g1879 ( .A(n_1511), .B(n_1877), .Y(n_1879) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
OAI221xp5_ASAP7_75t_L g1515 ( .A1(n_1516), .A2(n_1731), .B1(n_1733), .B2(n_1818), .C(n_1821), .Y(n_1515) );
NOR3xp33_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1711), .C(n_1725), .Y(n_1516) );
OAI221xp5_ASAP7_75t_L g1517 ( .A1(n_1518), .A2(n_1610), .B1(n_1632), .B2(n_1668), .C(n_1669), .Y(n_1517) );
OAI21xp5_ASAP7_75t_SL g1518 ( .A1(n_1519), .A2(n_1556), .B(n_1604), .Y(n_1518) );
OAI22xp5_ASAP7_75t_L g1727 ( .A1(n_1519), .A2(n_1583), .B1(n_1656), .B2(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
NAND2xp5_ASAP7_75t_SL g1520 ( .A(n_1521), .B(n_1551), .Y(n_1520) );
AOI211xp5_ASAP7_75t_L g1719 ( .A1(n_1521), .A2(n_1597), .B(n_1720), .C(n_1721), .Y(n_1719) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
OR2x2_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1538), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1523), .B(n_1576), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1523), .B(n_1599), .Y(n_1615) );
CKINVDCx5p33_ASAP7_75t_R g1623 ( .A(n_1523), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1523), .B(n_1635), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1523), .B(n_1655), .Y(n_1654) );
OAI21xp5_ASAP7_75t_SL g1724 ( .A1(n_1523), .A2(n_1655), .B(n_1721), .Y(n_1724) );
INVx4_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
OR2x2_ASAP7_75t_L g1603 ( .A(n_1524), .B(n_1567), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1524), .B(n_1612), .Y(n_1611) );
INVx4_ASAP7_75t_L g1620 ( .A(n_1524), .Y(n_1620) );
NOR2xp33_ASAP7_75t_L g1626 ( .A(n_1524), .B(n_1569), .Y(n_1626) );
NOR2xp33_ASAP7_75t_L g1630 ( .A(n_1524), .B(n_1631), .Y(n_1630) );
AOI322xp5_ASAP7_75t_L g1636 ( .A1(n_1524), .A2(n_1637), .A3(n_1639), .B1(n_1641), .B2(n_1643), .C1(n_1644), .C2(n_1646), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1524), .B(n_1572), .Y(n_1643) );
NAND2xp5_ASAP7_75t_SL g1663 ( .A(n_1524), .B(n_1567), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1524), .B(n_1551), .Y(n_1710) );
AND2x4_ASAP7_75t_SL g1524 ( .A(n_1525), .B(n_1533), .Y(n_1524) );
AND2x4_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1528), .Y(n_1526) );
AND2x6_ASAP7_75t_L g1531 ( .A(n_1527), .B(n_1532), .Y(n_1531) );
AND2x6_ASAP7_75t_L g1534 ( .A(n_1527), .B(n_1535), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1527), .B(n_1537), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1527), .B(n_1537), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1527), .B(n_1528), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1527), .B(n_1537), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1530), .Y(n_1528) );
INVx2_ASAP7_75t_L g1592 ( .A(n_1531), .Y(n_1592) );
HB1xp67_ASAP7_75t_L g1876 ( .A(n_1532), .Y(n_1876) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1538), .Y(n_1720) );
OR2x2_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1543), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1539), .B(n_1572), .Y(n_1571) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_1539), .B(n_1581), .Y(n_1580) );
OR2x2_ASAP7_75t_L g1680 ( .A(n_1539), .B(n_1545), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1539), .B(n_1626), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1541), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1567 ( .A(n_1540), .B(n_1541), .Y(n_1567) );
OR2x2_ASAP7_75t_L g1616 ( .A(n_1543), .B(n_1566), .Y(n_1616) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1543), .Y(n_1648) );
OR2x2_ASAP7_75t_L g1662 ( .A(n_1543), .B(n_1663), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_1543), .B(n_1697), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1548), .Y(n_1543) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1545), .B(n_1548), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1545), .B(n_1573), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1545), .B(n_1548), .Y(n_1576) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1545), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_1545), .B(n_1567), .Y(n_1667) );
NAND3xp33_ASAP7_75t_L g1671 ( .A(n_1545), .B(n_1587), .C(n_1607), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1547), .Y(n_1545) );
INVx2_ASAP7_75t_L g1573 ( .A(n_1548), .Y(n_1573) );
OR2x2_ASAP7_75t_L g1707 ( .A(n_1548), .B(n_1567), .Y(n_1707) );
NAND2x1p5_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1550), .Y(n_1548) );
AOI221xp5_ASAP7_75t_L g1610 ( .A1(n_1551), .A2(n_1583), .B1(n_1611), .B2(n_1613), .C(n_1624), .Y(n_1610) );
NAND2xp5_ASAP7_75t_L g1729 ( .A(n_1551), .B(n_1622), .Y(n_1729) );
INVx2_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1552), .B(n_1559), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1552), .B(n_1620), .Y(n_1666) );
OAI322xp33_ASAP7_75t_L g1681 ( .A1(n_1552), .A2(n_1564), .A3(n_1604), .B1(n_1682), .B2(n_1685), .C1(n_1686), .C2(n_1689), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1693 ( .A(n_1552), .B(n_1606), .Y(n_1693) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1578 ( .A(n_1553), .B(n_1559), .Y(n_1578) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1553), .Y(n_1600) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
OAI211xp5_ASAP7_75t_L g1556 ( .A1(n_1557), .A2(n_1563), .B(n_1574), .C(n_1596), .Y(n_1556) );
NOR2xp33_ASAP7_75t_L g1661 ( .A(n_1557), .B(n_1662), .Y(n_1661) );
OAI21xp5_ASAP7_75t_L g1730 ( .A1(n_1557), .A2(n_1578), .B(n_1644), .Y(n_1730) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
AOI21xp5_ASAP7_75t_L g1629 ( .A1(n_1558), .A2(n_1586), .B(n_1630), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1558), .B(n_1601), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1558), .B(n_1674), .Y(n_1673) );
INVx2_ASAP7_75t_L g1583 ( .A(n_1559), .Y(n_1583) );
OAI21xp33_ASAP7_75t_L g1584 ( .A1(n_1559), .A2(n_1585), .B(n_1586), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1559), .B(n_1607), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1656 ( .A(n_1559), .B(n_1600), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1685 ( .A(n_1559), .B(n_1607), .Y(n_1685) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1559), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1559), .B(n_1606), .Y(n_1723) );
INVx2_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1560), .B(n_1600), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1562), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1570), .Y(n_1563) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1565), .B(n_1623), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1566), .B(n_1568), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1566), .B(n_1572), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1566), .B(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1567), .B(n_1576), .Y(n_1575) );
OR2x2_ASAP7_75t_L g1631 ( .A(n_1567), .B(n_1573), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1567), .B(n_1640), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1567), .B(n_1573), .Y(n_1702) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1568), .B(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1568), .B(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1602 ( .A(n_1569), .B(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1572), .B(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1572), .Y(n_1697) );
OAI211xp5_ASAP7_75t_L g1705 ( .A1(n_1572), .A2(n_1706), .B(n_1708), .C(n_1709), .Y(n_1705) );
NAND3xp33_ASAP7_75t_L g1718 ( .A(n_1572), .B(n_1605), .C(n_1615), .Y(n_1718) );
AOI221xp5_ASAP7_75t_L g1574 ( .A1(n_1575), .A2(n_1577), .B1(n_1579), .B2(n_1582), .C(n_1584), .Y(n_1574) );
NAND2x1_ASAP7_75t_L g1645 ( .A(n_1575), .B(n_1620), .Y(n_1645) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1576), .Y(n_1581) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
OR2x2_ASAP7_75t_L g1650 ( .A(n_1578), .B(n_1651), .Y(n_1650) );
OAI21xp33_ASAP7_75t_L g1678 ( .A1(n_1579), .A2(n_1649), .B(n_1679), .Y(n_1678) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
NOR2x1_ASAP7_75t_L g1619 ( .A(n_1581), .B(n_1620), .Y(n_1619) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1586), .Y(n_1668) );
OAI321xp33_ASAP7_75t_L g1699 ( .A1(n_1586), .A2(n_1685), .A3(n_1700), .B1(n_1701), .B2(n_1704), .C(n_1705), .Y(n_1699) );
OAI221xp5_ASAP7_75t_L g1711 ( .A1(n_1586), .A2(n_1712), .B1(n_1719), .B2(n_1722), .C(n_1724), .Y(n_1711) );
INVx2_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1588), .B(n_1605), .Y(n_1604) );
NOR2xp33_ASAP7_75t_SL g1708 ( .A(n_1588), .B(n_1607), .Y(n_1708) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
OAI221xp5_ASAP7_75t_L g1589 ( .A1(n_1590), .A2(n_1591), .B1(n_1592), .B2(n_1593), .C(n_1594), .Y(n_1589) );
CKINVDCx20_ASAP7_75t_R g1732 ( .A(n_1592), .Y(n_1732) );
INVxp67_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1601), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1598), .B(n_1618), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1598), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
OR2x2_ASAP7_75t_L g1638 ( .A(n_1599), .B(n_1606), .Y(n_1638) );
NOR3xp33_ASAP7_75t_L g1676 ( .A(n_1599), .B(n_1662), .C(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
AOI221xp5_ASAP7_75t_L g1691 ( .A1(n_1602), .A2(n_1637), .B1(n_1689), .B2(n_1692), .C(n_1694), .Y(n_1691) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1603), .Y(n_1690) );
AOI31xp33_ASAP7_75t_L g1694 ( .A1(n_1605), .A2(n_1684), .A3(n_1695), .B(n_1698), .Y(n_1694) );
NOR2xp33_ASAP7_75t_L g1721 ( .A(n_1605), .B(n_1616), .Y(n_1721) );
CKINVDCx14_ASAP7_75t_R g1605 ( .A(n_1606), .Y(n_1605) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1606), .B(n_1628), .Y(n_1642) );
OR2x2_ASAP7_75t_L g1659 ( .A(n_1606), .B(n_1656), .Y(n_1659) );
OAI21xp5_ASAP7_75t_L g1701 ( .A1(n_1606), .A2(n_1702), .B(n_1703), .Y(n_1701) );
INVx3_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1607), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1607), .B(n_1688), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1612), .Y(n_1627) );
OAI211xp5_ASAP7_75t_L g1613 ( .A1(n_1614), .A2(n_1616), .B(n_1617), .C(n_1621), .Y(n_1613) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1616), .Y(n_1635) );
O2A1O1Ixp33_ASAP7_75t_SL g1725 ( .A1(n_1616), .A2(n_1726), .B(n_1727), .C(n_1730), .Y(n_1725) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1619), .Y(n_1658) );
O2A1O1Ixp33_ASAP7_75t_L g1712 ( .A1(n_1619), .A2(n_1637), .B(n_1713), .C(n_1715), .Y(n_1712) );
CKINVDCx5p33_ASAP7_75t_R g1674 ( .A(n_1620), .Y(n_1674) );
NOR2xp33_ASAP7_75t_L g1679 ( .A(n_1620), .B(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1623), .B(n_1667), .Y(n_1716) );
A2O1A1Ixp33_ASAP7_75t_L g1624 ( .A1(n_1625), .A2(n_1627), .B(n_1628), .C(n_1629), .Y(n_1624) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
OAI211xp5_ASAP7_75t_SL g1633 ( .A1(n_1628), .A2(n_1634), .B(n_1636), .C(n_1647), .Y(n_1633) );
CKINVDCx5p33_ASAP7_75t_R g1698 ( .A(n_1628), .Y(n_1698) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_1630), .B(n_1646), .Y(n_1717) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1631), .Y(n_1703) );
NOR5xp2_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1652), .C(n_1657), .D(n_1661), .E(n_1664), .Y(n_1632) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1643), .Y(n_1700) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1646), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1648), .B(n_1649), .Y(n_1647) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1654), .Y(n_1704) );
CKINVDCx5p33_ASAP7_75t_R g1655 ( .A(n_1656), .Y(n_1655) );
OAI21xp33_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1659), .B(n_1660), .Y(n_1657) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1663), .Y(n_1684) );
NOR2xp33_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1667), .Y(n_1664) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
NOR4xp25_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1681), .C(n_1691), .D(n_1699), .Y(n_1669) );
OAI211xp5_ASAP7_75t_SL g1670 ( .A1(n_1671), .A2(n_1672), .B(n_1675), .C(n_1678), .Y(n_1670) );
INVxp67_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
INVxp67_ASAP7_75t_SL g1675 ( .A(n_1676), .Y(n_1675) );
OAI211xp5_ASAP7_75t_L g1715 ( .A1(n_1686), .A2(n_1716), .B(n_1717), .C(n_1718), .Y(n_1715) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1708), .Y(n_1726) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
INVxp67_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
CKINVDCx20_ASAP7_75t_R g1731 ( .A(n_1732), .Y(n_1731) );
HB1xp67_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
AND4x1_ASAP7_75t_L g1735 ( .A(n_1736), .B(n_1771), .C(n_1796), .D(n_1813), .Y(n_1735) );
OAI21xp33_ASAP7_75t_L g1736 ( .A1(n_1737), .A2(n_1756), .B(n_1769), .Y(n_1736) );
INVx2_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
AOI22xp33_ASAP7_75t_L g1741 ( .A1(n_1742), .A2(n_1743), .B1(n_1745), .B2(n_1746), .Y(n_1741) );
AOI22xp33_ASAP7_75t_L g1813 ( .A1(n_1742), .A2(n_1745), .B1(n_1814), .B2(n_1817), .Y(n_1813) );
BUFx6f_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
AOI21xp5_ASAP7_75t_L g1747 ( .A1(n_1748), .A2(n_1752), .B(n_1754), .Y(n_1747) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1755), .Y(n_1764) );
INVx2_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
INVx4_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
INVx2_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx2_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
NOR2x1_ASAP7_75t_L g1762 ( .A(n_1763), .B(n_1764), .Y(n_1762) );
HB1xp67_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
NOR3xp33_ASAP7_75t_L g1771 ( .A(n_1772), .B(n_1777), .C(n_1789), .Y(n_1771) );
AND2x4_ASAP7_75t_SL g1793 ( .A(n_1773), .B(n_1794), .Y(n_1793) );
AND2x4_ASAP7_75t_L g1773 ( .A(n_1774), .B(n_1775), .Y(n_1773) );
OR2x2_ASAP7_75t_L g1802 ( .A(n_1774), .B(n_1803), .Y(n_1802) );
OAI21xp5_ASAP7_75t_L g1778 ( .A1(n_1779), .A2(n_1780), .B(n_1781), .Y(n_1778) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1793), .Y(n_1792) );
INVx2_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
AOI21xp5_ASAP7_75t_L g1796 ( .A1(n_1797), .A2(n_1804), .B(n_1805), .Y(n_1796) );
INVx8_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
AND2x4_ASAP7_75t_L g1798 ( .A(n_1799), .B(n_1802), .Y(n_1798) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1800), .Y(n_1816) );
AND2x4_ASAP7_75t_L g1806 ( .A(n_1807), .B(n_1808), .Y(n_1806) );
OR2x6_ASAP7_75t_L g1810 ( .A(n_1811), .B(n_1812), .Y(n_1810) );
AND2x4_ASAP7_75t_L g1814 ( .A(n_1815), .B(n_1816), .Y(n_1814) );
CKINVDCx5p33_ASAP7_75t_R g1818 ( .A(n_1819), .Y(n_1818) );
HB1xp67_ASAP7_75t_SL g1822 ( .A(n_1823), .Y(n_1822) );
BUFx3_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVxp33_ASAP7_75t_SL g1825 ( .A(n_1826), .Y(n_1825) );
HB1xp67_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
NOR4xp25_ASAP7_75t_L g1828 ( .A(n_1829), .B(n_1845), .C(n_1858), .D(n_1867), .Y(n_1828) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
INVx3_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
INVx2_ASAP7_75t_SL g1873 ( .A(n_1874), .Y(n_1873) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1875), .Y(n_1874) );
OAI21xp5_ASAP7_75t_L g1875 ( .A1(n_1876), .A2(n_1877), .B(n_1878), .Y(n_1875) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1879), .Y(n_1878) );
endmodule