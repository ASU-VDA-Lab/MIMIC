module fake_jpeg_13728_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_2),
.B(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_1),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_64),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_4),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_45),
.B1(n_43),
.B2(n_48),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_77),
.B1(n_8),
.B2(n_9),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR4xp25_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_46),
.C(n_51),
.D(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_4),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_46),
.B1(n_53),
.B2(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_64),
.B1(n_48),
.B2(n_44),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_88),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_49),
.B1(n_5),
.B2(n_6),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_12),
.B(n_13),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_17),
.C(n_25),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_18),
.B1(n_32),
.B2(n_31),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_7),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_67),
.B1(n_21),
.B2(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_9),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_24),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_11),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_10),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_109),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_102),
.C(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_11),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_82),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_15),
.C(n_16),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_116),
.B(n_117),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_115),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_87),
.C(n_90),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_26),
.C(n_27),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_107),
.B1(n_95),
.B2(n_108),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_101),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_123),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_113),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_121),
.A3(n_120),
.B1(n_114),
.B2(n_107),
.C1(n_98),
.C2(n_38),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_29),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_114),
.Y(n_129)
);


endmodule