module real_jpeg_5877_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_87),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_1),
.A2(n_100),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_57),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_221),
.B(n_224),
.C(n_227),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_1),
.B(n_235),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_1),
.B(n_52),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_1),
.B(n_34),
.C(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_1),
.B(n_139),
.C(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_1),
.B(n_93),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_2),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_2),
.A2(n_37),
.B1(n_78),
.B2(n_134),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_3),
.A2(n_65),
.B1(n_157),
.B2(n_161),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_5),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_7),
.Y(n_223)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_27),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_9),
.A2(n_27),
.B1(n_144),
.B2(n_149),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_9),
.A2(n_27),
.B1(n_71),
.B2(n_233),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_205),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_204),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_187),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_153),
.C(n_169),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_16),
.B(n_153),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_17),
.B(n_85),
.C(n_117),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_62),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_18),
.A2(n_19),
.B1(n_62),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_18),
.A2(n_19),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_18),
.A2(n_19),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_19),
.B(n_231),
.C(n_269),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_19),
.B(n_290),
.C(n_292),
.Y(n_303)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_29),
.B1(n_51),
.B2(n_53),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_21),
.B(n_52),
.Y(n_182)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_25),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_25),
.Y(n_260)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_26),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_29),
.B(n_51),
.Y(n_309)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_30),
.B(n_54),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_30),
.A2(n_52),
.B1(n_156),
.B2(n_198),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_49),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_52),
.A2(n_156),
.B(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_54),
.B(n_309),
.Y(n_308)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_62),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_74),
.B2(n_81),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_64),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_69),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_69),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_70),
.A2(n_176),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_70),
.A2(n_176),
.B1(n_232),
.B2(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_71),
.Y(n_248)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_75),
.B(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_77),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_77),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_116),
.B1(n_117),
.B2(n_152),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_85),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_85),
.B(n_199),
.C(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_85),
.A2(n_152),
.B1(n_199),
.B2(n_298),
.Y(n_322)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B1(n_112),
.B2(n_115),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_86),
.A2(n_92),
.B1(n_112),
.B2(n_115),
.Y(n_186)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_92),
.A2(n_112),
.B(n_115),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_100),
.Y(n_226)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_116),
.A2(n_117),
.B1(n_181),
.B2(n_258),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_116),
.B(n_258),
.C(n_277),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_116),
.A2(n_117),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_117),
.B(n_186),
.C(n_308),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_132),
.B2(n_143),
.Y(n_117)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_118),
.A2(n_121),
.B1(n_132),
.B2(n_143),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_119),
.A2(n_222),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_121),
.B(n_132),
.Y(n_185)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_128),
.Y(n_280)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_132),
.Y(n_270)
);

AOI22x1_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_164),
.B2(n_168),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_164),
.Y(n_194)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_168),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_165),
.B(n_176),
.Y(n_283)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_183),
.C(n_186),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_181),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_172),
.A2(n_181),
.B1(n_258),
.B2(n_325),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_172),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_181),
.A2(n_258),
.B1(n_259),
.B2(n_263),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_186),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_186),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_186),
.A2(n_214),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_202),
.B2(n_203),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_195),
.B1(n_196),
.B2(n_201),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_199),
.B(n_200),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_199),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_199),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_199),
.Y(n_298)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_236),
.B(n_336),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_208),
.B(n_210),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.C(n_218),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_212),
.B(n_216),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_218),
.B(n_332),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_219),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_220),
.A2(n_230),
.B1(n_231),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_220),
.Y(n_316)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_231),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_253),
.Y(n_254)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_318),
.B(n_333),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_302),
.B(n_317),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_287),
.B(n_301),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_274),
.B(n_286),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_265),
.B(n_273),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_255),
.B(n_264),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_252),
.B(n_254),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_256),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_256),
.B(n_296),
.C(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_263),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_259),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_272),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_283),
.B2(n_284),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_284),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_300),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_300),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_292),
.B1(n_293),
.B2(n_299),
.Y(n_288)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_313),
.C(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_328),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_327),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_326),
.C(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule