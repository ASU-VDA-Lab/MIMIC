module real_jpeg_28874_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_0),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_50),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_2),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_168),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_168),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_2),
.A2(n_50),
.B1(n_52),
.B2(n_168),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_157),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_157),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_3),
.A2(n_50),
.B1(n_52),
.B2(n_157),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_26),
.B1(n_55),
.B2(n_56),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_7),
.A2(n_26),
.B1(n_50),
.B2(n_52),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_8),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_94),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_94),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_8),
.A2(n_50),
.B1(n_52),
.B2(n_94),
.Y(n_238)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_9),
.A2(n_52),
.A3(n_55),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_10),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_11),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_11),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_126),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_12),
.A2(n_50),
.B1(n_52),
.B2(n_126),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_126),
.Y(n_271)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_31),
.B(n_62),
.C(n_65),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_96),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_96),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_15),
.A2(n_50),
.B1(n_52),
.B2(n_96),
.Y(n_182)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_17),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_17),
.A2(n_28),
.B(n_32),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_17),
.B(n_30),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_17),
.A2(n_55),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_17),
.B(n_55),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_17),
.B(n_68),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_17),
.A2(n_84),
.B1(n_88),
.B2(n_250),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_17),
.A2(n_31),
.B(n_267),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_335),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_76),
.B(n_331),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_21),
.B(n_37),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_21),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_25),
.A2(n_34),
.B(n_166),
.C(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_27),
.A2(n_30),
.B1(n_93),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_27),
.A2(n_30),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_27),
.A2(n_30),
.B1(n_125),
.B2(n_197),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_27),
.A2(n_30),
.B(n_35),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_63),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g275 ( 
.A1(n_31),
.A2(n_56),
.A3(n_63),
.B1(n_268),
.B2(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_32),
.B(n_166),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_38),
.A2(n_39),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_40),
.B(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_46),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_46),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_46),
.A2(n_58),
.B1(n_135),
.B2(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_47),
.A2(n_53),
.B1(n_57),
.B2(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_47),
.A2(n_53),
.B1(n_102),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_47),
.A2(n_53),
.B1(n_121),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_47),
.A2(n_53),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_47),
.A2(n_53),
.B1(n_224),
.B2(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_47),
.B(n_166),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_47),
.A2(n_53),
.B1(n_162),
.B2(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_49),
.B(n_50),
.Y(n_228)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_50),
.B(n_255),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_55),
.B(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_58),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_68),
.B1(n_111),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_60),
.A2(n_68),
.B1(n_156),
.B2(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_60),
.A2(n_68),
.B1(n_123),
.B2(n_200),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_65),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_65),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_61),
.A2(n_65),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_61),
.A2(n_65),
.B1(n_158),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_61),
.A2(n_65),
.B1(n_180),
.B2(n_266),
.Y(n_265)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_69),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_75),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_73),
.A2(n_75),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_324),
.B(n_330),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_138),
.A3(n_147),
.B1(n_322),
.B2(n_323),
.C(n_341),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_127),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_79),
.B(n_127),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_108),
.C(n_115),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_80),
.B(n_108),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_97),
.B1(n_98),
.B2(n_107),
.Y(n_80)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_90),
.B2(n_91),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_82),
.A2(n_91),
.B(n_97),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_82),
.A2(n_83),
.B1(n_99),
.B2(n_100),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_86),
.B1(n_89),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_84),
.A2(n_86),
.B1(n_119),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_84),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_84),
.A2(n_86),
.B1(n_244),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_84),
.A2(n_86),
.B1(n_238),
.B2(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_85),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_85),
.A2(n_87),
.B1(n_173),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_85),
.A2(n_174),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g239 ( 
.A(n_87),
.Y(n_239)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_103),
.A2(n_106),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_103),
.A2(n_106),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B(n_114),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_113),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_128),
.CI(n_137),
.CON(n_127),
.SN(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_128),
.C(n_137),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_115),
.A2(n_116),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_124),
.Y(n_116)
);

FAx1_ASAP7_75t_L g305 ( 
.A(n_117),
.B(n_122),
.CI(n_124),
.CON(n_305),
.SN(n_305)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_118),
.B(n_120),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_127),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_136),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_130),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.C(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_130),
.B(n_145),
.C(n_146),
.Y(n_325)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_139),
.B(n_140),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_303),
.A3(n_311),
.B1(n_316),
.B2(n_321),
.C(n_342),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_202),
.C(n_214),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_184),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_150),
.B(n_184),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_169),
.C(n_176),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_151),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_164),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_159),
.B2(n_160),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_160),
.C(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_166),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_169),
.A2(n_176),
.B1(n_177),
.B2(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_169),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_178),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_181),
.B(n_183),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_182),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_191),
.C(n_192),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_189),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_201),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_198),
.C(n_201),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_203),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_204),
.B(n_205),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_207),
.B(n_208),
.C(n_213),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_297),
.B(n_302),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_283),
.B(n_296),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_261),
.B(n_282),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_240),
.B(n_260),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_229),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_219),
.B(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_259),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_242),
.B(n_246),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_252),
.B(n_258),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_251),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_274),
.B1(n_280),
.B2(n_281),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_264)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_273),
.C(n_281),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_271),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_274),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_292),
.C(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_305),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_312),
.A2(n_317),
.B(n_320),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule