module fake_netlist_6_2678_n_34 (n_7, n_6, n_12, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_11, n_8, n_10, n_34);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_34;

wire n_16;
wire n_18;
wire n_21;
wire n_24;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_32;
wire n_22;
wire n_26;
wire n_13;
wire n_28;
wire n_17;
wire n_23;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_31;
wire n_25;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_1),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

AND3x1_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_1),
.C(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_18),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_18),
.B1(n_16),
.B2(n_13),
.Y(n_23)
);

OAI22x1_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_21),
.B1(n_15),
.B2(n_20),
.Y(n_25)
);

OR2x6_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_25),
.Y(n_29)
);

AOI221x1_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_27),
.B1(n_22),
.B2(n_5),
.C(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_20),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_20),
.C(n_4),
.Y(n_33)
);

OAI221xp5_ASAP7_75t_R g34 ( 
.A1(n_33),
.A2(n_32),
.B1(n_6),
.B2(n_11),
.C(n_12),
.Y(n_34)
);


endmodule