module fake_jpeg_1860_n_194 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_194);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_40),
.A2(n_27),
.B1(n_28),
.B2(n_8),
.Y(n_92)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_13),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_57),
.Y(n_100)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_29),
.B(n_4),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_25),
.B(n_6),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_66),
.Y(n_87)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_19),
.B1(n_18),
.B2(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_99),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_14),
.B1(n_34),
.B2(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_37),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_97),
.B1(n_88),
.B2(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_7),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_65),
.B(n_46),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_87),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_98),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_110),
.B1(n_85),
.B2(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_108),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_95),
.B1(n_90),
.B2(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_114),
.Y(n_132)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_115),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_80),
.B(n_93),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_117),
.Y(n_140)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_74),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_74),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_72),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_78),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_144),
.B(n_127),
.C(n_143),
.Y(n_155)
);

OAI22x1_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_85),
.B1(n_101),
.B2(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_108),
.C(n_105),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_150),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_114),
.B(n_118),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_157),
.B(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_111),
.C(n_110),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_138),
.Y(n_156)
);

NOR4xp25_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_138),
.C(n_136),
.D(n_144),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_117),
.A3(n_103),
.B1(n_104),
.B2(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NAND2x1_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_139),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_165),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_113),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_148),
.C(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.C(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_161),
.Y(n_179)
);

OAI321xp33_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_146),
.A3(n_147),
.B1(n_135),
.B2(n_127),
.C(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_147),
.B1(n_143),
.B2(n_140),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_178),
.B1(n_174),
.B2(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_179),
.C(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_170),
.B(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_159),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_183),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_173),
.B1(n_166),
.B2(n_171),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_107),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_120),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_103),
.B(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

AOI211xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_181),
.B(n_121),
.C(n_122),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_187),
.C(n_190),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_192),
.Y(n_194)
);


endmodule