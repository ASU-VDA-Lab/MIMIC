module fake_jpeg_26503_n_59 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_1),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_3),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_24),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_4),
.C(n_5),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_51),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_50),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_27),
.B1(n_5),
.B2(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_9),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_7),
.B(n_8),
.Y(n_51)
);

OAI211xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_48),
.B(n_36),
.C(n_45),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B(n_36),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_46),
.Y(n_56)
);

AOI332xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_54),
.A3(n_10),
.B1(n_9),
.B2(n_12),
.B3(n_11),
.C1(n_15),
.C2(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_14),
.Y(n_59)
);


endmodule