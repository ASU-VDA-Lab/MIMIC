module fake_jpeg_17793_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_80),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_51),
.B1(n_48),
.B2(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_77),
.B1(n_43),
.B2(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_48),
.B1(n_41),
.B2(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_85),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_47),
.B1(n_54),
.B2(n_52),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_57),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_89),
.B(n_87),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_98),
.Y(n_113)
);

O2A1O1Ixp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_47),
.B(n_23),
.C(n_37),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_22),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_55),
.C(n_53),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_50),
.C(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_115),
.Y(n_122)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_102),
.B(n_103),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_118),
.C(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_116),
.B1(n_111),
.B2(n_114),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_110),
.B1(n_115),
.B2(n_108),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_108),
.B1(n_56),
.B2(n_101),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_121),
.C(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_130),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_3),
.B(n_4),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_131),
.B1(n_5),
.B2(n_6),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.C(n_5),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_4),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_18),
.B(n_32),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_14),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_19),
.B(n_31),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_12),
.B(n_30),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_11),
.B(n_29),
.C(n_26),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_9),
.Y(n_145)
);


endmodule