module fake_jpeg_11438_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_58),
.B(n_46),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_2),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_48),
.B1(n_42),
.B2(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_81),
.B1(n_65),
.B2(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_57),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_56),
.B1(n_52),
.B2(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_94),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_98),
.B1(n_3),
.B2(n_5),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_90),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_20),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_92),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_80),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_96),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_47),
.B1(n_46),
.B2(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_81),
.B1(n_77),
.B2(n_6),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_104),
.B1(n_110),
.B2(n_113),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_31),
.B1(n_35),
.B2(n_41),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_18),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_114),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_22),
.B1(n_39),
.B2(n_36),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_92),
.B1(n_86),
.B2(n_84),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_8),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_11),
.Y(n_120)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_120),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_126),
.B1(n_127),
.B2(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_125),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_15),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_16),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B1(n_111),
.B2(n_124),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_132),
.B1(n_134),
.B2(n_105),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_133),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_132),
.A3(n_110),
.B1(n_103),
.B2(n_119),
.C1(n_108),
.C2(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_119),
.B1(n_110),
.B2(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);


endmodule