module fake_jpeg_6357_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_5),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_5),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_22),
.A2(n_15),
.B1(n_37),
.B2(n_24),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_106)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_23),
.B(n_10),
.CON(n_43),
.SN(n_43)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_30),
.B1(n_37),
.B2(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_45),
.Y(n_64)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_10),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_35),
.Y(n_89)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_31),
.B1(n_27),
.B2(n_10),
.Y(n_111)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_66),
.Y(n_113)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_111),
.B1(n_3),
.B2(n_12),
.Y(n_136)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_78),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_73),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_22),
.B1(n_34),
.B2(n_29),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_77),
.B1(n_86),
.B2(n_107),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_90),
.Y(n_131)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_41),
.B(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_60),
.B1(n_59),
.B2(n_62),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_102),
.B1(n_106),
.B2(n_4),
.Y(n_120)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_21),
.B1(n_35),
.B2(n_18),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_33),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_98),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_95),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_62),
.B1(n_61),
.B2(n_50),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_31),
.B1(n_27),
.B2(n_12),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_50),
.B(n_18),
.Y(n_95)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_103),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_101),
.B(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_42),
.B(n_38),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_49),
.A2(n_36),
.B1(n_32),
.B2(n_17),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_41),
.B(n_11),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_119),
.B1(n_143),
.B2(n_97),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_31),
.B1(n_27),
.B2(n_2),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_81),
.B1(n_74),
.B2(n_94),
.Y(n_159)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_133),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_4),
.B1(n_13),
.B2(n_12),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_63),
.B1(n_108),
.B2(n_92),
.Y(n_157)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_138),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_63),
.B1(n_108),
.B2(n_92),
.Y(n_156)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_79),
.A2(n_14),
.B(n_13),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_74),
.C(n_81),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_153),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_145),
.B(n_149),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_79),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_132),
.C(n_93),
.Y(n_197)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_151),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_98),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_172),
.C(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_90),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_90),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_139),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_84),
.B(n_127),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_162),
.B1(n_177),
.B2(n_125),
.Y(n_187)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_163),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_159),
.A2(n_164),
.B1(n_13),
.B2(n_14),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_91),
.B1(n_87),
.B2(n_80),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_165),
.B1(n_170),
.B2(n_124),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_131),
.B1(n_121),
.B2(n_122),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_70),
.B1(n_64),
.B2(n_104),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_71),
.B1(n_69),
.B2(n_101),
.Y(n_170)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_174),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_109),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_65),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_78),
.B1(n_85),
.B2(n_68),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_182),
.B(n_184),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_199),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_114),
.B(n_117),
.C(n_128),
.D(n_129),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_188),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_93),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_192),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_153),
.A2(n_134),
.B(n_96),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_193),
.A2(n_206),
.B(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_188),
.C(n_190),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_208),
.B1(n_148),
.B2(n_138),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_149),
.B(n_133),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_155),
.A2(n_178),
.B(n_151),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_127),
.B1(n_118),
.B2(n_75),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_146),
.A2(n_169),
.B1(n_170),
.B2(n_158),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_154),
.B1(n_14),
.B2(n_1),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_118),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_220),
.B(n_222),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_174),
.B(n_1),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_171),
.B(n_163),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_234),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_235),
.B1(n_185),
.B2(n_207),
.Y(n_258)
);

BUFx4f_ASAP7_75t_SL g227 ( 
.A(n_201),
.Y(n_227)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_196),
.B(n_182),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_233),
.B(n_185),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_197),
.C(n_199),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_180),
.B(n_204),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_195),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_206),
.B(n_184),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_242),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_212),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_251),
.B(n_255),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_250),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_243),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_244),
.Y(n_261)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx11_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_230),
.C(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_205),
.C(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_217),
.B(n_228),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_256),
.B(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_233),
.B(n_186),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_218),
.B1(n_237),
.B2(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_213),
.B1(n_231),
.B2(n_191),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_253),
.A2(n_237),
.B1(n_221),
.B2(n_213),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_271),
.A2(n_273),
.B1(n_222),
.B2(n_257),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_226),
.B1(n_236),
.B2(n_189),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_256),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_282),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_252),
.B1(n_219),
.B2(n_245),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_276),
.B(n_235),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_278),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_250),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_274),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_271),
.B1(n_260),
.B2(n_239),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_268),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_249),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_245),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_259),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_251),
.C(n_217),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_290),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_259),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_220),
.B1(n_254),
.B2(n_198),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_264),
.B1(n_239),
.B2(n_208),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_235),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_287),
.B(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_270),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_300),
.B(n_248),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_276),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_300),
.B(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_306),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_203),
.B1(n_210),
.B2(n_192),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_308),
.B(n_209),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_311),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_266),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_214),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_304),
.C(n_289),
.Y(n_318)
);

AOI321xp33_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_319),
.A3(n_302),
.B1(n_299),
.B2(n_228),
.C(n_314),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_309),
.B(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_314),
.C(n_315),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_179),
.Y(n_323)
);


endmodule