module fake_jpeg_27550_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_26),
.Y(n_60)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_36),
.B1(n_34),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_45),
.B1(n_38),
.B2(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_36),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_32),
.B1(n_34),
.B2(n_28),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_32),
.B1(n_28),
.B2(n_23),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_87),
.B1(n_89),
.B2(n_63),
.Y(n_99)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

FAx1_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_45),
.CI(n_44),
.CON(n_79),
.SN(n_79)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_21),
.CI(n_37),
.CON(n_104),
.SN(n_104)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_46),
.C(n_11),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_82),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_85),
.B1(n_92),
.B2(n_41),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_44),
.B1(n_46),
.B2(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_96),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_24),
.B1(n_19),
.B2(n_43),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_35),
.B(n_42),
.C(n_19),
.Y(n_90)
);

AOI22x1_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_63),
.B1(n_37),
.B2(n_38),
.Y(n_98)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_42),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_66),
.C(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_99),
.B1(n_35),
.B2(n_39),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_43),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_38),
.B1(n_41),
.B2(n_37),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_53),
.B1(n_66),
.B2(n_64),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_84),
.A3(n_76),
.B1(n_93),
.B2(n_35),
.Y(n_134)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_112),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_21),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_122),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_84),
.B1(n_91),
.B2(n_72),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_43),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_33),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_65),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_35),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_41),
.B1(n_52),
.B2(n_33),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_96),
.B1(n_74),
.B2(n_70),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_90),
.B(n_39),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_39),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_33),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_130),
.A2(n_137),
.B1(n_138),
.B2(n_108),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_100),
.B(n_105),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_94),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_105),
.B1(n_117),
.B2(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_146),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_150),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_120),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_109),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_100),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_119),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_181),
.B1(n_168),
.B2(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_139),
.B(n_144),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_146),
.B1(n_147),
.B2(n_133),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_173),
.B1(n_115),
.B2(n_149),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_103),
.C(n_119),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_135),
.C(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_104),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_126),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_113),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_18),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_126),
.B1(n_108),
.B2(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_182),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_184),
.C(n_191),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_135),
.C(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_190),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_213),
.B1(n_176),
.B2(n_174),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_152),
.C(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_194),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_12),
.C(n_16),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_160),
.C(n_158),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_210),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_202),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_205),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_152),
.B(n_106),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_204),
.B(n_177),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_111),
.B(n_102),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_18),
.B(n_25),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_142),
.B(n_1),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_181),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_167),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_18),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_142),
.C(n_66),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_53),
.Y(n_238)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_218),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_231),
.B1(n_232),
.B2(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_193),
.B(n_182),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_156),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_230),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_238),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_212),
.B1(n_210),
.B2(n_200),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_201),
.B1(n_53),
.B2(n_30),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_0),
.B(n_1),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_0),
.B(n_1),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_191),
.C(n_184),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_246),
.C(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_195),
.C(n_183),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_209),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_202),
.C(n_200),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_201),
.C(n_203),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_260),
.C(n_219),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_29),
.B1(n_64),
.B2(n_25),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

XOR2x2_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_25),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_240),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_64),
.C(n_31),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_25),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_257),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_279),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_222),
.B1(n_220),
.B2(n_230),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_266),
.B(n_268),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_273),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_214),
.B1(n_224),
.B2(n_229),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_215),
.B1(n_217),
.B2(n_225),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_9),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_35),
.C(n_11),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_262),
.C(n_260),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_7),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_280),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_11),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_256),
.B1(n_247),
.B2(n_242),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_3),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_244),
.C(n_280),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_251),
.B(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_279),
.B1(n_264),
.B2(n_2),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_4),
.C(n_14),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_302),
.C(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_4),
.C(n_14),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_303),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_3),
.C(n_4),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_3),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_294),
.C(n_282),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_293),
.C(n_286),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_319),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_307),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_295),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_298),
.Y(n_322)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_299),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_313),
.A2(n_304),
.B1(n_301),
.B2(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_296),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_328),
.C(n_316),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_305),
.C(n_291),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_314),
.B(n_12),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_331),
.B(n_321),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_321),
.A3(n_327),
.B1(n_329),
.B2(n_332),
.C1(n_325),
.C2(n_15),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_2),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_334),
.C2(n_333),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_13),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_338),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_15),
.Y(n_340)
);


endmodule