module fake_jpeg_925_n_77 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_32),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_1),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_23),
.B1(n_32),
.B2(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_33),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_25),
.B1(n_28),
.B2(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_32),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_29),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_44),
.B(n_45),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_31),
.B(n_33),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_46),
.B(n_39),
.Y(n_53)
);

OAI22x1_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_31),
.B(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_37),
.B1(n_32),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_12),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_13),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_54),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_60),
.Y(n_61)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_49),
.B(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_66),
.Y(n_68)
);

FAx1_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_4),
.CI(n_6),
.CON(n_64),
.SN(n_64)
);

NOR3xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_59),
.C(n_7),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_15),
.C(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_69),
.Y(n_71)
);

AO221x1_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_65),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_6),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_61),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_68),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_71),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_63),
.C(n_67),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_11),
.B(n_16),
.Y(n_76)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.C(n_10),
.Y(n_77)
);


endmodule