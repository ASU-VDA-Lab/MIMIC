module fake_jpeg_10795_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_15),
.B(n_50),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_22),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_87),
.Y(n_91)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_88),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_77),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_53),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_59),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_77),
.B1(n_76),
.B2(n_67),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_59),
.B(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_62),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_115),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_32),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_75),
.C(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_61),
.B1(n_69),
.B2(n_68),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_103),
.B1(n_106),
.B2(n_10),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_78),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_120),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_121),
.B(n_7),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_79),
.B1(n_57),
.B2(n_74),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_56),
.B1(n_2),
.B2(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_0),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_70),
.B1(n_66),
.B2(n_60),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_23),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_56),
.A3(n_59),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_135),
.B(n_141),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_136),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_9),
.B1(n_49),
.B2(n_13),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_27),
.B(n_47),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_5),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_26),
.B(n_46),
.C(n_45),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_7),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_29),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_9),
.B(n_10),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_151),
.C(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_12),
.B1(n_18),
.B2(n_20),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_21),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_31),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_156),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_155),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_40),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_151),
.C(n_159),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_153),
.B1(n_150),
.B2(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_166),
.C(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_171),
.Y(n_177)
);


endmodule