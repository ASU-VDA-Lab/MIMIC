module fake_jpeg_29247_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_19),
.Y(n_46)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

OR2x4_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_21),
.B1(n_29),
.B2(n_15),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_49),
.C(n_45),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_68),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_37),
.B(n_39),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_37),
.CI(n_36),
.CON(n_68),
.SN(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_85),
.B1(n_28),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_40),
.B1(n_34),
.B2(n_36),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_78),
.B1(n_20),
.B2(n_23),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_20),
.Y(n_99)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_74),
.B1(n_22),
.B2(n_30),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_27),
.B(n_34),
.C(n_28),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_33),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_21),
.B1(n_29),
.B2(n_33),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_22),
.B1(n_30),
.B2(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_15),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_15),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_93),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_96),
.B1(n_97),
.B2(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_62),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

OR2x4_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_16),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_71),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_70),
.B1(n_85),
.B2(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_9),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_11),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_116),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_126),
.B1(n_97),
.B2(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_125),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_65),
.B1(n_68),
.B2(n_61),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_124),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_63),
.B1(n_82),
.B2(n_77),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_96),
.B1(n_102),
.B2(n_110),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_18),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_18),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_10),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_129),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_73),
.B(n_84),
.C(n_74),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_104),
.B(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_18),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_107),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_112),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_107),
.B1(n_105),
.B2(n_108),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_143),
.B(n_115),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_R g143 ( 
.A1(n_116),
.A2(n_104),
.B(n_4),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_1),
.B(n_5),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_118),
.B(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_113),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_156),
.B(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_120),
.C(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_153),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_144),
.B1(n_131),
.B2(n_13),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_116),
.C(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_12),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_116),
.C(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_128),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_136),
.B1(n_133),
.B2(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_133),
.B1(n_138),
.B2(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_146),
.B(n_151),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_14),
.B(n_6),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_151),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_169),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_1),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_12),
.C(n_13),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_165),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_172),
.A2(n_157),
.B1(n_160),
.B2(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_161),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_176),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_168),
.B(n_170),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_167),
.C(n_169),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_1),
.B(n_8),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

OAI211xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_181),
.B(n_180),
.C(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_8),
.C(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_8),
.Y(n_187)
);


endmodule