module fake_jpeg_29151_n_494 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_33),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_65),
.Y(n_128)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_9),
.C(n_14),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_35),
.C(n_25),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_15),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_68),
.B(n_69),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_16),
.B(n_12),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_77),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_12),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_11),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_23),
.B(n_11),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_92),
.Y(n_150)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_94),
.Y(n_122)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_97),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_48),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_99),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_105),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_31),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_84),
.B1(n_97),
.B2(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_110),
.B1(n_138),
.B2(n_22),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_39),
.B1(n_43),
.B2(n_35),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_53),
.B(n_18),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_41),
.C(n_1),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_64),
.B(n_24),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_119),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_67),
.A2(n_91),
.B1(n_71),
.B2(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_115),
.A2(n_126),
.B1(n_44),
.B2(n_22),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_25),
.B1(n_47),
.B2(n_23),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_31),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_24),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_45),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_29),
.B1(n_30),
.B2(n_21),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_76),
.B(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_148),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_47),
.B1(n_21),
.B2(n_18),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_18),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_122),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_58),
.A2(n_44),
.B1(n_21),
.B2(n_45),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_41),
.B1(n_45),
.B2(n_92),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_46),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_69),
.B(n_48),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_0),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_166),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_94),
.B1(n_96),
.B2(n_62),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_158),
.A2(n_180),
.B1(n_124),
.B2(n_130),
.Y(n_244)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_164),
.Y(n_206)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_162),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_45),
.B1(n_22),
.B2(n_44),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_165),
.A2(n_153),
.B1(n_100),
.B2(n_151),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_45),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_174),
.Y(n_218)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_183),
.B1(n_187),
.B2(n_189),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_115),
.A2(n_89),
.B1(n_82),
.B2(n_10),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_117),
.B1(n_124),
.B2(n_103),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_0),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_204),
.C(n_197),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_105),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_128),
.B(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_186),
.Y(n_236)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_110),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_188)
);

AO22x1_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_204),
.B1(n_180),
.B2(n_193),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_194),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_11),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_10),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_151),
.A2(n_41),
.B1(n_10),
.B2(n_2),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_124),
.Y(n_212)
);

INVx6_ASAP7_75t_SL g200 ( 
.A(n_123),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_SL g202 ( 
.A(n_118),
.B(n_0),
.C(n_1),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_202),
.B(n_203),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_208),
.A2(n_229),
.B1(n_234),
.B2(n_238),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_112),
.A3(n_140),
.B1(n_111),
.B2(n_136),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_204),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_156),
.A2(n_153),
.B1(n_131),
.B2(n_125),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_210),
.A2(n_244),
.B1(n_177),
.B2(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_212),
.B(n_113),
.Y(n_280)
);

NOR2x1p5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_152),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_227),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_123),
.B(n_139),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_231),
.B(n_130),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_130),
.B1(n_131),
.B2(n_125),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_139),
.B(n_122),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_173),
.B(n_140),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_237),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_173),
.B1(n_175),
.B2(n_159),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_175),
.B(n_122),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_179),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_166),
.A2(n_100),
.B1(n_145),
.B2(n_143),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_152),
.B1(n_145),
.B2(n_143),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_262),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_274),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_226),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_159),
.C(n_179),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_251),
.C(n_240),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_199),
.C(n_158),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_261),
.B1(n_279),
.B2(n_229),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_151),
.B1(n_163),
.B2(n_167),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_254),
.A2(n_258),
.A3(n_271),
.B1(n_269),
.B2(n_283),
.Y(n_300)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_188),
.B(n_149),
.C(n_147),
.D(n_137),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_266),
.B(n_206),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_185),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_257),
.Y(n_297)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_236),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_260),
.B(n_277),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_222),
.A2(n_224),
.B1(n_244),
.B2(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_172),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_264),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_181),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_188),
.B(n_201),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_271),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_208),
.A2(n_147),
.B(n_186),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_171),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_273),
.B1(n_271),
.B2(n_216),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_215),
.B(n_188),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_224),
.A2(n_149),
.B1(n_113),
.B2(n_162),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_171),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_205),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_235),
.A2(n_137),
.B(n_160),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_206),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_224),
.A2(n_127),
.B1(n_109),
.B2(n_189),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_212),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_236),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_285),
.A2(n_248),
.B1(n_187),
.B2(n_220),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_259),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_292),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_213),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_245),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_225),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_303),
.C(n_318),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_304),
.A2(n_252),
.B1(n_312),
.B2(n_279),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_308),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_313),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_271),
.A2(n_209),
.B1(n_211),
.B2(n_241),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_262),
.B1(n_249),
.B2(n_255),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_225),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_225),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_216),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_214),
.C(n_220),
.Y(n_318)
);

OAI22x1_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_265),
.B1(n_256),
.B2(n_273),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_320),
.A2(n_325),
.B1(n_314),
.B2(n_213),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_251),
.CI(n_250),
.CON(n_323),
.SN(n_323)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_323),
.B(n_340),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_272),
.B1(n_281),
.B2(n_248),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_298),
.A2(n_254),
.A3(n_276),
.B1(n_280),
.B2(n_256),
.Y(n_329)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_330),
.A2(n_332),
.B1(n_350),
.B2(n_310),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_285),
.A2(n_276),
.B1(n_266),
.B2(n_281),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_331),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_310),
.A2(n_278),
.B1(n_238),
.B2(n_275),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_334),
.A2(n_320),
.B(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_268),
.B1(n_267),
.B2(n_235),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_272),
.B1(n_243),
.B2(n_183),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_286),
.A2(n_232),
.B(n_223),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_341),
.Y(n_356)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_342),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_319),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_343),
.Y(n_359)
);

AND2x2_ASAP7_75t_SL g344 ( 
.A(n_298),
.B(n_216),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_344),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_297),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_347),
.B(n_294),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_223),
.C(n_232),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_302),
.C(n_291),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_286),
.A2(n_243),
.B1(n_157),
.B2(n_226),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_351),
.Y(n_358)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_363),
.A2(n_338),
.B1(n_337),
.B2(n_330),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_313),
.C(n_291),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_366),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_367),
.C(n_369),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_318),
.C(n_305),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_368),
.A2(n_336),
.B1(n_349),
.B2(n_293),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_296),
.C(n_286),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_287),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_345),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_287),
.C(n_284),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_373),
.C(n_376),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_284),
.C(n_290),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_374),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_300),
.C(n_315),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_375),
.B(n_340),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_332),
.B(n_316),
.C(n_314),
.Y(n_376)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_380),
.B1(n_381),
.B2(n_350),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_331),
.A2(n_293),
.B1(n_295),
.B2(n_217),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_327),
.A2(n_293),
.B1(n_295),
.B2(n_217),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_383),
.A2(n_387),
.B1(n_392),
.B2(n_396),
.Y(n_408)
);

AOI222xp33_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_335),
.B1(n_344),
.B2(n_329),
.C1(n_322),
.C2(n_326),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_404),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_363),
.A2(n_344),
.B1(n_351),
.B2(n_334),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_366),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_362),
.A2(n_361),
.B1(n_352),
.B2(n_360),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_395),
.B1(n_398),
.B2(n_407),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_335),
.B1(n_326),
.B2(n_344),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_339),
.B1(n_321),
.B2(n_324),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_367),
.C(n_364),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_373),
.C(n_356),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_379),
.A2(n_324),
.B1(n_321),
.B2(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_399),
.Y(n_411)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_403),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_342),
.Y(n_402)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_354),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_406),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_381),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_389),
.A2(n_372),
.B(n_376),
.Y(n_409)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_415),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_369),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_370),
.B1(n_368),
.B2(n_358),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_416),
.A2(n_418),
.B1(n_421),
.B2(n_423),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_383),
.A2(n_387),
.B1(n_392),
.B2(n_399),
.Y(n_417)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_417),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_398),
.A2(n_395),
.B1(n_386),
.B2(n_390),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_358),
.B1(n_380),
.B2(n_356),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_422),
.B(n_393),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_385),
.A2(n_374),
.B1(n_217),
.B2(n_226),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_384),
.B(n_207),
.C(n_239),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_384),
.C(n_400),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_207),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_168),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_207),
.B(n_239),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_2),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_430),
.C(n_433),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_393),
.C(n_382),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_438),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_391),
.C(n_388),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_410),
.A2(n_396),
.B1(n_403),
.B2(n_182),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_435),
.A2(n_436),
.B1(n_419),
.B2(n_420),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_410),
.A2(n_127),
.B1(n_109),
.B2(n_170),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_114),
.C(n_129),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_442),
.C(n_414),
.Y(n_455)
);

OAI221xp5_ASAP7_75t_L g440 ( 
.A1(n_412),
.A2(n_129),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_440)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_440),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_409),
.C(n_416),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_413),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_427),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_426),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_428),
.A2(n_408),
.B1(n_417),
.B2(n_420),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_450),
.Y(n_462)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_428),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_452),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_437),
.A2(n_418),
.B1(n_423),
.B2(n_421),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_451),
.A2(n_436),
.B1(n_441),
.B2(n_429),
.Y(n_466)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_457),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_434),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_434),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_437),
.B(n_427),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_464),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_408),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_455),
.C(n_450),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_471),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_453),
.A2(n_439),
.B(n_430),
.Y(n_467)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_467),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_441),
.B(n_4),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_470),
.A2(n_4),
.B(n_5),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_4),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_473),
.B(n_480),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_454),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_477),
.Y(n_481)
);

AOI21xp33_ASAP7_75t_L g475 ( 
.A1(n_469),
.A2(n_446),
.B(n_448),
.Y(n_475)
);

O2A1O1Ixp33_ASAP7_75t_SL g482 ( 
.A1(n_475),
.A2(n_478),
.B(n_461),
.C(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_458),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_463),
.A2(n_445),
.B(n_4),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_484),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_462),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_472),
.B(n_462),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_476),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_487),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_465),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_488),
.A2(n_476),
.B(n_483),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_SL g492 ( 
.A(n_491),
.B(n_489),
.C(n_478),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_492),
.A2(n_5),
.B(n_489),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_5),
.Y(n_494)
);


endmodule