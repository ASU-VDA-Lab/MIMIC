module fake_jpeg_7125_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx24_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.C(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_34),
.B1(n_19),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_52),
.B1(n_30),
.B2(n_37),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_15),
.B1(n_22),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_19),
.B1(n_26),
.B2(n_24),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_30),
.B1(n_24),
.B2(n_17),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_27),
.B1(n_35),
.B2(n_25),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_17),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_27),
.B(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_64),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_45),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_36),
.C(n_33),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_67),
.C(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_70),
.B1(n_75),
.B2(n_72),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_18),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_39),
.B1(n_38),
.B2(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_2),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_32),
.B(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_43),
.A3(n_32),
.B1(n_41),
.B2(n_25),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_41),
.B1(n_46),
.B2(n_43),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_85),
.B1(n_90),
.B2(n_93),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_32),
.A3(n_51),
.B1(n_54),
.B2(n_16),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_51),
.B(n_54),
.C(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_42),
.B1(n_16),
.B2(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_103),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_58),
.B1(n_70),
.B2(n_66),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_110),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_68),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_22),
.B(n_95),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_18),
.B(n_68),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_83),
.B(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_18),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_74),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_100),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_93),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_124),
.B(n_127),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_85),
.B(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_97),
.B1(n_104),
.B2(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_79),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_82),
.C(n_81),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_126),
.C(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_81),
.C(n_74),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_95),
.B(n_22),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_5),
.Y(n_141)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_97),
.B1(n_102),
.B2(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_133),
.B1(n_140),
.B2(n_6),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_101),
.B1(n_98),
.B2(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_138),
.C(n_117),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_101),
.C(n_98),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_111),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_118),
.B(n_120),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_103),
.B1(n_22),
.B2(n_7),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_121),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_126),
.B(n_115),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_146),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_117),
.C(n_116),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_153),
.Y(n_160)
);

BUFx12f_ASAP7_75t_SL g146 ( 
.A(n_141),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_13),
.C(n_7),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_13),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_151),
.A2(n_130),
.B1(n_134),
.B2(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_161),
.B1(n_156),
.B2(n_148),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_160),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_165),
.C(n_6),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_159),
.A2(n_146),
.B1(n_145),
.B2(n_149),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_157),
.B1(n_7),
.B2(n_8),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_170),
.B(n_171),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_157),
.C(n_167),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_162),
.B1(n_10),
.B2(n_11),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_163),
.B(n_168),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_177),
.B(n_175),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_8),
.C(n_10),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_11),
.Y(n_180)
);


endmodule