module real_aes_2583_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g526 ( .A(n_0), .B(n_223), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_1), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g157 ( .A(n_2), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_3), .B(n_529), .Y(n_548) );
NAND2xp33_ASAP7_75t_SL g519 ( .A(n_4), .B(n_178), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_5), .B(n_191), .Y(n_214) );
INVx1_ASAP7_75t_L g511 ( .A(n_6), .Y(n_511) );
INVx1_ASAP7_75t_L g248 ( .A(n_7), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_8), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_9), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_10), .Y(n_265) );
AND2x2_ASAP7_75t_L g546 ( .A(n_11), .B(n_147), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_12), .A2(n_793), .B1(n_800), .B2(n_802), .Y(n_799) );
INVx2_ASAP7_75t_L g148 ( .A(n_13), .Y(n_148) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_14), .B(n_113), .C(n_115), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_14), .Y(n_128) );
INVx1_ASAP7_75t_L g224 ( .A(n_15), .Y(n_224) );
AOI221x1_ASAP7_75t_L g514 ( .A1(n_16), .A2(n_180), .B1(n_515), .B2(n_517), .C(n_518), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_17), .B(n_529), .Y(n_582) );
INVx1_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
INVx1_ASAP7_75t_L g221 ( .A(n_19), .Y(n_221) );
INVx1_ASAP7_75t_SL g169 ( .A(n_20), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_21), .B(n_172), .Y(n_194) );
AOI33xp33_ASAP7_75t_L g239 ( .A1(n_22), .A2(n_49), .A3(n_154), .B1(n_165), .B2(n_240), .B3(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_23), .A2(n_517), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_24), .B(n_223), .Y(n_551) );
AOI221xp5_ASAP7_75t_SL g591 ( .A1(n_25), .A2(n_40), .B1(n_517), .B2(n_529), .C(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g258 ( .A(n_26), .Y(n_258) );
OR2x2_ASAP7_75t_L g149 ( .A(n_27), .B(n_91), .Y(n_149) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_27), .A2(n_91), .B(n_148), .Y(n_182) );
INVxp67_ASAP7_75t_L g513 ( .A(n_28), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_29), .B(n_226), .Y(n_586) );
AND2x2_ASAP7_75t_L g540 ( .A(n_30), .B(n_146), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_31), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_32), .A2(n_517), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_33), .B(n_226), .Y(n_593) );
AND2x2_ASAP7_75t_L g159 ( .A(n_34), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g164 ( .A(n_34), .Y(n_164) );
AND2x2_ASAP7_75t_L g178 ( .A(n_34), .B(n_157), .Y(n_178) );
INVxp67_ASAP7_75t_L g115 ( .A(n_35), .Y(n_115) );
OR2x6_ASAP7_75t_L g130 ( .A(n_35), .B(n_109), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_36), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_37), .B(n_152), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_38), .A2(n_181), .B1(n_187), .B2(n_191), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_39), .B(n_196), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_41), .A2(n_83), .B1(n_162), .B2(n_517), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_42), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_43), .B(n_223), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_44), .B(n_198), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_45), .B(n_172), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_46), .Y(n_190) );
AND2x2_ASAP7_75t_L g530 ( .A(n_47), .B(n_146), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_48), .B(n_146), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_50), .B(n_172), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_51), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_51), .A2(n_63), .B1(n_437), .B2(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g155 ( .A(n_52), .Y(n_155) );
INVx1_ASAP7_75t_L g174 ( .A(n_52), .Y(n_174) );
AOI22x1_ASAP7_75t_L g793 ( .A1(n_53), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_53), .Y(n_794) );
AND2x2_ASAP7_75t_L g290 ( .A(n_54), .B(n_146), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_55), .A2(n_76), .B1(n_152), .B2(n_162), .C(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_56), .B(n_152), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_57), .B(n_529), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_58), .A2(n_805), .B(n_820), .Y(n_804) );
INVx1_ASAP7_75t_L g823 ( .A(n_58), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_59), .B(n_181), .Y(n_267) );
AOI21xp5_ASAP7_75t_SL g203 ( .A1(n_60), .A2(n_162), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g567 ( .A(n_61), .B(n_146), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_62), .B(n_226), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_63), .Y(n_818) );
INVx1_ASAP7_75t_L g217 ( .A(n_64), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_65), .B(n_223), .Y(n_565) );
AND2x2_ASAP7_75t_SL g587 ( .A(n_66), .B(n_147), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_67), .A2(n_517), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g288 ( .A(n_68), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_69), .B(n_226), .Y(n_552) );
AND2x2_ASAP7_75t_SL g559 ( .A(n_70), .B(n_198), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_71), .A2(n_103), .B1(n_797), .B2(n_798), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_71), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_72), .A2(n_162), .B(n_287), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_73), .A2(n_816), .B1(n_817), .B2(n_819), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_73), .Y(n_816) );
INVx1_ASAP7_75t_L g160 ( .A(n_74), .Y(n_160) );
INVx1_ASAP7_75t_L g176 ( .A(n_74), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_75), .B(n_152), .Y(n_242) );
AND2x2_ASAP7_75t_L g179 ( .A(n_77), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g218 ( .A(n_78), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_79), .A2(n_162), .B(n_168), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_80), .A2(n_162), .B(n_193), .C(n_197), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_81), .A2(n_86), .B1(n_152), .B2(n_529), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_82), .B(n_529), .Y(n_566) );
INVx1_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_85), .B(n_180), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_87), .A2(n_162), .B1(n_237), .B2(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_88), .B(n_223), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_89), .B(n_223), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_90), .A2(n_517), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g205 ( .A(n_92), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_93), .B(n_226), .Y(n_564) );
AND2x2_ASAP7_75t_L g243 ( .A(n_94), .B(n_180), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_95), .A2(n_256), .B(n_257), .C(n_259), .Y(n_255) );
INVxp67_ASAP7_75t_L g516 ( .A(n_96), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_97), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_98), .B(n_226), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_99), .A2(n_517), .B(n_584), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_100), .Y(n_125) );
BUFx2_ASAP7_75t_L g121 ( .A(n_101), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_102), .B(n_172), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_103), .Y(n_798) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_116), .B(n_827), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_107), .B(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_112), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OA22x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_131), .B1(n_804), .B2(n_825), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
CKINVDCx11_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g826 ( .A(n_119), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_124), .A2(n_821), .B(n_822), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g824 ( .A(n_126), .Y(n_824) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g808 ( .A(n_127), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x6_ASAP7_75t_SL g501 ( .A(n_128), .B(n_130), .Y(n_501) );
OR2x6_ASAP7_75t_SL g792 ( .A(n_128), .B(n_129), .Y(n_792) );
OR2x2_ASAP7_75t_L g803 ( .A(n_128), .B(n_130), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_793), .B(n_799), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_500), .B1(n_502), .B2(n_790), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_135), .A2(n_500), .B1(n_503), .B2(n_801), .Y(n_800) );
AND3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_494), .C(n_497), .Y(n_135) );
NAND5xp2_ASAP7_75t_L g136 ( .A(n_137), .B(n_394), .C(n_424), .D(n_438), .E(n_464), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_138), .A2(n_437), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g812 ( .A(n_138), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_343), .Y(n_138) );
NOR3xp33_ASAP7_75t_SL g139 ( .A(n_140), .B(n_291), .C(n_325), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_208), .B(n_230), .C(n_269), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_183), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_143), .B(n_281), .Y(n_346) );
AND2x2_ASAP7_75t_L g433 ( .A(n_143), .B(n_211), .Y(n_433) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OR2x2_ASAP7_75t_L g229 ( .A(n_144), .B(n_200), .Y(n_229) );
INVx1_ASAP7_75t_L g271 ( .A(n_144), .Y(n_271) );
INVx2_ASAP7_75t_L g276 ( .A(n_144), .Y(n_276) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_144), .Y(n_304) );
INVx1_ASAP7_75t_L g318 ( .A(n_144), .Y(n_318) );
AND2x2_ASAP7_75t_L g322 ( .A(n_144), .B(n_213), .Y(n_322) );
AND2x2_ASAP7_75t_L g403 ( .A(n_144), .B(n_212), .Y(n_403) );
AO21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_150), .B(n_179), .Y(n_144) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_145), .A2(n_534), .B(n_540), .Y(n_533) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_145), .A2(n_561), .B(n_567), .Y(n_560) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_145), .A2(n_534), .B(n_540), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_146), .Y(n_145) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_146), .A2(n_591), .B(n_595), .Y(n_590) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x4_ASAP7_75t_L g191 ( .A(n_148), .B(n_149), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_161), .Y(n_150) );
INVx1_ASAP7_75t_L g268 ( .A(n_152), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_152), .A2(n_162), .B1(n_510), .B2(n_512), .Y(n_509) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_158), .Y(n_152) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
OR2x6_ASAP7_75t_L g170 ( .A(n_154), .B(n_166), .Y(n_170) );
INVxp33_ASAP7_75t_L g240 ( .A(n_154), .Y(n_240) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g167 ( .A(n_155), .B(n_157), .Y(n_167) );
AND2x4_ASAP7_75t_L g226 ( .A(n_155), .B(n_175), .Y(n_226) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x6_ASAP7_75t_L g517 ( .A(n_159), .B(n_167), .Y(n_517) );
INVx2_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
AND2x6_ASAP7_75t_L g223 ( .A(n_160), .B(n_173), .Y(n_223) );
INVxp67_ASAP7_75t_L g266 ( .A(n_162), .Y(n_266) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_167), .Y(n_162) );
NOR2x1p5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx1_ASAP7_75t_L g241 ( .A(n_165), .Y(n_241) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_177), .Y(n_168) );
INVx2_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_177), .B(n_205), .C(n_206), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_170), .A2(n_217), .B1(n_218), .B2(n_219), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_170), .A2(n_177), .B(n_248), .C(n_249), .Y(n_247) );
INVxp67_ASAP7_75t_L g256 ( .A(n_170), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_170), .A2(n_177), .B(n_288), .C(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
AND2x4_ASAP7_75t_L g529 ( .A(n_172), .B(n_178), .Y(n_529) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_177), .A2(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_177), .B(n_191), .Y(n_227) );
INVx1_ASAP7_75t_L g237 ( .A(n_177), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_177), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_177), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_177), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_177), .A2(n_564), .B(n_565), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_177), .A2(n_585), .B(n_586), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_177), .A2(n_593), .B(n_594), .Y(n_592) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_178), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_180), .A2(n_255), .B1(n_260), .B2(n_261), .Y(n_254) );
INVx3_ASAP7_75t_L g261 ( .A(n_180), .Y(n_261) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_181), .B(n_264), .Y(n_263) );
AOI21x1_ASAP7_75t_L g522 ( .A1(n_181), .A2(n_523), .B(n_530), .Y(n_522) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx4f_ASAP7_75t_L g198 ( .A(n_182), .Y(n_198) );
AND2x4_ASAP7_75t_SL g183 ( .A(n_184), .B(n_199), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
AND2x2_ASAP7_75t_L g272 ( .A(n_185), .B(n_213), .Y(n_272) );
AND2x2_ASAP7_75t_L g293 ( .A(n_185), .B(n_200), .Y(n_293) );
INVx1_ASAP7_75t_L g316 ( .A(n_185), .Y(n_316) );
AND2x4_ASAP7_75t_L g383 ( .A(n_185), .B(n_212), .Y(n_383) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_192), .Y(n_185) );
NOR3xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .C(n_190), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_191), .A2(n_203), .B(n_207), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_191), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_191), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_191), .B(n_516), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_191), .B(n_219), .C(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_191), .A2(n_548), .B(n_549), .Y(n_547) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_197), .A2(n_235), .B(n_243), .Y(n_234) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_197), .A2(n_235), .B(n_243), .Y(n_298) );
AOI21x1_ASAP7_75t_L g555 ( .A1(n_197), .A2(n_556), .B(n_559), .Y(n_555) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_198), .A2(n_246), .B(n_250), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_198), .A2(n_582), .B(n_583), .Y(n_581) );
AND2x4_ASAP7_75t_L g399 ( .A(n_199), .B(n_316), .Y(n_399) );
OR2x2_ASAP7_75t_L g440 ( .A(n_199), .B(n_441), .Y(n_440) );
NOR2xp67_ASAP7_75t_SL g459 ( .A(n_199), .B(n_332), .Y(n_459) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_199), .B(n_391), .Y(n_477) );
INVx4_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2x1_ASAP7_75t_SL g277 ( .A(n_200), .B(n_213), .Y(n_277) );
AND2x4_ASAP7_75t_L g315 ( .A(n_200), .B(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_200), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_200), .B(n_275), .Y(n_353) );
INVx2_ASAP7_75t_L g367 ( .A(n_200), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_200), .B(n_319), .Y(n_389) );
AND2x2_ASAP7_75t_L g481 ( .A(n_200), .B(n_339), .Y(n_481) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2x1_ASAP7_75t_L g209 ( .A(n_210), .B(n_229), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_211), .B(n_318), .Y(n_332) );
AND2x2_ASAP7_75t_SL g341 ( .A(n_211), .B(n_321), .Y(n_341) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_228), .Y(n_211) );
INVx1_ASAP7_75t_L g319 ( .A(n_212), .Y(n_319) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g339 ( .A(n_213), .Y(n_339) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B(n_227), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_219), .B(n_258), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B1(n_224), .B2(n_225), .Y(n_220) );
INVxp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g372 ( .A(n_228), .Y(n_372) );
INVx2_ASAP7_75t_SL g417 ( .A(n_229), .Y(n_417) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_251), .Y(n_231) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_232), .B(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g363 ( .A(n_232), .Y(n_363) );
AND2x2_ASAP7_75t_L g487 ( .A(n_232), .B(n_312), .Y(n_487) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_244), .Y(n_232) );
AND2x4_ASAP7_75t_L g300 ( .A(n_233), .B(n_282), .Y(n_300) );
INVx1_ASAP7_75t_L g311 ( .A(n_233), .Y(n_311) );
AND2x2_ASAP7_75t_L g342 ( .A(n_233), .B(n_297), .Y(n_342) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_234), .B(n_245), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_234), .B(n_283), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_236), .B(n_242), .Y(n_235) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g280 ( .A(n_245), .Y(n_280) );
AND2x4_ASAP7_75t_L g348 ( .A(n_245), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g360 ( .A(n_245), .Y(n_360) );
INVx1_ASAP7_75t_L g402 ( .A(n_245), .Y(n_402) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_245), .Y(n_414) );
AND2x2_ASAP7_75t_L g430 ( .A(n_245), .B(n_253), .Y(n_430) );
BUFx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g377 ( .A(n_252), .B(n_335), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_252), .Y(n_379) );
AND2x2_ASAP7_75t_L g400 ( .A(n_252), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g279 ( .A(n_253), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g307 ( .A(n_253), .Y(n_307) );
INVx2_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_253), .B(n_283), .Y(n_328) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_262), .Y(n_253) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_261), .A2(n_284), .B(n_290), .Y(n_283) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_261), .A2(n_284), .B(n_290), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B1(n_267), .B2(n_268), .Y(n_262) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_273), .B(n_278), .Y(n_269) );
INVx1_ASAP7_75t_L g409 ( .A(n_270), .Y(n_409) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g329 ( .A(n_272), .Y(n_329) );
AND2x2_ASAP7_75t_L g385 ( .A(n_272), .B(n_321), .Y(n_385) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_274), .B(n_315), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_274), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g406 ( .A(n_274), .B(n_399), .Y(n_406) );
AND2x2_ASAP7_75t_L g480 ( .A(n_274), .B(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_275), .Y(n_468) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_276), .Y(n_388) );
AND2x2_ASAP7_75t_L g301 ( .A(n_277), .B(n_302), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_277), .A2(n_490), .B(n_492), .Y(n_489) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx3_ASAP7_75t_L g375 ( .A(n_279), .Y(n_375) );
NAND2x1_ASAP7_75t_SL g419 ( .A(n_279), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g422 ( .A(n_279), .B(n_300), .Y(n_422) );
AND2x2_ASAP7_75t_L g334 ( .A(n_281), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g471 ( .A(n_281), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g482 ( .A(n_281), .B(n_430), .Y(n_482) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_282), .B(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g413 ( .A(n_283), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
OAI21xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_305), .B(n_308), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B1(n_300), .B2(n_301), .Y(n_292) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_299), .Y(n_294) );
AND2x2_ASAP7_75t_L g323 ( .A(n_295), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g429 ( .A(n_295), .B(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_295), .A2(n_448), .B1(n_449), .B2(n_450), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_295), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_297), .B(n_313), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_297), .B(n_313), .Y(n_393) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_297), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g349 ( .A(n_298), .Y(n_349) );
AND2x2_ASAP7_75t_L g357 ( .A(n_298), .B(n_313), .Y(n_357) );
INVx1_ASAP7_75t_L g420 ( .A(n_298), .Y(n_420) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2x1_ASAP7_75t_L g338 ( .A(n_303), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g450 ( .A(n_306), .B(n_335), .Y(n_450) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g324 ( .A(n_307), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_307), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g435 ( .A(n_307), .B(n_342), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_314), .B1(n_320), .B2(n_323), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g443 ( .A(n_310), .B(n_444), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g473 ( .A(n_313), .B(n_360), .Y(n_473) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_L g340 ( .A(n_315), .Y(n_340) );
OAI21xp33_ASAP7_75t_SL g486 ( .A1(n_315), .A2(n_487), .B(n_488), .Y(n_486) );
AND2x4_ASAP7_75t_SL g317 ( .A(n_318), .B(n_319), .Y(n_317) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_318), .Y(n_476) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_SL g418 ( .A1(n_321), .A2(n_419), .B(n_421), .C(n_423), .Y(n_418) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_322), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g423 ( .A(n_322), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_322), .B(n_399), .Y(n_463) );
INVx1_ASAP7_75t_SL g330 ( .A(n_323), .Y(n_330) );
AND2x2_ASAP7_75t_L g411 ( .A(n_324), .B(n_348), .Y(n_411) );
INVx1_ASAP7_75t_L g456 ( .A(n_324), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_330), .B2(n_331), .C(n_333), .Y(n_325) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_326), .Y(n_445) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g493 ( .A(n_328), .B(n_336), .Y(n_493) );
OR2x2_ASAP7_75t_L g352 ( .A(n_329), .B(n_353), .Y(n_352) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_329), .B(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_329), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g491 ( .A(n_329), .B(n_388), .Y(n_491) );
BUFx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI32xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_337), .A3(n_340), .B1(n_341), .B2(n_342), .Y(n_333) );
INVx1_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_337), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g449 ( .A(n_338), .Y(n_449) );
OAI22xp33_ASAP7_75t_SL g431 ( .A1(n_340), .A2(n_432), .B1(n_434), .B2(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g462 ( .A(n_341), .Y(n_462) );
AOI211x1_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_350), .B(n_351), .C(n_368), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_345), .B(n_430), .Y(n_436) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g392 ( .A(n_348), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g458 ( .A(n_348), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B1(n_355), .B2(n_361), .C1(n_362), .C2(n_364), .Y(n_351) );
INVxp67_ASAP7_75t_L g448 ( .A(n_352), .Y(n_448) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_356), .B(n_441), .Y(n_488) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g404 ( .A(n_357), .B(n_401), .Y(n_404) );
INVx3_ASAP7_75t_L g444 ( .A(n_359), .Y(n_444) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_367), .B(n_383), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B1(n_376), .B2(n_381), .C(n_384), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_370), .A2(n_427), .B(n_429), .Y(n_426) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g380 ( .A(n_374), .Y(n_380) );
OR2x2_ASAP7_75t_L g484 ( .A(n_375), .B(n_420), .Y(n_484) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_378), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_381), .A2(n_410), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_382), .A2(n_454), .B(n_461), .Y(n_460) );
INVx4_ASAP7_75t_L g391 ( .A(n_383), .Y(n_391) );
OAI31xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_386), .A3(n_390), .B(n_392), .Y(n_384) );
INVx1_ASAP7_75t_L g442 ( .A(n_386), .Y(n_442) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_407), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_395), .B(n_407), .C(n_426), .D(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_405), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B1(n_403), .B2(n_404), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g467 ( .A(n_399), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_400), .B(n_420), .Y(n_428) );
INVx1_ASAP7_75t_SL g441 ( .A(n_403), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_418), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_412), .B2(n_415), .Y(n_408) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_417), .A2(n_480), .B1(n_482), .B2(n_483), .Y(n_479) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_431), .C(n_437), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g496 ( .A(n_431), .Y(n_496) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_437), .A2(n_498), .B(n_499), .Y(n_497) );
INVxp33_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
AND2x2_ASAP7_75t_L g811 ( .A(n_438), .B(n_464), .Y(n_811) );
NOR2xp67_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_443), .A2(n_466), .B(n_469), .Y(n_465) );
INVx2_ASAP7_75t_L g453 ( .A(n_444), .Y(n_453) );
NAND3xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_451), .C(n_460), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B1(n_457), .B2(n_459), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVxp33_ASAP7_75t_SL g499 ( .A(n_464), .Y(n_499) );
NOR3x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_478), .C(n_485), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_486), .B(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g813 ( .A(n_495), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_667), .Y(n_503) );
NOR4xp25_ASAP7_75t_L g504 ( .A(n_505), .B(n_610), .C(n_649), .D(n_656), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_531), .B1(n_568), .B2(n_577), .C(n_596), .Y(n_505) );
OR2x2_ASAP7_75t_L g740 ( .A(n_506), .B(n_602), .Y(n_740) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g655 ( .A(n_507), .B(n_580), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_507), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_507), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
AND2x4_ASAP7_75t_SL g579 ( .A(n_508), .B(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g601 ( .A(n_508), .Y(n_601) );
AND2x2_ASAP7_75t_L g636 ( .A(n_508), .B(n_609), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_508), .B(n_521), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_508), .B(n_603), .Y(n_688) );
OR2x2_ASAP7_75t_L g766 ( .A(n_508), .B(n_580), .Y(n_766) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g588 ( .A(n_521), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_521), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g614 ( .A(n_521), .Y(n_614) );
OR2x2_ASAP7_75t_L g619 ( .A(n_521), .B(n_603), .Y(n_619) );
AND2x2_ASAP7_75t_L g632 ( .A(n_521), .B(n_590), .Y(n_632) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_521), .Y(n_635) );
INVx1_ASAP7_75t_L g647 ( .A(n_521), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_521), .B(n_601), .Y(n_712) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_541), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g576 ( .A(n_533), .B(n_560), .Y(n_576) );
AND2x4_ASAP7_75t_L g606 ( .A(n_533), .B(n_545), .Y(n_606) );
INVx2_ASAP7_75t_L g640 ( .A(n_533), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_533), .B(n_560), .Y(n_698) );
AND2x2_ASAP7_75t_L g745 ( .A(n_533), .B(n_574), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
AOI222xp33_ASAP7_75t_L g733 ( .A1(n_541), .A2(n_605), .B1(n_648), .B2(n_708), .C1(n_734), .C2(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_553), .Y(n_542) );
AND2x2_ASAP7_75t_L g652 ( .A(n_543), .B(n_572), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_543), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g781 ( .A(n_543), .B(n_621), .Y(n_781) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_544), .A2(n_612), .B(n_616), .Y(n_611) );
AND2x2_ASAP7_75t_L g692 ( .A(n_544), .B(n_575), .Y(n_692) );
OR2x2_ASAP7_75t_L g717 ( .A(n_544), .B(n_576), .Y(n_717) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx5_ASAP7_75t_L g571 ( .A(n_545), .Y(n_571) );
AND2x2_ASAP7_75t_L g658 ( .A(n_545), .B(n_640), .Y(n_658) );
AND2x2_ASAP7_75t_L g684 ( .A(n_545), .B(n_560), .Y(n_684) );
OR2x2_ASAP7_75t_L g687 ( .A(n_545), .B(n_574), .Y(n_687) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_545), .Y(n_705) );
AND2x4_ASAP7_75t_SL g762 ( .A(n_545), .B(n_639), .Y(n_762) );
OR2x2_ASAP7_75t_L g771 ( .A(n_545), .B(n_598), .Y(n_771) );
OR2x6_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g604 ( .A(n_553), .Y(n_604) );
AOI221xp5_ASAP7_75t_SL g722 ( .A1(n_553), .A2(n_606), .B1(n_723), .B2(n_725), .C(n_726), .Y(n_722) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_560), .Y(n_553) );
OR2x2_ASAP7_75t_L g661 ( .A(n_554), .B(n_631), .Y(n_661) );
OR2x2_ASAP7_75t_L g671 ( .A(n_554), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g697 ( .A(n_554), .B(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g703 ( .A(n_554), .B(n_622), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_554), .B(n_686), .Y(n_715) );
INVx2_ASAP7_75t_L g728 ( .A(n_554), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_554), .B(n_606), .Y(n_749) );
AND2x2_ASAP7_75t_L g753 ( .A(n_554), .B(n_575), .Y(n_753) );
AND2x2_ASAP7_75t_L g761 ( .A(n_554), .B(n_762), .Y(n_761) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g574 ( .A(n_555), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_560), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g605 ( .A(n_560), .B(n_574), .Y(n_605) );
INVx2_ASAP7_75t_L g622 ( .A(n_560), .Y(n_622) );
AND2x4_ASAP7_75t_L g639 ( .A(n_560), .B(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_560), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g751 ( .A(n_570), .B(n_573), .Y(n_751) );
AND2x4_ASAP7_75t_L g597 ( .A(n_571), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g638 ( .A(n_571), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g665 ( .A(n_571), .B(n_605), .Y(n_665) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g769 ( .A(n_573), .B(n_770), .Y(n_769) );
BUFx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g621 ( .A(n_574), .B(n_622), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_575), .A2(n_642), .B(n_648), .Y(n_641) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_588), .Y(n_578) );
INVx1_ASAP7_75t_SL g695 ( .A(n_579), .Y(n_695) );
AND2x2_ASAP7_75t_L g725 ( .A(n_579), .B(n_635), .Y(n_725) );
AND2x4_ASAP7_75t_L g736 ( .A(n_579), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g602 ( .A(n_580), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g609 ( .A(n_580), .Y(n_609) );
AND2x4_ASAP7_75t_L g615 ( .A(n_580), .B(n_601), .Y(n_615) );
INVx2_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
INVx1_ASAP7_75t_L g675 ( .A(n_580), .Y(n_675) );
OR2x2_ASAP7_75t_L g696 ( .A(n_580), .B(n_680), .Y(n_696) );
OR2x2_ASAP7_75t_L g710 ( .A(n_580), .B(n_590), .Y(n_710) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_580), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_580), .B(n_632), .Y(n_782) );
OR2x6_ASAP7_75t_L g580 ( .A(n_581), .B(n_587), .Y(n_580) );
INVx1_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
AND2x2_ASAP7_75t_L g760 ( .A(n_588), .B(n_626), .Y(n_760) );
AND2x2_ASAP7_75t_L g785 ( .A(n_588), .B(n_615), .Y(n_785) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g603 ( .A(n_590), .Y(n_603) );
BUFx3_ASAP7_75t_L g645 ( .A(n_590), .Y(n_645) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_590), .Y(n_672) );
INVx1_ASAP7_75t_L g681 ( .A(n_590), .Y(n_681) );
AOI33xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .A3(n_604), .B1(n_605), .B2(n_606), .B3(n_607), .Y(n_596) );
AOI21x1_ASAP7_75t_SL g699 ( .A1(n_597), .A2(n_621), .B(n_683), .Y(n_699) );
INVx2_ASAP7_75t_L g729 ( .A(n_597), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_597), .B(n_728), .Y(n_735) );
AND2x2_ASAP7_75t_L g683 ( .A(n_598), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g646 ( .A(n_601), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g747 ( .A(n_602), .Y(n_747) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_603), .Y(n_737) );
OAI32xp33_ASAP7_75t_L g786 ( .A1(n_604), .A2(n_606), .A3(n_782), .B1(n_787), .B2(n_789), .Y(n_786) );
AND2x2_ASAP7_75t_L g704 ( .A(n_605), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g694 ( .A(n_606), .Y(n_694) );
AND2x2_ASAP7_75t_L g759 ( .A(n_606), .B(n_703), .Y(n_759) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_620), .B1(n_623), .B2(n_637), .C(n_641), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_614), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_615), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_615), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_615), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g664 ( .A(n_619), .Y(n_664) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .C(n_633), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_625), .A2(n_687), .B1(n_727), .B2(n_730), .Y(n_726) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g630 ( .A(n_626), .Y(n_630) );
NOR2x1p5_ASAP7_75t_L g644 ( .A(n_626), .B(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_626), .Y(n_666) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI322xp33_ASAP7_75t_L g693 ( .A1(n_629), .A2(n_671), .A3(n_694), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_699), .Y(n_693) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_631), .A2(n_650), .B(n_651), .C(n_653), .Y(n_649) );
OR2x2_ASAP7_75t_L g741 ( .A(n_631), .B(n_695), .Y(n_741) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g648 ( .A(n_632), .B(n_636), .Y(n_648) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g654 ( .A(n_638), .B(n_655), .Y(n_654) );
INVx3_ASAP7_75t_SL g686 ( .A(n_639), .Y(n_686) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_643), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_SL g690 ( .A(n_646), .Y(n_690) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_647), .Y(n_732) );
OR2x6_ASAP7_75t_SL g787 ( .A(n_650), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g777 ( .A1(n_655), .A2(n_778), .B(n_779), .C(n_786), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_659), .B(n_662), .C(n_666), .Y(n_656) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_657), .A2(n_669), .B(n_676), .C(n_700), .Y(n_668) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_713), .C(n_757), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_672), .Y(n_764) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g719 ( .A(n_675), .Y(n_719) );
NOR3xp33_ASAP7_75t_SL g676 ( .A(n_677), .B(n_689), .C(n_693), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_682), .B1(n_685), .B2(n_688), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g721 ( .A(n_681), .Y(n_721) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_681), .Y(n_788) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_SL g774 ( .A(n_687), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
OR2x2_ASAP7_75t_L g724 ( .A(n_690), .B(n_710), .Y(n_724) );
OR2x2_ASAP7_75t_L g775 ( .A(n_690), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g773 ( .A(n_698), .Y(n_773) );
OR2x2_ASAP7_75t_L g789 ( .A(n_698), .B(n_728), .Y(n_789) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B(n_706), .Y(n_700) );
OAI31xp33_ASAP7_75t_L g714 ( .A1(n_701), .A2(n_715), .A3(n_716), .B(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g746 ( .A(n_711), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND4xp25_ASAP7_75t_SL g713 ( .A(n_714), .B(n_722), .C(n_733), .D(n_738), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_721), .Y(n_756) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_742), .B1(n_746), .B2(n_748), .C(n_750), .Y(n_738) );
NAND2xp33_ASAP7_75t_SL g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g783 ( .A(n_742), .Y(n_783) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_743), .B(n_745), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI21xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g778 ( .A(n_752), .Y(n_778) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_758), .B(n_777), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_763), .C(n_767), .Y(n_758) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
AOI21xp33_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_772), .B(n_775), .Y(n_767) );
INVxp33_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_791), .Y(n_801) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_SL g821 ( .A(n_809), .Y(n_821) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .Y(n_809) );
NAND3x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .C(n_813), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g819 ( .A(n_817), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
endmodule