module fake_jpeg_24395_n_90 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_90);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_25),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_48),
.B1(n_21),
.B2(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_25),
.B(n_22),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_42),
.B(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_32),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_22),
.C(n_25),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_51),
.C(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_25),
.B1(n_22),
.B2(n_27),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_52),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_32),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_59),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_60),
.C(n_15),
.Y(n_62)
);

NOR4xp25_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_51),
.C(n_33),
.D(n_44),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_45),
.B(n_20),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_41),
.C(n_33),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_57),
.B(n_33),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_72),
.B(n_20),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_39),
.B1(n_32),
.B2(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_31),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_12),
.A3(n_13),
.B1(n_37),
.B2(n_17),
.C1(n_18),
.C2(n_31),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_13),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_78),
.C(n_28),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_75),
.A2(n_19),
.B1(n_70),
.B2(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.C(n_69),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_37),
.C(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_7),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_4),
.Y(n_88)
);

AOI221xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_3),
.B1(n_4),
.B2(n_10),
.C(n_89),
.Y(n_90)
);


endmodule