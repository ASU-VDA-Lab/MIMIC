module fake_netlist_6_4439_n_1628 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1628);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1628;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g145 ( 
.A(n_33),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_8),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_61),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_10),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_59),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_50),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_28),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_85),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_46),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_17),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_112),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_46),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_67),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_23),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_51),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_48),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_30),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_29),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_6),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_54),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_72),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_53),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_12),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_141),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_6),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_124),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_43),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_137),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_47),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_101),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_83),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_79),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_45),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_18),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_40),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_41),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_82),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_36),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_42),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_4),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_120),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_52),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_18),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_133),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_0),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_144),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_130),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_66),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_123),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_142),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_92),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_106),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_81),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_21),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_17),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_89),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_78),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_107),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_74),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_93),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_33),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_13),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_42),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_29),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_30),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_99),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_11),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_108),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_71),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_139),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_111),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_114),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_129),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_19),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_91),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_96),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_116),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_119),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_90),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_21),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_20),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_11),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_16),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_31),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_103),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_64),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_69),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_73),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_98),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_122),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_55),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_94),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_14),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_80),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_269),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_158),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_182),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_146),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_154),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_184),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_178),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_178),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_158),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_211),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_211),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_166),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_171),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_161),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_156),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_172),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_180),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_186),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_189),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_145),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_161),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_148),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_194),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_181),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_196),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_173),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_168),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_184),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_190),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_186),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_193),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_197),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_201),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_212),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_231),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_199),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_250),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_173),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_149),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_150),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_152),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_184),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_202),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_151),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_175),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_170),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_170),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_225),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_203),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_163),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_204),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_296),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_214),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_214),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_288),
.A2(n_195),
.B1(n_174),
.B2(n_268),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_311),
.A2(n_174),
.B1(n_195),
.B2(n_268),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_324),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_240),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

AND2x2_ASAP7_75t_SL g367 ( 
.A(n_349),
.B(n_225),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_298),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_210),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_284),
.B(n_210),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_312),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_300),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_302),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_285),
.B(n_286),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_302),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_303),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_303),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_304),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_289),
.B(n_343),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_307),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_309),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_290),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_294),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_291),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_314),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_317),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_285),
.B(n_210),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_286),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_353),
.A2(n_261),
.B(n_236),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_305),
.B(n_240),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_354),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_354),
.A2(n_261),
.B(n_236),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_291),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_346),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_346),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_292),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_292),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_320),
.B(n_160),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_351),
.B(n_264),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_301),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_326),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_322),
.B(n_327),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

NOR2x1p5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_163),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_329),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_378),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_264),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_301),
.Y(n_433)
);

BUFx6f_ASAP7_75t_SL g434 ( 
.A(n_367),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_365),
.B(n_306),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_367),
.A2(n_357),
.B1(n_355),
.B2(n_348),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_425),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_367),
.A2(n_368),
.B1(n_376),
.B2(n_405),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_369),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_365),
.B(n_306),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_410),
.B(n_313),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_370),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_368),
.A2(n_376),
.B1(n_385),
.B2(n_313),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_415),
.B(n_315),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_419),
.B(n_315),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_287),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_373),
.A2(n_357),
.B1(n_355),
.B2(n_348),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_153),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_372),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_408),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

AND3x2_ASAP7_75t_L g476 ( 
.A(n_408),
.B(n_283),
.C(n_293),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_377),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_406),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_420),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_372),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_417),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_406),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_359),
.B(n_181),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_L g492 ( 
.A(n_359),
.B(n_181),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_383),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_372),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_423),
.A2(n_283),
.B1(n_335),
.B2(n_341),
.Y(n_497)
);

CKINVDCx6p67_ASAP7_75t_R g498 ( 
.A(n_420),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_381),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_381),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_377),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_381),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_422),
.B(n_323),
.C(n_319),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_422),
.B(n_319),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_393),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_395),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_423),
.A2(n_331),
.B1(n_332),
.B2(n_340),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_395),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_372),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_412),
.B(n_323),
.Y(n_517)
);

NOR2x1p5_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_282),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_384),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_395),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_372),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_360),
.B(n_325),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_375),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_393),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_360),
.B(n_325),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_375),
.Y(n_530)
);

CKINVDCx6p67_ASAP7_75t_R g531 ( 
.A(n_384),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_412),
.A2(n_336),
.B1(n_259),
.B2(n_175),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_397),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_421),
.B(n_336),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_397),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_362),
.A2(n_259),
.B1(n_218),
.B2(n_221),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_407),
.B(n_333),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_375),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_396),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_363),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_426),
.B(n_218),
.Y(n_545)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_423),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_396),
.B(n_162),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_402),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_375),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_402),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_398),
.B(n_328),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_402),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_409),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_363),
.Y(n_555)
);

NOR2x1p5_ASAP7_75t_L g556 ( 
.A(n_418),
.B(n_282),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_399),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_375),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_382),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_402),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_403),
.B(n_347),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_409),
.B(n_334),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_364),
.B(n_147),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_364),
.B(n_157),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_403),
.B(n_337),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_418),
.B(n_235),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_375),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_404),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_404),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_478),
.B(n_366),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_427),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_427),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_520),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_478),
.B(n_366),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_435),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_525),
.B(n_277),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_502),
.B(n_529),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_160),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_502),
.B(n_342),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_517),
.B(n_164),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_520),
.B(n_366),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_428),
.B(n_371),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_433),
.B(n_164),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_428),
.B(n_371),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_449),
.B(n_181),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_441),
.B(n_371),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_441),
.B(n_402),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_442),
.B(n_402),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_432),
.B(n_165),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_546),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_537),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_546),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_458),
.B(n_206),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_539),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_442),
.B(n_413),
.Y(n_596)
);

OAI21xp33_ASAP7_75t_L g597 ( 
.A1(n_552),
.A2(n_338),
.B(n_339),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_436),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_461),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_562),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_445),
.B(n_206),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_455),
.B(n_206),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_444),
.B(n_413),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_498),
.B(n_207),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_444),
.B(n_413),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_450),
.B(n_453),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_519),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_519),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_519),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_500),
.B(n_206),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_473),
.B(n_350),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_463),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_531),
.Y(n_616)
);

BUFx8_ASAP7_75t_L g617 ( 
.A(n_434),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_548),
.Y(n_618)
);

INVx8_ASAP7_75t_L g619 ( 
.A(n_434),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_430),
.B(n_220),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_437),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_548),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_450),
.B(n_413),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_475),
.B(n_213),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_453),
.B(n_413),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_434),
.A2(n_208),
.B1(n_205),
.B2(n_191),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_557),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_509),
.A2(n_234),
.B1(n_188),
.B2(n_187),
.Y(n_628)
);

BUFx5_ASAP7_75t_L g629 ( 
.A(n_432),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_556),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_457),
.B(n_413),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_500),
.B(n_237),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_544),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_447),
.A2(n_215),
.B1(n_209),
.B2(n_200),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_500),
.B(n_506),
.Y(n_636)
);

BUFx5_ASAP7_75t_L g637 ( 
.A(n_432),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_457),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_506),
.B(n_237),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_472),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_472),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_508),
.A2(n_222),
.B1(n_255),
.B2(n_198),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_567),
.B(n_224),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_506),
.B(n_237),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_535),
.B(n_224),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_456),
.B(n_216),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_563),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_474),
.B(n_413),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_569),
.B(n_233),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_437),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_482),
.B(n_382),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_569),
.B(n_241),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_465),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_482),
.B(n_382),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_532),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_546),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_439),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_563),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_531),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_483),
.B(n_382),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_483),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_545),
.A2(n_185),
.B1(n_281),
.B2(n_280),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_566),
.B(n_407),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_485),
.B(n_382),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_485),
.B(n_382),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_487),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_545),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_487),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_493),
.B(n_503),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_546),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_382),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_544),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_503),
.B(n_388),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_505),
.B(n_388),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_510),
.B(n_237),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_547),
.B(n_242),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_566),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_510),
.B(n_253),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_570),
.B(n_411),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_439),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_563),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_440),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_505),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_510),
.B(n_253),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_518),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_521),
.B(n_253),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_518),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_521),
.B(n_467),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_570),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_507),
.B(n_244),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_521),
.B(n_253),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_507),
.B(n_512),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_512),
.B(n_388),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_467),
.B(n_265),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_467),
.B(n_265),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_527),
.B(n_388),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_527),
.B(n_542),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_429),
.A2(n_248),
.B1(n_179),
.B2(n_183),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_542),
.B(n_388),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_494),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_443),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_431),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_494),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_570),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_443),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_446),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_497),
.A2(n_155),
.B1(n_167),
.B2(n_176),
.C(n_177),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_432),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_460),
.B(n_260),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_446),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_554),
.B(n_265),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_538),
.B(n_279),
.C(n_278),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_554),
.B(n_564),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_429),
.A2(n_251),
.B1(n_169),
.B2(n_217),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_499),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_499),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_565),
.B(n_501),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_563),
.A2(n_159),
.B1(n_192),
.B2(n_230),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_501),
.B(n_388),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_504),
.B(n_265),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_504),
.B(n_389),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_498),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_555),
.A2(n_409),
.B1(n_274),
.B2(n_243),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_511),
.B(n_252),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_462),
.B(n_226),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_692),
.B(n_511),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_577),
.A2(n_480),
.B1(n_543),
.B2(n_489),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_L g728 ( 
.A1(n_712),
.A2(n_555),
.B1(n_480),
.B2(n_514),
.C(n_273),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_702),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_577),
.B(n_448),
.C(n_227),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_692),
.B(n_513),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_609),
.B(n_513),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_586),
.A2(n_523),
.B1(n_534),
.B2(n_515),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_638),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_647),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_586),
.A2(n_594),
.B(n_667),
.C(n_635),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_679),
.B(n_219),
.Y(n_737)
);

OR2x4_ASAP7_75t_L g738 ( 
.A(n_709),
.B(n_476),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_656),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_688),
.A2(n_526),
.B(n_438),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_580),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_669),
.B(n_515),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_640),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_697),
.B(n_641),
.Y(n_744)
);

NAND2x1p5_ASAP7_75t_L g745 ( 
.A(n_656),
.B(n_479),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_661),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_R g747 ( 
.A(n_689),
.B(n_228),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_666),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_647),
.B(n_522),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_683),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_614),
.Y(n_752)
);

BUFx4f_ASAP7_75t_L g753 ( 
.A(n_619),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_655),
.A2(n_266),
.B1(n_229),
.B2(n_239),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_620),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_656),
.B(n_670),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_578),
.B(n_254),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_581),
.B(n_522),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_592),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_599),
.Y(n_760)
);

AOI211xp5_ASAP7_75t_L g761 ( 
.A1(n_643),
.A2(n_492),
.B(n_491),
.C(n_257),
.Y(n_761)
);

INVx6_ASAP7_75t_L g762 ( 
.A(n_617),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_599),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_704),
.B(n_256),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_658),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_606),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_700),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_676),
.A2(n_495),
.B1(n_489),
.B2(n_523),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_618),
.B(n_528),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_615),
.B(n_526),
.Y(n_771)
);

NAND2x1p5_ASAP7_75t_L g772 ( 
.A(n_656),
.B(n_495),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_670),
.Y(n_773)
);

AND2x4_ASAP7_75t_SL g774 ( 
.A(n_610),
.B(n_223),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_703),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_670),
.B(n_438),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_601),
.B(n_526),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_223),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_619),
.B(n_528),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_658),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_715),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_595),
.B(n_559),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_716),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_622),
.B(n_534),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_600),
.B(n_624),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_627),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_605),
.B(n_559),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_634),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_688),
.A2(n_438),
.B(n_477),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_630),
.B(n_536),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_723),
.A2(n_536),
.B1(n_454),
.B2(n_459),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_663),
.B(n_466),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_634),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_670),
.B(n_452),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_574),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_583),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_685),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_723),
.A2(n_454),
.B1(n_459),
.B2(n_464),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_585),
.Y(n_799)
);

OR2x2_ASAP7_75t_SL g800 ( 
.A(n_653),
.B(n_223),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_616),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_676),
.B(n_584),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_687),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_636),
.A2(n_477),
.B(n_541),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_617),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_681),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_584),
.B(n_272),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_681),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_591),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_619),
.B(n_466),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_631),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_579),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_646),
.B(n_275),
.Y(n_813)
);

NOR2x1_ASAP7_75t_L g814 ( 
.A(n_607),
.B(n_481),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_672),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_594),
.B(n_491),
.C(n_492),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_649),
.B(n_652),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_659),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_636),
.B(n_451),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_587),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_717),
.B(n_468),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_672),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_649),
.B(n_568),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_725),
.B(n_468),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_652),
.B(n_232),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_680),
.B(n_469),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_680),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_722),
.B(n_276),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_611),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_612),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_705),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_705),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_SL g833 ( 
.A(n_591),
.B(n_452),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_593),
.B(n_477),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_579),
.B(n_232),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_706),
.B(n_469),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_SL g837 ( 
.A1(n_643),
.A2(n_232),
.B1(n_258),
.B2(n_7),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_571),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_593),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_575),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_R g841 ( 
.A(n_709),
.B(n_568),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_613),
.B(n_471),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_626),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_613),
.B(n_471),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_633),
.B(n_484),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_646),
.B(n_524),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_572),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_645),
.B(n_464),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_645),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_690),
.B(n_568),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_628),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_690),
.B(n_530),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_573),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_576),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_713),
.B(n_530),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_602),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_R g857 ( 
.A(n_590),
.B(n_481),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_598),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_708),
.B(n_698),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_714),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_662),
.B(n_496),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_629),
.B(n_452),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_582),
.B(n_561),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_621),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_650),
.B(n_657),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_718),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_682),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_642),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_701),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_629),
.B(n_452),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_629),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_633),
.B(n_561),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_588),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_639),
.B(n_560),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_597),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_602),
.B(n_560),
.C(n_488),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_710),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_603),
.Y(n_878)
);

NOR2x2_ASAP7_75t_L g879 ( 
.A(n_603),
.B(n_258),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_724),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_639),
.B(n_481),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_724),
.B(n_553),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_629),
.B(n_558),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_644),
.B(n_486),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_711),
.A2(n_486),
.B1(n_553),
.B2(n_551),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_651),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_629),
.B(n_558),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_589),
.B(n_484),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_694),
.B(n_488),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_629),
.B(n_558),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_637),
.B(n_558),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_SL g892 ( 
.A(n_694),
.B(n_558),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_644),
.A2(n_551),
.B(n_549),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_637),
.B(n_541),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_654),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_817),
.B(n_675),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_802),
.A2(n_678),
.B(n_675),
.C(n_684),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_752),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_868),
.A2(n_707),
.B1(n_678),
.B2(n_691),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_734),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_840),
.B(n_684),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_SL g902 ( 
.A1(n_800),
.A2(n_812),
.B1(n_849),
.B2(n_805),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_815),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_755),
.B(n_686),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_739),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_871),
.A2(n_794),
.B(n_789),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_755),
.B(n_686),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_815),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_744),
.B(n_691),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_744),
.B(n_596),
.Y(n_910)
);

OR2x6_ASAP7_75t_L g911 ( 
.A(n_762),
.B(n_604),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_871),
.A2(n_695),
.B(n_711),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_726),
.A2(n_695),
.B1(n_608),
.B2(n_623),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_859),
.A2(n_648),
.B1(n_632),
.B2(n_625),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_785),
.B(n_671),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_873),
.A2(n_637),
.B(n_660),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_741),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_838),
.B(n_665),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_796),
.B(n_664),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_799),
.B(n_673),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_727),
.B(n_674),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_825),
.B(n_693),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_866),
.A2(n_720),
.B(n_699),
.C(n_696),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_814),
.B(n_721),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_875),
.A2(n_720),
.B(n_719),
.C(n_549),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_730),
.B(n_637),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_729),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_835),
.B(n_524),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_736),
.A2(n_823),
.B(n_880),
.C(n_851),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_820),
.B(n_637),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_740),
.A2(n_541),
.B(n_524),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_860),
.B(n_541),
.Y(n_932)
);

OR2x6_ASAP7_75t_SL g933 ( 
.A(n_848),
.B(n_1),
.Y(n_933)
);

OA21x2_ASAP7_75t_L g934 ( 
.A1(n_893),
.A2(n_490),
.B(n_541),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_809),
.A2(n_524),
.B(n_550),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_779),
.B(n_56),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_809),
.A2(n_524),
.B(n_550),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_861),
.A2(n_389),
.B(n_516),
.C(n_470),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_801),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_743),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_779),
.B(n_117),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_726),
.A2(n_490),
.B1(n_516),
.B2(n_550),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_728),
.A2(n_389),
.B(n_516),
.C(n_470),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_818),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_809),
.A2(n_550),
.B(n_516),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_746),
.B(n_490),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_809),
.A2(n_550),
.B(n_516),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_748),
.B(n_490),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_829),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_754),
.A2(n_389),
.B1(n_5),
.B2(n_9),
.C(n_10),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_782),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_753),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_843),
.B(n_1),
.Y(n_953)
);

BUFx5_ASAP7_75t_L g954 ( 
.A(n_750),
.Y(n_954)
);

CKINVDCx8_ASAP7_75t_R g955 ( 
.A(n_739),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_759),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_760),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_738),
.B(n_14),
.Y(n_958)
);

CKINVDCx6p67_ASAP7_75t_R g959 ( 
.A(n_779),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_804),
.A2(n_102),
.B(n_143),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_797),
.B(n_97),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_811),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_808),
.Y(n_963)
);

AO32x2_ASAP7_75t_L g964 ( 
.A1(n_798),
.A2(n_15),
.A3(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_964)
);

BUFx5_ASAP7_75t_L g965 ( 
.A(n_750),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_839),
.A2(n_389),
.B(n_135),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_749),
.B(n_15),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_751),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_813),
.A2(n_807),
.B(n_757),
.C(n_737),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_SL g970 ( 
.A1(n_771),
.A2(n_134),
.B(n_121),
.C(n_118),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_808),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_738),
.B(n_22),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_786),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_859),
.A2(n_87),
.B1(n_86),
.B2(n_63),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_830),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_763),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_856),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_SL g978 ( 
.A(n_753),
.B(n_57),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_777),
.B(n_31),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_803),
.B(n_32),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_764),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_773),
.B(n_34),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_792),
.B(n_35),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_778),
.B(n_795),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_767),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_839),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_758),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_987)
);

O2A1O1Ixp5_ASAP7_75t_L g988 ( 
.A1(n_846),
.A2(n_892),
.B(n_852),
.C(n_850),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_770),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_821),
.A2(n_43),
.B(n_44),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_782),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_821),
.A2(n_742),
.B(n_732),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_774),
.B(n_44),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_762),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_788),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_R g996 ( 
.A(n_765),
.B(n_806),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_886),
.B(n_895),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_756),
.B(n_808),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_837),
.B(n_787),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_878),
.B(n_847),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_793),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_731),
.B(n_768),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_881),
.A2(n_816),
.B(n_761),
.C(n_775),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_816),
.A2(n_761),
.B(n_783),
.C(n_781),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_810),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_828),
.B(n_810),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_747),
.B(n_877),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_784),
.A2(n_790),
.B1(n_889),
.B2(n_780),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_735),
.B(n_780),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_735),
.A2(n_766),
.B1(n_806),
.B2(n_889),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_854),
.A2(n_864),
.B(n_867),
.C(n_869),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_841),
.B(n_766),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_862),
.A2(n_894),
.B(n_887),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_853),
.B(n_858),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_870),
.A2(n_891),
.B(n_890),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_853),
.B(n_858),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_827),
.B(n_832),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_SL g1018 ( 
.A(n_769),
.B(n_857),
.C(n_879),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_SL g1019 ( 
.A(n_950),
.B(n_756),
.C(n_865),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_915),
.B(n_888),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_929),
.A2(n_883),
.B(n_884),
.C(n_872),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_906),
.A2(n_893),
.B(n_885),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_992),
.A2(n_834),
.B(n_776),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_896),
.A2(n_876),
.B(n_884),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1002),
.B(n_888),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_904),
.A2(n_745),
.B1(n_772),
.B2(n_810),
.Y(n_1026)
);

BUFx8_ASAP7_75t_SL g1027 ( 
.A(n_927),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1003),
.A2(n_876),
.B(n_842),
.Y(n_1028)
);

AOI221x1_ASAP7_75t_L g1029 ( 
.A1(n_897),
.A2(n_885),
.B1(n_798),
.B2(n_791),
.C(n_833),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_SL g1030 ( 
.A1(n_958),
.A2(n_824),
.B(n_733),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_931),
.A2(n_836),
.B(n_826),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_952),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_938),
.A2(n_791),
.A3(n_855),
.B(n_872),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_SL g1034 ( 
.A1(n_909),
.A2(n_819),
.B(n_874),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1004),
.A2(n_745),
.B(n_772),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_831),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_912),
.A2(n_960),
.B(n_916),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_989),
.B(n_910),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_997),
.B(n_863),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_922),
.A2(n_844),
.B(n_845),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_921),
.B(n_822),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_SL g1042 ( 
.A1(n_972),
.A2(n_844),
.B(n_842),
.Y(n_1042)
);

CKINVDCx11_ASAP7_75t_R g1043 ( 
.A(n_933),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_940),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_917),
.B(n_882),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_SL g1046 ( 
.A1(n_969),
.A2(n_882),
.B(n_990),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_1013),
.A2(n_1015),
.B(n_1010),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_968),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_955),
.Y(n_1049)
);

CKINVDCx11_ASAP7_75t_R g1050 ( 
.A(n_994),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_SL g1051 ( 
.A(n_987),
.B(n_1007),
.C(n_984),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_928),
.A2(n_988),
.B(n_926),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_919),
.B(n_920),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_944),
.B(n_991),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_899),
.A2(n_901),
.B(n_914),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_SL g1056 ( 
.A1(n_902),
.A2(n_979),
.B1(n_977),
.B2(n_973),
.C(n_967),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_991),
.B(n_951),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_975),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_930),
.A2(n_913),
.B(n_1008),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1008),
.A2(n_937),
.B(n_935),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1006),
.B(n_1005),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_918),
.A2(n_923),
.B(n_932),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1018),
.A2(n_983),
.B(n_982),
.C(n_907),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_963),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_943),
.A2(n_942),
.A3(n_1009),
.B(n_974),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_SL g1066 ( 
.A1(n_936),
.A2(n_941),
.B(n_971),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_936),
.B(n_941),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_998),
.A2(n_1012),
.B(n_925),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1006),
.B(n_911),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_998),
.A2(n_1016),
.B(n_1014),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_962),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_970),
.A2(n_993),
.B(n_999),
.C(n_1011),
.Y(n_1072)
);

BUFx8_ASAP7_75t_L g1073 ( 
.A(n_949),
.Y(n_1073)
);

AO32x2_ASAP7_75t_L g1074 ( 
.A1(n_902),
.A2(n_964),
.A3(n_934),
.B1(n_965),
.B2(n_954),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_945),
.A2(n_947),
.B(n_946),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1000),
.B(n_924),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_948),
.A2(n_1017),
.B(n_966),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_963),
.Y(n_1078)
);

OAI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_978),
.A2(n_980),
.B(n_961),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_980),
.Y(n_1080)
);

AO32x2_ASAP7_75t_L g1081 ( 
.A1(n_964),
.A2(n_965),
.A3(n_954),
.B1(n_959),
.B2(n_996),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_963),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_911),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_903),
.A2(n_908),
.A3(n_1001),
.B(n_995),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_956),
.A2(n_976),
.B(n_981),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_957),
.A2(n_985),
.B(n_961),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_971),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_905),
.B(n_965),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_954),
.A2(n_965),
.B(n_964),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_954),
.B(n_965),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_900),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_917),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_900),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_927),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1006),
.B(n_1005),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_L g1099 ( 
.A1(n_979),
.A2(n_817),
.B(n_802),
.C(n_581),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_939),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_969),
.A2(n_817),
.B(n_802),
.C(n_736),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_906),
.A2(n_871),
.B(n_992),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_969),
.A2(n_817),
.B(n_802),
.C(n_736),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_897),
.A2(n_938),
.A3(n_1003),
.B(n_1008),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_897),
.A2(n_988),
.B(n_938),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_953),
.A2(n_817),
.B(n_802),
.C(n_581),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_905),
.Y(n_1107)
);

BUFx2_ASAP7_75t_SL g1108 ( 
.A(n_955),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_SL g1109 ( 
.A(n_986),
.B(n_809),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1110)
);

NAND2x1_ASAP7_75t_L g1111 ( 
.A(n_963),
.B(n_739),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_915),
.B(n_817),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_915),
.B(n_817),
.Y(n_1113)
);

AO32x2_ASAP7_75t_L g1114 ( 
.A1(n_913),
.A2(n_1008),
.A3(n_902),
.B1(n_635),
.B2(n_718),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_898),
.B(n_817),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_929),
.A2(n_817),
.B(n_802),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_915),
.B(n_817),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_900),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_SL g1119 ( 
.A1(n_969),
.A2(n_736),
.B(n_990),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_906),
.A2(n_871),
.B(n_992),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_979),
.A2(n_817),
.B(n_802),
.C(n_581),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_955),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_927),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_898),
.B(n_817),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_900),
.Y(n_1127)
);

NAND4xp25_ASAP7_75t_L g1128 ( 
.A(n_953),
.B(n_362),
.C(n_538),
.D(n_555),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_L g1130 ( 
.A(n_1018),
.B(n_578),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_906),
.A2(n_931),
.B(n_912),
.Y(n_1131)
);

AOI221x1_ASAP7_75t_L g1132 ( 
.A1(n_897),
.A2(n_817),
.B1(n_802),
.B2(n_929),
.C(n_979),
.Y(n_1132)
);

AOI211x1_ASAP7_75t_L g1133 ( 
.A1(n_997),
.A2(n_802),
.B(n_744),
.C(n_990),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_898),
.B(n_817),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_897),
.A2(n_938),
.A3(n_1003),
.B(n_1008),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_915),
.B(n_817),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_939),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_927),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1106),
.B(n_1121),
.C(n_1099),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1069),
.B(n_1067),
.Y(n_1140)
);

BUFx4f_ASAP7_75t_SL g1141 ( 
.A(n_1032),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1037),
.Y(n_1142)
);

OA21x2_ASAP7_75t_L g1143 ( 
.A1(n_1059),
.A2(n_1029),
.B(n_1132),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1091),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_1116),
.C(n_1136),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1112),
.B(n_1113),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1092),
.A2(n_1098),
.B(n_1096),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1117),
.A2(n_1130),
.B(n_1062),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1130),
.A2(n_1055),
.B(n_1068),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_1070),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1049),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1102),
.A2(n_1120),
.B(n_1023),
.Y(n_1152)
);

OAI222xp33_ASAP7_75t_L g1153 ( 
.A1(n_1053),
.A2(n_1038),
.B1(n_1134),
.B2(n_1063),
.C1(n_1025),
.C2(n_1020),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1110),
.A2(n_1123),
.B(n_1125),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1044),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1041),
.A2(n_1072),
.B(n_1042),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1022),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1047),
.A2(n_1060),
.B(n_1077),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1048),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1066),
.B(n_1035),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1090),
.A2(n_1028),
.B(n_1046),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1069),
.B(n_1067),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1107),
.B(n_1083),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1094),
.Y(n_1164)
);

BUFx10_ASAP7_75t_L g1165 ( 
.A(n_1124),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1027),
.B(n_1138),
.Y(n_1166)
);

AO21x2_ASAP7_75t_L g1167 ( 
.A1(n_1119),
.A2(n_1089),
.B(n_1024),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1064),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1115),
.A2(n_1126),
.B1(n_1079),
.B2(n_1076),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1026),
.A2(n_1133),
.A3(n_1105),
.B(n_1104),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1040),
.A2(n_1088),
.B(n_1085),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_1079),
.B(n_1108),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1056),
.A2(n_1042),
.B(n_1128),
.C(n_1030),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1128),
.B(n_1030),
.C(n_1133),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1039),
.B(n_1036),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1049),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1057),
.B(n_1054),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1034),
.A2(n_1019),
.B(n_1086),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1049),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1122),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1118),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1064),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1127),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1061),
.B(n_1097),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1061),
.B(n_1097),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1034),
.A2(n_1021),
.B(n_1109),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_1045),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1111),
.A2(n_1082),
.B(n_1087),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1084),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1100),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1080),
.A2(n_1122),
.B1(n_1043),
.B2(n_1071),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1050),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_1104),
.A2(n_1135),
.B(n_1074),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1058),
.B(n_1093),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1107),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1122),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1107),
.A2(n_1135),
.B(n_1104),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1137),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_SL g1199 ( 
.A(n_1078),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1095),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1033),
.A2(n_1135),
.B(n_1065),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1033),
.A2(n_1065),
.B(n_1114),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1074),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1081),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1033),
.A2(n_1065),
.B(n_1114),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1081),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1081),
.A2(n_1073),
.B(n_1095),
.Y(n_1208)
);

NOR3xp33_ASAP7_75t_L g1209 ( 
.A(n_1073),
.B(n_817),
.C(n_1106),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1059),
.A2(n_1029),
.B(n_1132),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1037),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1132),
.A2(n_1029),
.A3(n_1059),
.B(n_897),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1128),
.A2(n_817),
.B1(n_577),
.B2(n_425),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1049),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1051),
.B(n_817),
.C(n_1018),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1106),
.A2(n_817),
.B(n_1116),
.C(n_1099),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1049),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_1101),
.A2(n_1103),
.B(n_802),
.C(n_1106),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1099),
.A2(n_817),
.B(n_1121),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1112),
.B(n_817),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1059),
.A2(n_1029),
.B(n_1132),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1037),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1054),
.B(n_1057),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1064),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1091),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1091),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1099),
.A2(n_817),
.B(n_1121),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1112),
.A2(n_817),
.B1(n_1117),
.B2(n_1113),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1099),
.A2(n_817),
.B(n_1121),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1059),
.A2(n_1029),
.B(n_1132),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1059),
.A2(n_1029),
.B(n_1132),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1112),
.A2(n_817),
.B1(n_802),
.B2(n_1113),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1099),
.A2(n_817),
.B(n_1121),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1058),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1075),
.A2(n_1037),
.B(n_1031),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1112),
.A2(n_817),
.B1(n_802),
.B2(n_1113),
.Y(n_1236)
);

AO21x1_ASAP7_75t_L g1237 ( 
.A1(n_1106),
.A2(n_817),
.B(n_1116),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1069),
.B(n_1067),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1075),
.A2(n_1037),
.B(n_1031),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1099),
.A2(n_817),
.B(n_1121),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1037),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1112),
.B(n_817),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1091),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1091),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1106),
.A2(n_817),
.B(n_802),
.C(n_1099),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_817),
.B(n_1121),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1031),
.A2(n_1075),
.B(n_1037),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1049),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1112),
.B(n_1113),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1112),
.A2(n_817),
.B1(n_802),
.B2(n_1113),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1027),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1091),
.Y(n_1252)
);

BUFx2_ASAP7_75t_SL g1253 ( 
.A(n_1049),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1223),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1220),
.B(n_1242),
.Y(n_1255)
);

O2A1O1Ixp5_ASAP7_75t_L g1256 ( 
.A1(n_1237),
.A2(n_1216),
.B(n_1227),
.C(n_1246),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1152),
.A2(n_1218),
.B(n_1145),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1232),
.A2(n_1250),
.B1(n_1236),
.B2(n_1242),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1140),
.B(n_1162),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1232),
.A2(n_1236),
.B1(n_1250),
.B2(n_1220),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1195),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1216),
.A2(n_1218),
.B(n_1245),
.C(n_1209),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1150),
.A2(n_1160),
.B(n_1149),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1177),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1209),
.A2(n_1153),
.B(n_1215),
.C(n_1219),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1178),
.A2(n_1156),
.B(n_1186),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1228),
.B(n_1146),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1215),
.A2(n_1233),
.B(n_1240),
.C(n_1229),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1213),
.A2(n_1249),
.B1(n_1173),
.B2(n_1175),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1141),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1148),
.B(n_1173),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1174),
.A2(n_1169),
.B1(n_1172),
.B2(n_1139),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1187),
.B(n_1194),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1172),
.A2(n_1160),
.B1(n_1234),
.B2(n_1208),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1195),
.A2(n_1200),
.B(n_1238),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1251),
.Y(n_1276)
);

AND2x4_ASAP7_75t_SL g1277 ( 
.A(n_1165),
.B(n_1200),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1190),
.B(n_1226),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1143),
.B(n_1210),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1155),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1251),
.B(n_1191),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1202),
.A2(n_1197),
.B(n_1161),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1143),
.B(n_1210),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1140),
.B(n_1162),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1184),
.B(n_1185),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1143),
.B(n_1221),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1164),
.A2(n_1181),
.B1(n_1183),
.B2(n_1230),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1141),
.Y(n_1289)
);

CKINVDCx12_ASAP7_75t_R g1290 ( 
.A(n_1253),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1171),
.A2(n_1238),
.B(n_1203),
.C(n_1206),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1221),
.A2(n_1230),
.B1(n_1231),
.B2(n_1225),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1192),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1243),
.B(n_1252),
.Y(n_1294)
);

BUFx2_ASAP7_75t_R g1295 ( 
.A(n_1192),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1144),
.A2(n_1244),
.B(n_1196),
.C(n_1179),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1165),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1189),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1231),
.B(n_1212),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1235),
.A2(n_1239),
.B(n_1211),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1248),
.A2(n_1193),
.B1(n_1198),
.B2(n_1151),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1165),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1195),
.A2(n_1176),
.B(n_1180),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1235),
.A2(n_1239),
.B(n_1222),
.Y(n_1304)
);

AOI221x1_ASAP7_75t_SL g1305 ( 
.A1(n_1205),
.A2(n_1207),
.B1(n_1201),
.B2(n_1204),
.C(n_1212),
.Y(n_1305)
);

AOI211xp5_ASAP7_75t_L g1306 ( 
.A1(n_1151),
.A2(n_1217),
.B(n_1214),
.C(n_1180),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1163),
.B(n_1176),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1163),
.Y(n_1308)
);

AOI221x1_ASAP7_75t_SL g1309 ( 
.A1(n_1212),
.A2(n_1248),
.B1(n_1217),
.B2(n_1214),
.C(n_1193),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1168),
.B(n_1224),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1168),
.Y(n_1311)
);

INVx5_ASAP7_75t_L g1312 ( 
.A(n_1182),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1199),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1199),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1188),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_SL g1316 ( 
.A1(n_1193),
.A2(n_1170),
.B1(n_1166),
.B2(n_1206),
.C(n_1167),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1157),
.A2(n_1147),
.B1(n_1170),
.B2(n_1158),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1154),
.B(n_1142),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1241),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1247),
.B(n_1184),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1213),
.A2(n_902),
.B1(n_800),
.B2(n_1220),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1160),
.A2(n_1103),
.B(n_1101),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1232),
.A2(n_1113),
.B1(n_1117),
.B2(n_1112),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1251),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1156),
.B(n_1232),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1223),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1156),
.B(n_1232),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1151),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1216),
.A2(n_817),
.B(n_1106),
.C(n_802),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1298),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1299),
.B(n_1279),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1320),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1267),
.B(n_1325),
.Y(n_1333)
);

OR2x6_ASAP7_75t_L g1334 ( 
.A(n_1263),
.B(n_1322),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1258),
.A2(n_1260),
.B1(n_1269),
.B2(n_1327),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1315),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1266),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1291),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1257),
.B(n_1266),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1288),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1288),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1317),
.A2(n_1279),
.B(n_1284),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1283),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1299),
.B(n_1287),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1300),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1304),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1304),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1292),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1301),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1267),
.B(n_1325),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1319),
.Y(n_1351)
);

NOR2xp67_ASAP7_75t_L g1352 ( 
.A(n_1271),
.B(n_1272),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1301),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1280),
.B(n_1281),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1316),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1256),
.A2(n_1327),
.B(n_1318),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1273),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1318),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1272),
.A2(n_1274),
.B(n_1294),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1329),
.A2(n_1268),
.B(n_1262),
.Y(n_1360)
);

AND2x6_ASAP7_75t_L g1361 ( 
.A(n_1259),
.B(n_1285),
.Y(n_1361)
);

OAI321xp33_ASAP7_75t_L g1362 ( 
.A1(n_1258),
.A2(n_1260),
.A3(n_1265),
.B1(n_1269),
.B2(n_1321),
.C(n_1323),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1274),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1324),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1305),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1254),
.B(n_1326),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1264),
.B(n_1278),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1309),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1323),
.B(n_1255),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1296),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1308),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1312),
.Y(n_1372)
);

OAI21xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1275),
.A2(n_1303),
.B(n_1310),
.Y(n_1373)
);

NAND2x1_ASAP7_75t_L g1374 ( 
.A(n_1334),
.B(n_1285),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1330),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1330),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1342),
.B(n_1307),
.Y(n_1378)
);

AND2x4_ASAP7_75t_SL g1379 ( 
.A(n_1334),
.B(n_1261),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1361),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1362),
.B(n_1360),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1345),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1358),
.B(n_1312),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1331),
.B(n_1286),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1358),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1333),
.B(n_1306),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1372),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1333),
.B(n_1277),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1344),
.B(n_1261),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1345),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1354),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1357),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1342),
.B(n_1314),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1350),
.B(n_1328),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1351),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1336),
.B(n_1311),
.Y(n_1396)
);

OA222x2_ASAP7_75t_L g1397 ( 
.A1(n_1393),
.A2(n_1339),
.B1(n_1334),
.B2(n_1337),
.C1(n_1365),
.C2(n_1340),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1379),
.Y(n_1398)
);

OAI211xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1381),
.A2(n_1360),
.B(n_1335),
.C(n_1369),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1375),
.Y(n_1400)
);

AOI221xp5_ASAP7_75t_L g1401 ( 
.A1(n_1381),
.A2(n_1362),
.B1(n_1369),
.B2(n_1335),
.C(n_1365),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1375),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1392),
.B(n_1357),
.Y(n_1403)
);

NOR4xp25_ASAP7_75t_SL g1404 ( 
.A(n_1385),
.B(n_1338),
.C(n_1353),
.D(n_1363),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1384),
.B(n_1353),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1392),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1348),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_SL g1408 ( 
.A(n_1386),
.B(n_1297),
.Y(n_1408)
);

AOI222xp33_ASAP7_75t_L g1409 ( 
.A1(n_1386),
.A2(n_1352),
.B1(n_1355),
.B2(n_1368),
.C1(n_1350),
.C2(n_1338),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1388),
.A2(n_1334),
.B1(n_1352),
.B2(n_1355),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1384),
.B(n_1332),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1378),
.B(n_1348),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1389),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1376),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1393),
.B(n_1370),
.C(n_1334),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1378),
.B(n_1393),
.Y(n_1416)
);

AO21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1395),
.A2(n_1368),
.B(n_1349),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1376),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1377),
.Y(n_1419)
);

AOI222xp33_ASAP7_75t_L g1420 ( 
.A1(n_1394),
.A2(n_1363),
.B1(n_1349),
.B2(n_1370),
.C1(n_1341),
.C2(n_1340),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1395),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

OAI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1388),
.A2(n_1334),
.B1(n_1373),
.B2(n_1366),
.C(n_1367),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1396),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1389),
.B(n_1332),
.Y(n_1425)
);

NAND2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1374),
.B(n_1302),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1382),
.A2(n_1346),
.B(n_1347),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1380),
.B(n_1332),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1380),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1374),
.A2(n_1373),
.B1(n_1366),
.B2(n_1367),
.C(n_1289),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1389),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1426),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1427),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1400),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1400),
.Y(n_1435)
);

INVx4_ASAP7_75t_SL g1436 ( 
.A(n_1428),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1415),
.A2(n_1347),
.B(n_1343),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1402),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1397),
.B(n_1385),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1429),
.Y(n_1440)
);

INVx4_ASAP7_75t_SL g1441 ( 
.A(n_1428),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1421),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1420),
.B(n_1407),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1428),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1414),
.Y(n_1445)
);

AND2x6_ASAP7_75t_SL g1446 ( 
.A(n_1403),
.B(n_1295),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1399),
.B(n_1364),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1418),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1407),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1416),
.A2(n_1343),
.B(n_1390),
.Y(n_1450)
);

AND2x4_ASAP7_75t_SL g1451 ( 
.A(n_1398),
.B(n_1383),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1417),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1412),
.B(n_1391),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_SL g1454 ( 
.A(n_1417),
.B(n_1387),
.Y(n_1454)
);

INVx4_ASAP7_75t_SL g1455 ( 
.A(n_1424),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1436),
.B(n_1429),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1445),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1449),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1445),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1436),
.B(n_1397),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_L g1461 ( 
.A(n_1432),
.B(n_1430),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1449),
.B(n_1412),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1436),
.B(n_1405),
.Y(n_1463)
);

NAND4xp25_ASAP7_75t_L g1464 ( 
.A(n_1443),
.B(n_1401),
.C(n_1409),
.D(n_1410),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1436),
.B(n_1405),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1448),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1448),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1447),
.A2(n_1423),
.B(n_1363),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1442),
.B(n_1419),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1442),
.B(n_1422),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1439),
.B(n_1404),
.C(n_1408),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.B(n_1455),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1434),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_1411),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1452),
.B(n_1374),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1439),
.B(n_1411),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1446),
.B(n_1276),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1450),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1452),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1429),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1450),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1441),
.B(n_1425),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1450),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1450),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1452),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1434),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1446),
.B(n_1276),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1450),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1441),
.B(n_1425),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1435),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1433),
.Y(n_1492)
);

NAND4xp75_ASAP7_75t_L g1493 ( 
.A(n_1440),
.B(n_1359),
.C(n_1356),
.D(n_1282),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1478),
.B(n_1432),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1464),
.B(n_1444),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1472),
.B(n_1444),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1461),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1461),
.A2(n_1406),
.B(n_1440),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1487),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1472),
.B(n_1455),
.Y(n_1500)
);

NOR2x1_ASAP7_75t_L g1501 ( 
.A(n_1471),
.B(n_1452),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1487),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1475),
.B(n_1452),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1473),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1475),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1431),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1474),
.B(n_1455),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1474),
.B(n_1455),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1471),
.B(n_1452),
.C(n_1371),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1481),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1458),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1458),
.B(n_1453),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1457),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1473),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1491),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1492),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1457),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1492),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1491),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1459),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1474),
.B(n_1477),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1468),
.B(n_1413),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1488),
.B(n_1455),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1462),
.B(n_1438),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1459),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1477),
.B(n_1455),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1460),
.B(n_1451),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1462),
.B(n_1438),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1505),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1504),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1497),
.A2(n_1509),
.B(n_1498),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1501),
.B(n_1480),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1501),
.A2(n_1468),
.B1(n_1493),
.B2(n_1460),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1507),
.B(n_1456),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1504),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1511),
.B(n_1477),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1514),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1514),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1495),
.A2(n_1454),
.B1(n_1437),
.B2(n_1486),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1496),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1503),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1503),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1515),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1515),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1496),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1521),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1519),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1519),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1512),
.B(n_1506),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1521),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_1463),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1513),
.Y(n_1553)
);

AOI21xp33_ASAP7_75t_L g1554 ( 
.A1(n_1531),
.A2(n_1494),
.B(n_1510),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1533),
.A2(n_1523),
.B(n_1493),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1529),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1532),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1547),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1541),
.A2(n_1527),
.B1(n_1522),
.B2(n_1526),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1547),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1546),
.Y(n_1561)
);

OAI32xp33_ASAP7_75t_L g1562 ( 
.A1(n_1532),
.A2(n_1486),
.A3(n_1480),
.B1(n_1517),
.B2(n_1502),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1550),
.A2(n_1500),
.B(n_1508),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1551),
.Y(n_1564)
);

OAI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1540),
.A2(n_1512),
.B1(n_1500),
.B2(n_1508),
.C(n_1526),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1534),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1567)
);

AOI31xp33_ASAP7_75t_L g1568 ( 
.A1(n_1553),
.A2(n_1293),
.A3(n_1476),
.B(n_1313),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1551),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1520),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1535),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1558),
.Y(n_1573)
);

AOI222xp33_ASAP7_75t_L g1574 ( 
.A1(n_1556),
.A2(n_1536),
.B1(n_1548),
.B2(n_1545),
.C1(n_1544),
.C2(n_1549),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1567),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1560),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1566),
.B(n_1534),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1567),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1556),
.Y(n_1579)
);

NOR3xp33_ASAP7_75t_L g1580 ( 
.A(n_1554),
.B(n_1543),
.C(n_1538),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1561),
.B(n_1538),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1563),
.B(n_1543),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1568),
.B(n_1542),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1564),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1575),
.B(n_1569),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1579),
.B(n_1559),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1580),
.A2(n_1565),
.B1(n_1557),
.B2(n_1540),
.C(n_1571),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1581),
.B(n_1542),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1582),
.A2(n_1562),
.B1(n_1555),
.B2(n_1572),
.C(n_1570),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1577),
.A2(n_1476),
.B1(n_1456),
.B2(n_1463),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_SL g1591 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1578),
.A2(n_1570),
.B1(n_1539),
.B2(n_1537),
.C(n_1499),
.Y(n_1592)
);

OAI31xp33_ASAP7_75t_L g1593 ( 
.A1(n_1573),
.A2(n_1502),
.A3(n_1499),
.B(n_1520),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1576),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1585),
.Y(n_1595)
);

XNOR2x1_ASAP7_75t_L g1596 ( 
.A(n_1588),
.B(n_1584),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1591),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1586),
.Y(n_1598)
);

AOI211xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1587),
.A2(n_1525),
.B(n_1574),
.C(n_1518),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1589),
.A2(n_1456),
.B1(n_1476),
.B2(n_1525),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1596),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1595),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1597),
.B(n_1574),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1598),
.B(n_1599),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1600),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1596),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1604),
.B(n_1594),
.C(n_1592),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1601),
.Y(n_1608)
);

AOI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1606),
.A2(n_1593),
.B1(n_1590),
.B2(n_1518),
.C(n_1516),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1603),
.A2(n_1516),
.B1(n_1466),
.B2(n_1467),
.C(n_1492),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1605),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1608),
.Y(n_1612)
);

AOI211xp5_ASAP7_75t_L g1613 ( 
.A1(n_1607),
.A2(n_1602),
.B(n_1481),
.C(n_1456),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1611),
.Y(n_1614)
);

XNOR2x1_ASAP7_75t_L g1615 ( 
.A(n_1612),
.B(n_1609),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_1613),
.B1(n_1614),
.B2(n_1610),
.C(n_1476),
.Y(n_1616)
);

OAI22x1_ASAP7_75t_L g1617 ( 
.A1(n_1616),
.A2(n_1467),
.B1(n_1466),
.B2(n_1528),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_R g1618 ( 
.A1(n_1616),
.A2(n_1479),
.B1(n_1489),
.B2(n_1485),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1617),
.B(n_1524),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1618),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1620),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1619),
.A2(n_1270),
.B1(n_1290),
.B2(n_1528),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1622),
.Y(n_1623)
);

NAND2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1623),
.B(n_1621),
.Y(n_1624)
);

AND3x1_ASAP7_75t_L g1625 ( 
.A(n_1624),
.B(n_1490),
.C(n_1483),
.Y(n_1625)
);

OAI22x1_ASAP7_75t_L g1626 ( 
.A1(n_1625),
.A2(n_1524),
.B1(n_1440),
.B2(n_1465),
.Y(n_1626)
);

AOI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1626),
.A2(n_1479),
.B1(n_1482),
.B2(n_1489),
.C(n_1484),
.Y(n_1627)
);

AOI211xp5_ASAP7_75t_L g1628 ( 
.A1(n_1627),
.A2(n_1470),
.B(n_1469),
.C(n_1483),
.Y(n_1628)
);


endmodule