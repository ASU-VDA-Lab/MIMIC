module real_jpeg_19875_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_0),
.A2(n_30),
.B1(n_57),
.B2(n_58),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_70),
.B1(n_74),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_3),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_137),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_137),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_137),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_4),
.B(n_72),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_4),
.A2(n_14),
.B(n_29),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_125),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_83),
.B1(n_84),
.B2(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_4),
.B(n_57),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_4),
.A2(n_57),
.B(n_223),
.Y(n_227)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_36),
.B1(n_70),
.B2(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_7),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_8),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_75),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_75),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_75),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_70),
.B1(n_74),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_110),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_110),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_110),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_127)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_69),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_140),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_19),
.B(n_112),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_91),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_79),
.B2(n_80),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_37),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_25),
.A2(n_84),
.B(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_28),
.B(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_31),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_31),
.A2(n_35),
.B(n_102),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_33),
.A2(n_83),
.B1(n_183),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_34),
.A2(n_83),
.B(n_186),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_38),
.A2(n_48),
.B(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_38),
.A2(n_87),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_38),
.A2(n_44),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_38),
.A2(n_44),
.B1(n_194),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_38),
.A2(n_44),
.B1(n_214),
.B2(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_38),
.A2(n_230),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_40),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

AOI32xp33_ASAP7_75t_L g222 ( 
.A1(n_39),
.A2(n_55),
.A3(n_58),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_40),
.A2(n_45),
.B(n_125),
.C(n_190),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_40),
.B(n_53),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_44),
.A2(n_46),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_44),
.B(n_125),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_59),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_53),
.B(n_57),
.C(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_52),
.B(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_52),
.A2(n_61),
.B1(n_131),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_52),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_52),
.A2(n_61),
.B1(n_171),
.B2(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.Y(n_62)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_69),
.Y(n_123)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_58),
.A2(n_71),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_60),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_73),
.B(n_76),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_73),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_109),
.B1(n_111),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_68),
.A2(n_72),
.B1(n_124),
.B2(n_136),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_125),
.CON(n_124),
.SN(n_124)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_83),
.A2(n_100),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_84),
.B(n_125),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_89),
.B(n_150),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_103),
.C(n_107),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_93),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_119),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_113),
.A2(n_117),
.B1(n_118),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_113),
.Y(n_259)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_119),
.A2(n_120),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_129),
.C(n_133),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_126),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_174),
.B(n_254),
.C(n_260),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_159),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_142),
.B(n_159),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_155),
.B2(n_158),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_145),
.B(n_146),
.C(n_158),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_154),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_160),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_169),
.B(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_253),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_248),
.B(n_252),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_235),
.B(n_247),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_217),
.B(n_234),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_206),
.B(n_216),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_195),
.B(n_205),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_187),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_191),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_200),
.B(n_204),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_219),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_225),
.B1(n_232),
.B2(n_233),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_226),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_231),
.C(n_232),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_237),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_244),
.C(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);


endmodule