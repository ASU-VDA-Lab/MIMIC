module fake_ariane_3148_n_1382 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1382);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1382;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_169),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_185),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_181),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_254),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_160),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_70),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_71),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_106),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_213),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_2),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_111),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_252),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_153),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_69),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_103),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_75),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_101),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_266),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_47),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_212),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_269),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_286),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_315),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_172),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_268),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_229),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_36),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_238),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_83),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_54),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_215),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_115),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_236),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_150),
.Y(n_368)
);

BUFx2_ASAP7_75t_SL g369 ( 
.A(n_250),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_73),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_211),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_167),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_151),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_291),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_133),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_277),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_145),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_178),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_143),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_264),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_2),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_180),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_44),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_201),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_191),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_72),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_5),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_61),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_41),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_239),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_64),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_95),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_32),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_179),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_159),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_33),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_273),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_287),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_293),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_128),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_23),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_30),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_99),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_38),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_207),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_270),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_127),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_146),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_177),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_161),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_194),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_156),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_86),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_199),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_305),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_5),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_56),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_261),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_14),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_81),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_7),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_90),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_313),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_97),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_162),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_158),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_125),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_136),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_142),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_288),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_205),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_193),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_93),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_85),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_68),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_281),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_255),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_296),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_248),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_304),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_274),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_321),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_168),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_314),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_306),
.Y(n_448)
);

CKINVDCx11_ASAP7_75t_R g449 ( 
.A(n_307),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_55),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_208),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_198),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_39),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_200),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_11),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_3),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_122),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_59),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_138),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_45),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_272),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_9),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_189),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_282),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_182),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_311),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_82),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_15),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_107),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_183),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_187),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_4),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_76),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_309),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_230),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_114),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_20),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_329),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_192),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_249),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_224),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_26),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_108),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_109),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_131),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_34),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_104),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_23),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_197),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_36),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_102),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_251),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_290),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_80),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_84),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_126),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_223),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_144),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_14),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_279),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_37),
.Y(n_501)
);

BUFx8_ASAP7_75t_SL g502 ( 
.A(n_231),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_147),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_11),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_292),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_94),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_19),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_31),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_100),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_218),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_298),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_220),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_166),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_352),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_388),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_404),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_450),
.B(n_0),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_404),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_473),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_502),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_459),
.B(n_40),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_449),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_0),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_404),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_361),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_468),
.Y(n_530)
);

INVxp33_ASAP7_75t_SL g531 ( 
.A(n_462),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_398),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_337),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_499),
.Y(n_535)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_342),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_370),
.B(n_1),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_456),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_356),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_472),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_366),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_400),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_414),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_460),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_497),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_512),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_474),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_492),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_403),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_382),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_395),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_418),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_424),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_455),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_488),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_421),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_507),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_333),
.B(n_1),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_410),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_335),
.B(n_3),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_410),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_423),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_430),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_430),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_508),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_434),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_336),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_480),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_341),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_369),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_346),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_347),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_350),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_355),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_363),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_368),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_470),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_470),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_372),
.B(n_4),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_373),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_379),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_470),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_381),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_330),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_331),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_383),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_334),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_338),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_339),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_340),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_384),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_343),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_344),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_348),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_475),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_389),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_390),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_392),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_349),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_475),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_351),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_393),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_353),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_354),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_394),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_515),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_516),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_585),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_519),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_521),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_586),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_608),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_576),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_528),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_529),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_533),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_540),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_594),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_531),
.A2(n_443),
.B1(n_457),
.B2(n_401),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_542),
.Y(n_632)
);

CKINVDCx8_ASAP7_75t_R g633 ( 
.A(n_522),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_599),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_546),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_547),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_568),
.B(n_443),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_550),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_557),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_551),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_561),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_538),
.Y(n_650)
);

NAND2x1_ASAP7_75t_L g651 ( 
.A(n_569),
.B(n_475),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_575),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_523),
.B(n_345),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_544),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_613),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_554),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_535),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_527),
.A2(n_465),
.B1(n_433),
.B2(n_435),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_592),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_580),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_581),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_565),
.B(n_332),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_583),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_514),
.B(n_402),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_589),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_591),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_520),
.B(n_422),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_554),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_610),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_567),
.A2(n_444),
.B(n_425),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_590),
.B(n_454),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_588),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_555),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_603),
.B(n_463),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_534),
.B(n_539),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_570),
.B(n_442),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_579),
.B(n_578),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_572),
.B(n_464),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_520),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_537),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_564),
.B(n_357),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_518),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_518),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_593),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_574),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_598),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_602),
.B(n_513),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_SL g697 ( 
.A(n_600),
.B(n_466),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_614),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_648),
.B(n_556),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_615),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_693),
.B(n_536),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_633),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_695),
.B(n_607),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_643),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_654),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_648),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_636),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_687),
.B(n_609),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_643),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_619),
.B(n_611),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_696),
.B(n_558),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_626),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_627),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_630),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_653),
.A2(n_600),
.B1(n_601),
.B2(n_573),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_628),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_660),
.B(n_332),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_632),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_679),
.B(n_595),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_682),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_684),
.B(n_548),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_687),
.B(n_559),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_560),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_687),
.B(n_562),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_684),
.B(n_549),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_635),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_637),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_636),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_638),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_640),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_696),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_636),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_692),
.B(n_596),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_623),
.B(n_601),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_643),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_660),
.B(n_597),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_643),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_692),
.B(n_612),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_692),
.B(n_552),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_688),
.B(n_526),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_623),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_642),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_644),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_644),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_636),
.Y(n_746)
);

AND2x6_ASAP7_75t_L g747 ( 
.A(n_681),
.B(n_332),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_692),
.B(n_553),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_644),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_619),
.B(n_476),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_647),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_661),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_624),
.B(n_484),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_661),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_665),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_644),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_670),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_665),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_649),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_658),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_670),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_667),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_624),
.B(n_485),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_667),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_511),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_616),
.B(n_360),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_652),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_670),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_618),
.B(n_415),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_639),
.B(n_566),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_658),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_681),
.B(n_332),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_629),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_655),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_656),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_625),
.B(n_478),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_670),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_629),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_689),
.B(n_494),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_679),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_685),
.B(n_571),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_688),
.B(n_639),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_646),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_689),
.B(n_405),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_666),
.B(n_541),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_634),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_662),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_709),
.B(n_691),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_706),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_702),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_723),
.A2(n_653),
.B1(n_697),
.B2(n_677),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_713),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_714),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_722),
.B(n_694),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_705),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_SL g797 ( 
.A1(n_783),
.A2(n_551),
.B1(n_646),
.B2(n_545),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_724),
.B(n_677),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_725),
.B(n_680),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_705),
.B(n_645),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_719),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_727),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_780),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_735),
.B(n_674),
.Y(n_804)
);

AO22x2_ASAP7_75t_L g805 ( 
.A1(n_726),
.A2(n_770),
.B1(n_748),
.B2(n_739),
.Y(n_805)
);

AO22x2_ASAP7_75t_L g806 ( 
.A1(n_785),
.A2(n_737),
.B1(n_735),
.B2(n_782),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_782),
.B(n_699),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_728),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_732),
.B(n_690),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_730),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_734),
.A2(n_631),
.B1(n_680),
.B2(n_686),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_703),
.B(n_742),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_701),
.B(n_650),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_732),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_731),
.Y(n_815)
);

BUFx8_ASAP7_75t_L g816 ( 
.A(n_771),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_778),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_742),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_767),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_774),
.Y(n_821)
);

OR2x2_ASAP7_75t_SL g822 ( 
.A(n_715),
.B(n_741),
.Y(n_822)
);

NAND2x1p5_ASAP7_75t_L g823 ( 
.A(n_760),
.B(n_664),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_775),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_707),
.B(n_697),
.Y(n_825)
);

AO22x2_ASAP7_75t_L g826 ( 
.A1(n_781),
.A2(n_683),
.B1(n_659),
.B2(n_671),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_752),
.A2(n_683),
.B1(n_686),
.B2(n_641),
.Y(n_827)
);

OAI221xp5_ASAP7_75t_L g828 ( 
.A1(n_787),
.A2(n_675),
.B1(n_668),
.B2(n_672),
.C(n_669),
.Y(n_828)
);

AO22x2_ASAP7_75t_L g829 ( 
.A1(n_712),
.A2(n_678),
.B1(n_641),
.B2(n_634),
.Y(n_829)
);

AND2x2_ASAP7_75t_SL g830 ( 
.A(n_716),
.B(n_663),
.Y(n_830)
);

OR2x2_ASAP7_75t_SL g831 ( 
.A(n_720),
.B(n_657),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_754),
.Y(n_832)
);

OR2x6_ASAP7_75t_SL g833 ( 
.A(n_711),
.B(n_358),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_740),
.B(n_617),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_755),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_758),
.Y(n_836)
);

NOR2xp67_ASAP7_75t_L g837 ( 
.A(n_745),
.B(n_757),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_711),
.B(n_673),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_779),
.A2(n_663),
.B1(n_621),
.B2(n_620),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_749),
.B(n_761),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_698),
.B(n_651),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_764),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_751),
.B(n_676),
.Y(n_844)
);

OAI221xp5_ASAP7_75t_L g845 ( 
.A1(n_700),
.A2(n_510),
.B1(n_509),
.B2(n_506),
.C(n_505),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_779),
.B(n_359),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_759),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_765),
.B(n_362),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_773),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_786),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_750),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_750),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_768),
.B(n_405),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_718),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_745),
.B(n_364),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_765),
.B(n_365),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_757),
.A2(n_371),
.B1(n_374),
.B2(n_367),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_753),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_704),
.B(n_375),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_704),
.B(n_376),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_753),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_721),
.B(n_784),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_763),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_710),
.A2(n_378),
.B1(n_380),
.B2(n_377),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_778),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_763),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_708),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_784),
.B(n_6),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_710),
.A2(n_386),
.B1(n_387),
.B2(n_385),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_766),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_736),
.B(n_391),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_766),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_736),
.B(n_405),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_729),
.Y(n_875)
);

OAI221xp5_ASAP7_75t_L g876 ( 
.A1(n_769),
.A2(n_503),
.B1(n_498),
.B2(n_496),
.C(n_495),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_777),
.B(n_6),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_769),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_738),
.B(n_396),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_776),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_733),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_776),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_796),
.B(n_738),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_788),
.B(n_744),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_798),
.B(n_744),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_807),
.B(n_777),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_807),
.B(n_799),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_813),
.B(n_791),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_851),
.B(n_756),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_803),
.B(n_746),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_852),
.B(n_718),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_812),
.B(n_397),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_789),
.B(n_399),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_825),
.B(n_407),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_823),
.B(n_408),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_814),
.B(n_409),
.Y(n_896)
);

AND3x1_ASAP7_75t_L g897 ( 
.A(n_792),
.B(n_7),
.C(n_8),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_858),
.B(n_718),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_861),
.B(n_718),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_SL g900 ( 
.A(n_809),
.B(n_793),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_800),
.B(n_411),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_794),
.B(n_747),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_SL g903 ( 
.A(n_795),
.B(n_412),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_863),
.B(n_413),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_866),
.B(n_417),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_830),
.B(n_811),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_SL g907 ( 
.A(n_801),
.B(n_419),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_838),
.B(n_747),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_871),
.B(n_747),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_848),
.B(n_420),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_873),
.B(n_878),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_856),
.B(n_426),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_880),
.B(n_747),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_SL g914 ( 
.A(n_802),
.B(n_427),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_SL g915 ( 
.A(n_808),
.B(n_428),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_834),
.B(n_429),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_834),
.B(n_431),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_882),
.B(n_772),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_862),
.B(n_819),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_822),
.B(n_8),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_790),
.B(n_432),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_846),
.B(n_436),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_810),
.B(n_772),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_877),
.B(n_437),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_815),
.B(n_772),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_877),
.B(n_438),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_857),
.B(n_818),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_820),
.B(n_439),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_SL g929 ( 
.A(n_821),
.B(n_824),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_SL g930 ( 
.A(n_869),
.B(n_440),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_864),
.B(n_441),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_SL g932 ( 
.A(n_841),
.B(n_445),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_870),
.B(n_446),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_804),
.B(n_816),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_816),
.B(n_447),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_827),
.B(n_772),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_832),
.B(n_448),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_835),
.B(n_451),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_855),
.B(n_452),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_836),
.B(n_458),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_837),
.B(n_461),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_859),
.B(n_854),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_842),
.B(n_467),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_843),
.B(n_469),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_860),
.B(n_471),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_872),
.B(n_479),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_879),
.B(n_481),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_840),
.B(n_483),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_844),
.B(n_405),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_844),
.B(n_416),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_SL g951 ( 
.A(n_817),
.B(n_865),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_867),
.B(n_416),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_888),
.B(n_876),
.C(n_845),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_SL g954 ( 
.A(n_930),
.B(n_828),
.C(n_839),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_887),
.B(n_797),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_949),
.A2(n_874),
.B(n_868),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_949),
.A2(n_875),
.B(n_881),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_911),
.A2(n_885),
.B(n_892),
.Y(n_958)
);

NAND3x1_ASAP7_75t_L g959 ( 
.A(n_902),
.B(n_833),
.C(n_847),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_889),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_929),
.A2(n_912),
.B(n_910),
.Y(n_961)
);

NOR2x1_ASAP7_75t_SL g962 ( 
.A(n_942),
.B(n_849),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_920),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_SL g964 ( 
.A1(n_922),
.A2(n_850),
.B(n_831),
.C(n_829),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_906),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_927),
.B(n_805),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_919),
.B(n_805),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_886),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_934),
.B(n_883),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_916),
.A2(n_806),
.B1(n_826),
.B2(n_829),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_917),
.B(n_853),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_890),
.Y(n_972)
);

AO31x2_ASAP7_75t_L g973 ( 
.A1(n_936),
.A2(n_806),
.A3(n_826),
.B(n_489),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_891),
.A2(n_491),
.B(n_487),
.Y(n_974)
);

BUFx4_ASAP7_75t_SL g975 ( 
.A(n_935),
.Y(n_975)
);

NOR4xp25_ASAP7_75t_L g976 ( 
.A(n_894),
.B(n_9),
.C(n_10),
.D(n_12),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_924),
.B(n_10),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_923),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_926),
.B(n_12),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_898),
.A2(n_493),
.B(n_13),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_950),
.A2(n_43),
.B(n_42),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_900),
.A2(n_489),
.B(n_416),
.C(n_16),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_897),
.A2(n_489),
.B1(n_416),
.B2(n_16),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_899),
.A2(n_13),
.B(n_15),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_SL g985 ( 
.A1(n_950),
.A2(n_489),
.B(n_48),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_937),
.B(n_17),
.Y(n_986)
);

NOR4xp25_ASAP7_75t_L g987 ( 
.A(n_895),
.B(n_17),
.C(n_18),
.D(n_19),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_903),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_893),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_948),
.B(n_46),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_938),
.B(n_21),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_940),
.B(n_22),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_SL g993 ( 
.A1(n_921),
.A2(n_22),
.B(n_24),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_952),
.A2(n_50),
.B(n_49),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_909),
.A2(n_52),
.B(n_51),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_925),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_884),
.A2(n_57),
.B(n_53),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_945),
.A2(n_60),
.B(n_58),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_907),
.B(n_24),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_896),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_913),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_918),
.A2(n_63),
.B(n_62),
.Y(n_1002)
);

NAND3x1_ASAP7_75t_L g1003 ( 
.A(n_908),
.B(n_25),
.C(n_26),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_952),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_904),
.A2(n_25),
.B(n_27),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_SL g1006 ( 
.A1(n_905),
.A2(n_27),
.B(n_28),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_946),
.A2(n_66),
.B(n_65),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_901),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_951),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_928),
.B(n_28),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_932),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_943),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_941),
.A2(n_939),
.B(n_947),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_965),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_972),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_963),
.B(n_914),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1004),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_995),
.A2(n_1002),
.B(n_956),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_SL g1019 ( 
.A(n_953),
.B(n_931),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_969),
.B(n_944),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_953),
.A2(n_933),
.B1(n_915),
.B2(n_31),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_989),
.B(n_29),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_957),
.A2(n_74),
.B(n_67),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_981),
.A2(n_78),
.B(n_77),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_968),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_958),
.A2(n_87),
.B(n_79),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_997),
.A2(n_89),
.B(n_88),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_994),
.A2(n_219),
.B(n_327),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_967),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_988),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_SL g1031 ( 
.A1(n_962),
.A2(n_33),
.B(n_34),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_955),
.B(n_35),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_960),
.Y(n_1033)
);

OA21x2_ASAP7_75t_L g1034 ( 
.A1(n_984),
.A2(n_222),
.B(n_325),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_1007),
.A2(n_221),
.B(n_323),
.Y(n_1035)
);

BUFx2_ASAP7_75t_R g1036 ( 
.A(n_1000),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_966),
.B(n_1011),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_978),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_1001),
.A2(n_217),
.B(n_322),
.Y(n_1039)
);

INVx6_ASAP7_75t_L g1040 ( 
.A(n_972),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_996),
.A2(n_216),
.B(n_319),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1012),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_954),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_986),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_1006),
.A2(n_226),
.B(n_91),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_961),
.A2(n_227),
.B(n_92),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_991),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_977),
.B(n_39),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_992),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_979),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_982),
.A2(n_96),
.A3(n_98),
.B(n_105),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_972),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_983),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_998),
.A2(n_116),
.A3(n_117),
.B(n_118),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_974),
.A2(n_119),
.B(n_120),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_1010),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_983),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_969),
.Y(n_1058)
);

AO21x2_ASAP7_75t_L g1059 ( 
.A1(n_980),
.A2(n_129),
.B(n_130),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1011),
.B(n_328),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_1013),
.A2(n_132),
.B(n_134),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_973),
.A2(n_135),
.A3(n_137),
.B(n_139),
.Y(n_1062)
);

OA21x2_ASAP7_75t_L g1063 ( 
.A1(n_970),
.A2(n_140),
.B(n_141),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_964),
.A2(n_148),
.B(n_149),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_SL g1065 ( 
.A(n_993),
.B(n_999),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_977),
.B(n_318),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1005),
.A2(n_1009),
.B1(n_1008),
.B2(n_971),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_959),
.B(n_152),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_990),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_985),
.A2(n_154),
.B(n_155),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1029),
.B(n_973),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1017),
.B(n_973),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1017),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_1018),
.A2(n_1003),
.B(n_976),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1014),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1038),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1033),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1025),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1062),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1062),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1036),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1023),
.A2(n_987),
.B(n_163),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1062),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1042),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1058),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1061),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1037),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1054),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1056),
.B(n_975),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1054),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_1060),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1016),
.B(n_157),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1051),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1050),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1046),
.A2(n_164),
.B(n_165),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1052),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1044),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1043),
.A2(n_170),
.B(n_171),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1047),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1049),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1035),
.A2(n_173),
.B(n_174),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1048),
.B(n_175),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1040),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1067),
.B(n_176),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1054),
.Y(n_1105)
);

NAND2x1_ASAP7_75t_L g1106 ( 
.A(n_1019),
.B(n_184),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1021),
.A2(n_188),
.B1(n_190),
.B2(n_195),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1040),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1019),
.A2(n_316),
.B(n_202),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1060),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1015),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1020),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1039),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1020),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1031),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1051),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1041),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1051),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1055),
.A2(n_196),
.B(n_203),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1034),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1045),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1034),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1069),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1032),
.B(n_312),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1063),
.Y(n_1125)
);

INVx6_ASAP7_75t_L g1126 ( 
.A(n_1065),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1066),
.B(n_204),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1028),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1069),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1063),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1024),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1022),
.B(n_206),
.Y(n_1132)
);

OA21x2_ASAP7_75t_L g1133 ( 
.A1(n_1064),
.A2(n_1027),
.B(n_1026),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_1103),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_1081),
.B(n_1068),
.Y(n_1135)
);

INVxp33_ASAP7_75t_SL g1136 ( 
.A(n_1081),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1114),
.B(n_1057),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1111),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1114),
.B(n_1053),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1097),
.B(n_1065),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1075),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_R g1142 ( 
.A(n_1132),
.B(n_1092),
.Y(n_1142)
);

BUFx10_ASAP7_75t_L g1143 ( 
.A(n_1108),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1111),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_1099),
.Y(n_1145)
);

XOR2xp5_ASAP7_75t_L g1146 ( 
.A(n_1089),
.B(n_209),
.Y(n_1146)
);

BUFx8_ASAP7_75t_SL g1147 ( 
.A(n_1129),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1091),
.B(n_1070),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1078),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1091),
.B(n_1059),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1100),
.B(n_1094),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1129),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_1126),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1091),
.B(n_210),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1087),
.B(n_1030),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_1126),
.B(n_214),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_R g1157 ( 
.A(n_1110),
.B(n_225),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1087),
.B(n_228),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_1110),
.B(n_232),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1077),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1078),
.Y(n_1161)
);

NAND2xp33_ASAP7_75t_R g1162 ( 
.A(n_1110),
.B(n_233),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1075),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_R g1164 ( 
.A(n_1126),
.B(n_1123),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1084),
.B(n_234),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1073),
.B(n_235),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_R g1167 ( 
.A(n_1102),
.B(n_237),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1112),
.B(n_240),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1073),
.B(n_241),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1123),
.B(n_242),
.Y(n_1170)
);

NAND2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1106),
.B(n_243),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_R g1172 ( 
.A(n_1102),
.B(n_244),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1124),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_1126),
.B(n_245),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1123),
.Y(n_1175)
);

NAND2xp33_ASAP7_75t_R g1176 ( 
.A(n_1127),
.B(n_246),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1085),
.Y(n_1177)
);

NAND2xp33_ASAP7_75t_R g1178 ( 
.A(n_1127),
.B(n_247),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1096),
.B(n_253),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_1109),
.B(n_257),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1104),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1076),
.B(n_258),
.Y(n_1182)
);

XNOR2xp5_ASAP7_75t_L g1183 ( 
.A(n_1076),
.B(n_259),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1115),
.B(n_260),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1072),
.B(n_262),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1106),
.B(n_263),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_R g1187 ( 
.A(n_1109),
.B(n_265),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1072),
.B(n_267),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1071),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1071),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1074),
.B(n_271),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1098),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1152),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1144),
.B(n_1093),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1141),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1181),
.B(n_1122),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1145),
.B(n_1093),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1140),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1149),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1163),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1151),
.B(n_1118),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1161),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1177),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1160),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1189),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1138),
.B(n_1116),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1190),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1134),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1155),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1166),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1137),
.B(n_1118),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1143),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1150),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1148),
.B(n_1116),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1137),
.B(n_1088),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_1192),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1175),
.B(n_1116),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1139),
.B(n_1125),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1139),
.B(n_1074),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1165),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1173),
.B(n_1164),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1158),
.B(n_1122),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1169),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1153),
.B(n_1185),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1169),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1147),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1154),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1182),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1188),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1156),
.A2(n_1107),
.B1(n_1119),
.B2(n_1130),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1179),
.Y(n_1231)
);

NOR2x1_ASAP7_75t_L g1232 ( 
.A(n_1156),
.B(n_1121),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1179),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1186),
.A2(n_1125),
.B1(n_1130),
.B2(n_1133),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1154),
.B(n_1090),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1135),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1191),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1168),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1198),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1226),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1197),
.B(n_1088),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1197),
.B(n_1105),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1195),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1216),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1200),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1208),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1219),
.B(n_1090),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1209),
.B(n_1142),
.C(n_1176),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1199),
.Y(n_1249)
);

OAI222xp33_ASAP7_75t_L g1250 ( 
.A1(n_1230),
.A2(n_1183),
.B1(n_1178),
.B2(n_1167),
.C1(n_1172),
.C2(n_1105),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1204),
.B(n_1079),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1203),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1205),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1207),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1221),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1202),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1206),
.B(n_1121),
.Y(n_1257)
);

AOI211xp5_ASAP7_75t_L g1258 ( 
.A1(n_1230),
.A2(n_1174),
.B(n_1171),
.C(n_1159),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1194),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1237),
.B(n_1113),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1212),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1220),
.B(n_1184),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1201),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1218),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1213),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1218),
.B(n_1113),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1228),
.B(n_1136),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1194),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1214),
.B(n_1120),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1244),
.B(n_1217),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1245),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1239),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1268),
.B(n_1193),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1245),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1252),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1259),
.B(n_1193),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1255),
.B(n_1236),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1264),
.B(n_1211),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1246),
.B(n_1215),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1255),
.B(n_1236),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1263),
.B(n_1210),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1252),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1253),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1266),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1253),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1263),
.B(n_1234),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1254),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1266),
.B(n_1234),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1254),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1259),
.B(n_1214),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1272),
.B(n_1243),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1272),
.B(n_1287),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1289),
.A2(n_1248),
.B1(n_1258),
.B2(n_1162),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1277),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1270),
.B(n_1290),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1270),
.B(n_1262),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1290),
.B(n_1260),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1271),
.B(n_1260),
.Y(n_1299)
);

AO221x2_ASAP7_75t_L g1300 ( 
.A1(n_1274),
.A2(n_1250),
.B1(n_1267),
.B2(n_1240),
.C(n_1146),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1279),
.B(n_1251),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1284),
.A2(n_1157),
.B1(n_1231),
.B2(n_1233),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1280),
.B(n_1261),
.Y(n_1303)
);

AOI222xp33_ASAP7_75t_L g1304 ( 
.A1(n_1300),
.A2(n_1247),
.B1(n_1196),
.B2(n_1222),
.C1(n_1284),
.C2(n_1256),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1294),
.A2(n_1232),
.B1(n_1229),
.B2(n_1238),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1295),
.B(n_1240),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1303),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1296),
.B(n_1273),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1293),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1297),
.B(n_1285),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1292),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1301),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1299),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1298),
.B(n_1285),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1302),
.B(n_1275),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1303),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1294),
.A2(n_1273),
.B1(n_1276),
.B2(n_1291),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1293),
.B(n_1286),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1309),
.B(n_1288),
.C(n_1283),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1304),
.A2(n_1247),
.B1(n_1269),
.B2(n_1257),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1309),
.B(n_1282),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1305),
.A2(n_1269),
.B1(n_1257),
.B2(n_1281),
.Y(n_1322)
);

XNOR2xp5_ASAP7_75t_L g1323 ( 
.A(n_1317),
.B(n_1276),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1311),
.B(n_1278),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1306),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1306),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1314),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1315),
.A2(n_1251),
.B(n_1269),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1327),
.B(n_1313),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1326),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1321),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1324),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1325),
.B(n_1316),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1323),
.B(n_1316),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1333),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1329),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1330),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1329),
.Y(n_1338)
);

INVxp33_ASAP7_75t_SL g1339 ( 
.A(n_1334),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1332),
.Y(n_1340)
);

NAND4xp75_ASAP7_75t_L g1341 ( 
.A(n_1340),
.B(n_1331),
.C(n_1320),
.D(n_1328),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1335),
.A2(n_1319),
.B(n_1307),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1336),
.Y(n_1343)
);

AOI211xp5_ASAP7_75t_L g1344 ( 
.A1(n_1338),
.A2(n_1318),
.B(n_1322),
.C(n_1312),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1339),
.A2(n_1337),
.B(n_1308),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1339),
.A2(n_1312),
.B1(n_1305),
.B2(n_1222),
.Y(n_1346)
);

NOR3xp33_ASAP7_75t_L g1347 ( 
.A(n_1337),
.B(n_1170),
.C(n_1310),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1345),
.B(n_1308),
.Y(n_1348)
);

OAI211xp5_ASAP7_75t_L g1349 ( 
.A1(n_1342),
.A2(n_1180),
.B(n_1187),
.C(n_1082),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1341),
.A2(n_1224),
.B1(n_1227),
.B2(n_1265),
.Y(n_1350)
);

OAI211xp5_ASAP7_75t_L g1351 ( 
.A1(n_1343),
.A2(n_1082),
.B(n_1227),
.C(n_1133),
.Y(n_1351)
);

AOI32xp33_ASAP7_75t_L g1352 ( 
.A1(n_1344),
.A2(n_1223),
.A3(n_1225),
.B1(n_1095),
.B2(n_1265),
.Y(n_1352)
);

OAI211xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1347),
.A2(n_1131),
.B(n_1086),
.C(n_1117),
.Y(n_1353)
);

XNOR2xp5_ASAP7_75t_L g1354 ( 
.A(n_1348),
.B(n_1346),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1350),
.B(n_1227),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1353),
.Y(n_1356)
);

XNOR2x1_ASAP7_75t_L g1357 ( 
.A(n_1349),
.B(n_1101),
.Y(n_1357)
);

NOR2x1_ASAP7_75t_L g1358 ( 
.A(n_1351),
.B(n_1131),
.Y(n_1358)
);

NAND2xp33_ASAP7_75t_SL g1359 ( 
.A(n_1354),
.B(n_1352),
.Y(n_1359)
);

NAND2xp33_ASAP7_75t_SL g1360 ( 
.A(n_1357),
.B(n_1117),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_R g1361 ( 
.A(n_1356),
.B(n_275),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_R g1362 ( 
.A(n_1355),
.B(n_276),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_R g1363 ( 
.A(n_1358),
.B(n_278),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1359),
.Y(n_1364)
);

OAI211xp5_ASAP7_75t_L g1365 ( 
.A1(n_1362),
.A2(n_1095),
.B(n_1101),
.C(n_1133),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1361),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1363),
.A2(n_1196),
.B(n_1086),
.Y(n_1367)
);

OAI221xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1366),
.A2(n_1360),
.B1(n_1128),
.B2(n_1249),
.C(n_1120),
.Y(n_1368)
);

AND2x2_ASAP7_75t_SL g1369 ( 
.A(n_1366),
.B(n_1242),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1364),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1370),
.B(n_1367),
.Y(n_1371)
);

XOR2x2_ASAP7_75t_L g1372 ( 
.A(n_1369),
.B(n_1365),
.Y(n_1372)
);

AOI31xp33_ASAP7_75t_L g1373 ( 
.A1(n_1371),
.A2(n_1368),
.A3(n_283),
.B(n_284),
.Y(n_1373)
);

AOI31xp33_ASAP7_75t_L g1374 ( 
.A1(n_1372),
.A2(n_280),
.A3(n_285),
.B(n_289),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1374),
.A2(n_1249),
.B1(n_1242),
.B2(n_1241),
.Y(n_1375)
);

OAI322xp33_ASAP7_75t_L g1376 ( 
.A1(n_1373),
.A2(n_1128),
.A3(n_1083),
.B1(n_1080),
.B2(n_1079),
.C1(n_300),
.C2(n_301),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1376),
.A2(n_1242),
.B(n_1241),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1375),
.A2(n_1241),
.B1(n_1083),
.B2(n_1080),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1376),
.A2(n_1235),
.B1(n_295),
.B2(n_297),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1379),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1380),
.A2(n_1377),
.B1(n_1378),
.B2(n_1235),
.C(n_303),
.Y(n_1381)
);

AOI211xp5_ASAP7_75t_L g1382 ( 
.A1(n_1381),
.A2(n_294),
.B(n_299),
.C(n_302),
.Y(n_1382)
);


endmodule