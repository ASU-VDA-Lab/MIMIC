module fake_jpeg_8916_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_29),
.B1(n_21),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_54),
.B1(n_55),
.B2(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_60),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_42),
.B1(n_41),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_34),
.B1(n_39),
.B2(n_26),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_17),
.B1(n_23),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_17),
.B1(n_23),
.B2(n_26),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_1),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_1),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_16),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_64),
.Y(n_91)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_1),
.Y(n_109)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_74),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_38),
.B1(n_34),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_61),
.B1(n_49),
.B2(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_69),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_39),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_31),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_36),
.C(n_34),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_36),
.C(n_43),
.Y(n_113)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_80),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_74),
.B1(n_86),
.B2(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_99),
.B1(n_100),
.B2(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_57),
.B1(n_52),
.B2(n_56),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_66),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_79),
.B(n_20),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_52),
.C(n_45),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_78),
.C(n_65),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_118),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_84),
.B(n_67),
.C(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_130),
.B1(n_107),
.B2(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_75),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_75),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_121),
.C(n_93),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_135),
.B(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_126),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.C(n_8),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_76),
.B1(n_81),
.B2(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_27),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_134),
.B1(n_95),
.B2(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_145),
.B1(n_115),
.B2(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_144),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_149),
.C(n_152),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_106),
.B1(n_99),
.B2(n_93),
.C(n_97),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_111),
.B1(n_20),
.B2(n_7),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_103),
.C(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_43),
.C(n_33),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_121),
.C(n_119),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_120),
.C(n_122),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_150),
.C(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_139),
.C(n_120),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.C(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_147),
.C(n_137),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_24),
.B1(n_43),
.B2(n_7),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_122),
.C(n_118),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_141),
.C(n_144),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_177),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_176),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_164),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_146),
.B(n_135),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_178),
.B(n_5),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_117),
.A3(n_135),
.B1(n_32),
.B2(n_24),
.C1(n_43),
.C2(n_14),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_43),
.C(n_32),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_182),
.B(n_183),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_9),
.B(n_10),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_15),
.B1(n_11),
.B2(n_7),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_5),
.B(n_6),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_5),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_8),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_170),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_177),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_170),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_186),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_193),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_169),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_196),
.B(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_181),
.C(n_183),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_10),
.B(n_197),
.C(n_198),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_201),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_202),
.Y(n_205)
);


endmodule