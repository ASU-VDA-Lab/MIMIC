module real_jpeg_18655_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g83 ( 
.A(n_0),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_0),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_0),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_0),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_0),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_0),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_2),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_2),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_3),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_3),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_4),
.B(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_5),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_62),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g87 ( 
.A(n_6),
.B(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_6),
.B(n_98),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_6),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_134),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_7),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_8),
.B(n_81),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_8),
.B(n_42),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_8),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_8),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_9),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_9),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_9),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_9),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_9),
.B(n_160),
.Y(n_326)
);

BUFx2_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

NAND2x1_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_10),
.B(n_69),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_10),
.B(n_84),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_10),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_12),
.A2(n_15),
.B1(n_42),
.B2(n_46),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_12),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_12),
.B(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_12),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_14),
.Y(n_119)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_15),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_15),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_15),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_15),
.B(n_79),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_15),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_15),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_15),
.B(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_16),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_212),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_210),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_171),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_20),
.B(n_171),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.C(n_136),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_22),
.A2(n_23),
.B1(n_92),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_65),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_24),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.C(n_51),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_25),
.B(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_33),
.C(n_36),
.Y(n_75)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_35),
.Y(n_353)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_39),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_40),
.A2(n_41),
.B1(n_51),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_41),
.A2(n_232),
.B(n_236),
.Y(n_231)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_51),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.C(n_61),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_52),
.A2(n_53),
.B1(n_61),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_52),
.A2(n_53),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_57),
.B(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_64),
.Y(n_222)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_76),
.B1(n_90),
.B2(n_91),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_66),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_75),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_68),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_68),
.B(n_219),
.C(n_225),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_68),
.A2(n_200),
.B1(n_225),
.B2(n_226),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_70),
.Y(n_235)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_70),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_71),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_75),
.B(n_199),
.C(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_76),
.B(n_91),
.C(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.C(n_88),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_77),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.C(n_83),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_78),
.A2(n_83),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_78),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_78),
.B(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_80),
.B(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_83),
.Y(n_244)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_85),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_92),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_125),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_109),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_94),
.B(n_109),
.C(n_126),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.C(n_105),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_100),
.A2(n_105),
.B1(n_106),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_105),
.B(n_252),
.C(n_255),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_105),
.A2(n_106),
.B1(n_252),
.B2(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_107),
.Y(n_282)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_111),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_111),
.A2(n_120),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_116),
.C(n_121),
.Y(n_184)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_119),
.Y(n_292)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_129),
.C(n_133),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_137),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_164),
.C(n_168),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_138),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_153),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_140),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_143),
.B(n_153),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_144),
.B(n_150),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_154),
.A2(n_158),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_158),
.B(n_323),
.C(n_325),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_158),
.A2(n_249),
.B1(n_325),
.B2(n_326),
.Y(n_336)
);

XOR2x1_ASAP7_75t_L g246 ( 
.A(n_159),
.B(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_165),
.B(n_168),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_195),
.B1(n_208),
.B2(n_209),
.Y(n_174)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_179),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_377),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_268),
.C(n_273),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_260),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_216),
.B(n_260),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_245),
.C(n_258),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_217),
.B(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_230),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_218),
.B(n_231),
.C(n_241),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_219),
.B(n_367),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_SL g312 ( 
.A(n_220),
.B(n_223),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_220),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_220),
.A2(n_330),
.B1(n_331),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_243),
.B(n_280),
.C(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_245),
.B(n_258),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.C(n_256),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_246),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_251),
.B(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2x2_ASAP7_75t_SL g306 ( 
.A(n_255),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_263),
.C(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_269),
.Y(n_379)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_270),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_372),
.B(n_376),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_358),
.B(n_371),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_317),
.B(n_357),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_303),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_277),
.B(n_303),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.C(n_294),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_288),
.B1(n_294),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_289),
.B(n_293),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

AO22x1_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_302),
.B(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_306),
.C(n_309),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_327),
.B(n_356),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_322),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_323),
.A2(n_324),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_337),
.B(n_355),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_334),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_334),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_349),
.B(n_354),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_347),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_346),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_346),
.B(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_370),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_370),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_363),
.B2(n_364),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_365),
.C(n_369),
.Y(n_373)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_368),
.B2(n_369),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_374),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.C(n_380),
.Y(n_377)
);


endmodule