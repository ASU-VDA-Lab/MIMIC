module fake_ariane_2789_n_1109 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1109);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1109;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_244;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_940;
wire n_756;
wire n_466;
wire n_1016;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_222;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_254;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_246;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_258;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_211;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_SL g192 ( 
.A(n_146),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_6),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_91),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_86),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_17),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_96),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_9),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_84),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_76),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_116),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_178),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_81),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_129),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_19),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_180),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_11),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_34),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_14),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_176),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_181),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_55),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_78),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_23),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_18),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_64),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_65),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_121),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_92),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_5),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_18),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_24),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_105),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_111),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_45),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_70),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_97),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_173),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_82),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_15),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_72),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_123),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_134),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_29),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_107),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_61),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_102),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_191),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_19),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_184),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_32),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_220),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_242),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_193),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_201),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_215),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_219),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_248),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_231),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_197),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_239),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_240),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_216),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_253),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_192),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_275),
.A2(n_247),
.B1(n_264),
.B2(n_262),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_243),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_272),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_223),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_265),
.B(n_238),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_282),
.B(n_238),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_267),
.B(n_243),
.C(n_195),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_208),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_268),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_270),
.B(n_194),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_286),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

CKINVDCx6p67_ASAP7_75t_R g348 ( 
.A(n_279),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_196),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_298),
.B(n_198),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_200),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_203),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_287),
.A2(n_294),
.B1(n_271),
.B2(n_274),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_204),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_300),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_291),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_277),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_305),
.B(n_205),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_281),
.B(n_206),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_296),
.B(n_209),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_296),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_297),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_299),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_321),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_299),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_354),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_316),
.B(n_302),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_319),
.A2(n_301),
.B1(n_303),
.B2(n_295),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_322),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_295),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_302),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_304),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_346),
.A2(n_303),
.B1(n_301),
.B2(n_304),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_319),
.A2(n_280),
.B1(n_269),
.B2(n_312),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_367),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_312),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_354),
.B(n_306),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

BUFx6f_ASAP7_75t_SL g430 ( 
.A(n_346),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_318),
.B(n_280),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_340),
.A2(n_310),
.B1(n_309),
.B2(n_307),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_369),
.B(n_306),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_307),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_332),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_332),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_371),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_373),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_396),
.Y(n_449)
);

AO221x1_ASAP7_75t_L g450 ( 
.A1(n_399),
.A2(n_355),
.B1(n_309),
.B2(n_310),
.C(n_371),
.Y(n_450)
);

AO221x1_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_355),
.B1(n_371),
.B2(n_332),
.C(n_368),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_403),
.B(n_340),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_394),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_393),
.B(n_403),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_375),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_393),
.A2(n_369),
.B1(n_340),
.B2(n_349),
.Y(n_462)
);

AO221x1_ASAP7_75t_L g463 ( 
.A1(n_415),
.A2(n_342),
.B1(n_360),
.B2(n_368),
.C(n_338),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_394),
.B(n_343),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_369),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_362),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_403),
.B(n_344),
.Y(n_468)
);

AND2x6_ASAP7_75t_SL g469 ( 
.A(n_392),
.B(n_314),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_357),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_317),
.Y(n_472)
);

BUFx6f_ASAP7_75t_SL g473 ( 
.A(n_393),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

NOR3xp33_ASAP7_75t_L g476 ( 
.A(n_417),
.B(n_366),
.C(n_364),
.Y(n_476)
);

NOR3xp33_ASAP7_75t_L g477 ( 
.A(n_417),
.B(n_333),
.C(n_338),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_L g479 ( 
.A(n_392),
.B(n_345),
.C(n_342),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_418),
.B(n_317),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_393),
.B(n_317),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_377),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_377),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_413),
.B(n_317),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_372),
.B(n_345),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_376),
.B(n_356),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_435),
.B(n_320),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_386),
.B(n_339),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_408),
.B(n_339),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_424),
.B(n_356),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_441),
.B(n_360),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_426),
.B(n_363),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_428),
.B(n_363),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_380),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_426),
.B(n_365),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_383),
.B(n_365),
.C(n_347),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_426),
.B(n_384),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_430),
.B(n_326),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_437),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_384),
.Y(n_508)
);

BUFx6f_ASAP7_75t_SL g509 ( 
.A(n_430),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_430),
.B(n_337),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_383),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_437),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_437),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_426),
.B(n_337),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_384),
.B(n_347),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_442),
.B(n_352),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_432),
.B(n_352),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_385),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_384),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_442),
.B(n_358),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_442),
.B(n_358),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_384),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_387),
.B(n_320),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_384),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_409),
.B(n_361),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_443),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_455),
.B(n_320),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_511),
.A2(n_348),
.B1(n_320),
.B2(n_387),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_457),
.Y(n_534)
);

AO22x2_ASAP7_75t_L g535 ( 
.A1(n_451),
.A2(n_348),
.B1(n_315),
.B2(n_314),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_448),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_450),
.A2(n_315),
.B1(n_427),
.B2(n_425),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_449),
.A2(n_432),
.B1(n_427),
.B2(n_425),
.Y(n_540)
);

BUFx8_ASAP7_75t_L g541 ( 
.A(n_509),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_464),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

AO22x2_ASAP7_75t_L g544 ( 
.A1(n_474),
.A2(n_436),
.B1(n_438),
.B2(n_434),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_449),
.B(n_443),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_453),
.B(n_467),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_459),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_466),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_470),
.A2(n_436),
.B1(n_438),
.B2(n_434),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_452),
.B(n_361),
.Y(n_551)
);

AO22x2_ASAP7_75t_L g552 ( 
.A1(n_463),
.A2(n_439),
.B1(n_444),
.B2(n_440),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_455),
.A2(n_432),
.B1(n_440),
.B2(n_439),
.Y(n_554)
);

AO22x2_ASAP7_75t_L g555 ( 
.A1(n_465),
.A2(n_444),
.B1(n_446),
.B2(n_445),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_493),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_492),
.B(n_388),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_468),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_483),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_370),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_530),
.B(n_388),
.Y(n_561)
);

NAND2x1p5_ASAP7_75t_L g562 ( 
.A(n_526),
.B(n_388),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_492),
.B(n_370),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_486),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

AO22x2_ASAP7_75t_L g566 ( 
.A1(n_479),
.A2(n_446),
.B1(n_445),
.B2(n_402),
.Y(n_566)
);

OAI221xp5_ASAP7_75t_L g567 ( 
.A1(n_477),
.A2(n_405),
.B1(n_422),
.B2(n_421),
.C(n_406),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_488),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_512),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_526),
.B(n_388),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_475),
.B(n_390),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_519),
.A2(n_402),
.B1(n_405),
.B2(n_400),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_520),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_509),
.Y(n_574)
);

OAI221xp5_ASAP7_75t_L g575 ( 
.A1(n_462),
.A2(n_407),
.B1(n_422),
.B2(n_421),
.C(n_400),
.Y(n_575)
);

OR2x2_ASAP7_75t_SL g576 ( 
.A(n_469),
.B(n_378),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_457),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_461),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_492),
.A2(n_407),
.B1(n_406),
.B2(n_379),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_476),
.B(n_390),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_484),
.B(n_390),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_490),
.B(n_390),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_484),
.B(n_419),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_475),
.B(n_423),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_461),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_478),
.Y(n_586)
);

AO22x2_ASAP7_75t_L g587 ( 
.A1(n_478),
.A2(n_379),
.B1(n_381),
.B2(n_378),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_491),
.B(n_419),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_495),
.B(n_419),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g590 ( 
.A1(n_496),
.A2(n_419),
.B1(n_420),
.B2(n_423),
.C(n_416),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_488),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_510),
.B(n_409),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

AO32x2_ASAP7_75t_L g595 ( 
.A1(n_550),
.A2(n_503),
.A3(n_518),
.B1(n_487),
.B2(n_473),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_SL g596 ( 
.A1(n_548),
.A2(n_497),
.B(n_500),
.C(n_504),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_556),
.A2(n_485),
.B1(n_480),
.B2(n_472),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_558),
.A2(n_524),
.B(n_504),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_584),
.Y(n_600)
);

NOR2xp67_ASAP7_75t_L g601 ( 
.A(n_561),
.B(n_510),
.Y(n_601)
);

A2O1A1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_560),
.A2(n_485),
.B(n_505),
.C(n_515),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_542),
.B(n_473),
.Y(n_603)
);

AOI21xp33_ASAP7_75t_L g604 ( 
.A1(n_570),
.A2(n_525),
.B(n_515),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_545),
.A2(n_500),
.B(n_497),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_547),
.Y(n_606)
);

AOI21x1_ASAP7_75t_L g607 ( 
.A1(n_550),
.A2(n_529),
.B(n_516),
.Y(n_607)
);

OR2x6_ASAP7_75t_SL g608 ( 
.A(n_541),
.B(n_210),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_536),
.A2(n_481),
.B(n_498),
.C(n_518),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_589),
.A2(n_529),
.B(n_516),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_590),
.A2(n_521),
.B(n_508),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_538),
.A2(n_481),
.B1(n_528),
.B2(n_514),
.Y(n_612)
);

NOR3xp33_ASAP7_75t_L g613 ( 
.A(n_580),
.B(n_505),
.C(n_528),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_539),
.A2(n_513),
.B1(n_471),
.B2(n_454),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_535),
.A2(n_501),
.B1(n_502),
.B2(n_489),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_546),
.B(n_454),
.Y(n_616)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_593),
.A2(n_522),
.B(n_517),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_543),
.A2(n_471),
.B1(n_521),
.B2(n_508),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_575),
.A2(n_502),
.B(n_506),
.C(n_501),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_557),
.B(n_508),
.Y(n_620)
);

AO32x1_ASAP7_75t_L g621 ( 
.A1(n_534),
.A2(n_506),
.A3(n_507),
.B1(n_379),
.B2(n_381),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_582),
.A2(n_521),
.B(n_508),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_532),
.B(n_549),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_532),
.B(n_507),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_535),
.A2(n_523),
.B1(n_331),
.B2(n_381),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_541),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_557),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_553),
.B(n_521),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_574),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g630 ( 
.A1(n_587),
.A2(n_555),
.B(n_552),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_563),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_546),
.B(n_527),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_564),
.B(n_527),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_563),
.B(n_527),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_533),
.A2(n_331),
.B1(n_382),
.B2(n_378),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_588),
.A2(n_527),
.B(n_395),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_534),
.B(n_382),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_533),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_565),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_576),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_551),
.A2(n_395),
.B(n_382),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_592),
.B(n_395),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_569),
.B(n_398),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_592),
.A2(n_404),
.B(n_398),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_573),
.B(n_584),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_562),
.B(n_398),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_587),
.A2(n_555),
.B(n_552),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_581),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_567),
.A2(n_423),
.B(n_410),
.C(n_412),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_577),
.A2(n_410),
.B(n_404),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_578),
.A2(n_410),
.B(n_404),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_585),
.A2(n_420),
.B(n_416),
.C(n_414),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_601),
.B(n_540),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_603),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_638),
.B(n_586),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_599),
.B(n_537),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_627),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_623),
.B(n_537),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_627),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_602),
.A2(n_597),
.B(n_598),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_633),
.B(n_566),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_646),
.B(n_554),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_646),
.B(n_613),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_606),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_644),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_640),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_627),
.B(n_566),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_616),
.B(n_583),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_630),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_639),
.A2(n_544),
.B1(n_572),
.B2(n_568),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_648),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_641),
.A2(n_544),
.B1(n_572),
.B2(n_591),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_607),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_632),
.B(n_594),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_631),
.B(n_579),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_579),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_628),
.Y(n_678)
);

AND3x1_ASAP7_75t_SL g679 ( 
.A(n_608),
.B(n_0),
.C(n_1),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_635),
.B(n_412),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_595),
.B(n_412),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_649),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_595),
.B(n_414),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_643),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_629),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_600),
.B(n_571),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_631),
.B(n_414),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_617),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_634),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_621),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_621),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_621),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_595),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_631),
.B(n_416),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_619),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_615),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_596),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_626),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_647),
.A2(n_331),
.B1(n_409),
.B2(n_420),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_643),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_643),
.Y(n_701)
);

AND2x2_ASAP7_75t_SL g702 ( 
.A(n_636),
.B(n_625),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_620),
.B(n_331),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_643),
.A2(n_331),
.B1(n_409),
.B2(n_263),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_600),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_649),
.B(n_622),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_612),
.B(n_409),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_604),
.B(n_331),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_614),
.A2(n_331),
.B1(n_409),
.B2(n_261),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_645),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_661),
.A2(n_611),
.B(n_618),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_654),
.A2(n_605),
.B(n_697),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_667),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_662),
.B(n_0),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_667),
.B(n_609),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_705),
.B(n_637),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_678),
.Y(n_718)
);

O2A1O1Ixp5_ASAP7_75t_L g719 ( 
.A1(n_697),
.A2(n_610),
.B(n_650),
.C(n_642),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_662),
.B(n_1),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_702),
.A2(n_651),
.B1(n_652),
.B2(n_233),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_689),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_670),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_684),
.A2(n_653),
.B(n_212),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_689),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_655),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_665),
.B(n_2),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_684),
.A2(n_214),
.B(n_211),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_669),
.B(n_2),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_668),
.B(n_53),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_678),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_670),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_695),
.A2(n_221),
.B(n_218),
.Y(n_734)
);

AOI21x1_ASAP7_75t_L g735 ( 
.A1(n_688),
.A2(n_224),
.B(n_222),
.Y(n_735)
);

O2A1O1Ixp5_ASAP7_75t_L g736 ( 
.A1(n_709),
.A2(n_656),
.B(n_695),
.C(n_664),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_710),
.A2(n_227),
.B(n_225),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_705),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_680),
.B(n_3),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_701),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_680),
.B(n_3),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_708),
.A2(n_232),
.B(n_228),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_658),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_657),
.B(n_4),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_657),
.B(n_4),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_675),
.B(n_5),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_668),
.B(n_56),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_SL g748 ( 
.A1(n_700),
.A2(n_244),
.B(n_234),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_685),
.B(n_6),
.Y(n_749)
);

AND2x4_ASAP7_75t_SL g750 ( 
.A(n_655),
.B(n_57),
.Y(n_750)
);

INVx3_ASAP7_75t_SL g751 ( 
.A(n_685),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_701),
.B(n_58),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_681),
.B(n_683),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_701),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_708),
.A2(n_260),
.B(n_249),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_707),
.B(n_59),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_SL g757 ( 
.A1(n_700),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_711),
.A2(n_254),
.B(n_246),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_658),
.B(n_7),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_672),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_672),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_658),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_663),
.A2(n_258),
.B1(n_256),
.B2(n_255),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_658),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_658),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_666),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_660),
.B(n_8),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_660),
.B(n_10),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_660),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_681),
.B(n_10),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_674),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_655),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_711),
.A2(n_62),
.B(n_60),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_693),
.B(n_11),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_683),
.B(n_12),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_715),
.B(n_666),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_715),
.B(n_677),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_714),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_720),
.B(n_677),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_764),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_722),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_725),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_723),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_756),
.B(n_707),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_720),
.B(n_659),
.Y(n_785)
);

NAND2x1_ASAP7_75t_L g786 ( 
.A(n_729),
.B(n_707),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_730),
.B(n_660),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_660),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_766),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_712),
.A2(n_688),
.B(n_702),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_718),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_744),
.B(n_745),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_755),
.A2(n_702),
.B(n_704),
.C(n_693),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_718),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_SL g795 ( 
.A1(n_713),
.A2(n_691),
.B(n_690),
.C(n_692),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_745),
.B(n_706),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_738),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_716),
.A2(n_699),
.B(n_674),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_772),
.B(n_686),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_770),
.B(n_676),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_770),
.B(n_706),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_756),
.B(n_753),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_775),
.B(n_673),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_775),
.B(n_671),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_774),
.B(n_682),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_726),
.B(n_682),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_757),
.A2(n_687),
.B(n_694),
.C(n_703),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_723),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_751),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_756),
.B(n_686),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_760),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_751),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_774),
.B(n_696),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_719),
.A2(n_691),
.B(n_690),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_721),
.A2(n_696),
.B(n_686),
.C(n_703),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_738),
.A2(n_698),
.B1(n_679),
.B2(n_692),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_736),
.B(n_698),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_753),
.B(n_12),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_746),
.B(n_13),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_739),
.B(n_741),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_732),
.B(n_733),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_769),
.B(n_13),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_729),
.B(n_66),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_733),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_743),
.Y(n_825)
);

O2A1O1Ixp5_ASAP7_75t_L g826 ( 
.A1(n_735),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_750),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_827)
);

OA21x2_ASAP7_75t_L g828 ( 
.A1(n_771),
.A2(n_68),
.B(n_67),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_732),
.B(n_20),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_731),
.B(n_21),
.Y(n_830)
);

BUFx4_ASAP7_75t_R g831 ( 
.A(n_743),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_827),
.A2(n_749),
.B1(n_727),
.B2(n_729),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_SL g833 ( 
.A1(n_827),
.A2(n_750),
.B(n_763),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_783),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_803),
.A2(n_731),
.B1(n_747),
.B2(n_734),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_804),
.A2(n_785),
.B1(n_813),
.B2(n_800),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_819),
.A2(n_747),
.B1(n_731),
.B2(n_758),
.Y(n_837)
);

AOI222xp33_ASAP7_75t_L g838 ( 
.A1(n_793),
.A2(n_737),
.B1(n_747),
.B2(n_761),
.C1(n_771),
.C2(n_768),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_793),
.B(n_767),
.C(n_759),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_805),
.B(n_740),
.Y(n_840)
);

BUFx4f_ASAP7_75t_SL g841 ( 
.A(n_809),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_SL g842 ( 
.A1(n_816),
.A2(n_830),
.B(n_817),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_792),
.B(n_740),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_815),
.A2(n_742),
.B1(n_740),
.B2(n_754),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_SL g845 ( 
.A1(n_828),
.A2(n_752),
.B1(n_754),
.B2(n_773),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_790),
.A2(n_757),
.B1(n_717),
.B2(n_754),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_809),
.B(n_764),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_802),
.A2(n_724),
.B1(n_728),
.B2(n_752),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_791),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_817),
.A2(n_735),
.B1(n_752),
.B2(n_762),
.Y(n_850)
);

AOI222xp33_ASAP7_75t_L g851 ( 
.A1(n_820),
.A2(n_773),
.B1(n_765),
.B2(n_762),
.C1(n_764),
.C2(n_25),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_815),
.A2(n_765),
.B1(n_764),
.B2(n_748),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_797),
.A2(n_764),
.B1(n_748),
.B2(n_23),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_802),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_802),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_781),
.B(n_26),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_782),
.B(n_27),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_787),
.B(n_27),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_SL g859 ( 
.A1(n_818),
.A2(n_28),
.B(n_29),
.Y(n_859)
);

AOI222xp33_ASAP7_75t_L g860 ( 
.A1(n_777),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_801),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_L g862 ( 
.A(n_826),
.B(n_34),
.C(n_35),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_787),
.B(n_776),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_828),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_812),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_780),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_808),
.B(n_38),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_811),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_824),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_779),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_828),
.A2(n_810),
.B1(n_784),
.B2(n_796),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_778),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_812),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_810),
.A2(n_784),
.B1(n_799),
.B2(n_788),
.Y(n_874)
);

AOI222xp33_ASAP7_75t_L g875 ( 
.A1(n_829),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.C1(n_46),
.C2(n_47),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_784),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_834),
.B(n_821),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_843),
.B(n_825),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_869),
.B(n_780),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_868),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_868),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_841),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_858),
.Y(n_883)
);

NAND4xp25_ASAP7_75t_L g884 ( 
.A(n_860),
.B(n_822),
.C(n_795),
.D(n_814),
.Y(n_884)
);

CKINVDCx8_ASAP7_75t_R g885 ( 
.A(n_847),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_859),
.A2(n_799),
.B(n_798),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_839),
.B(n_807),
.C(n_789),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_863),
.B(n_840),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_864),
.A2(n_823),
.B(n_806),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_872),
.B(n_780),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_867),
.B(n_780),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_842),
.A2(n_823),
.B(n_795),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_867),
.B(n_786),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_872),
.B(n_810),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_836),
.B(n_823),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_866),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_866),
.B(n_831),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_874),
.B(n_791),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_866),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_871),
.B(n_794),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_856),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_833),
.A2(n_831),
.B(n_794),
.C(n_50),
.Y(n_902)
);

OAI211xp5_ASAP7_75t_L g903 ( 
.A1(n_875),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_903)
);

NAND4xp25_ASAP7_75t_SL g904 ( 
.A(n_838),
.B(n_48),
.C(n_49),
.D(n_51),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_857),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_849),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_832),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_865),
.A2(n_52),
.B1(n_69),
.B2(n_71),
.C(n_73),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_877),
.B(n_849),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_880),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_846),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_880),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_897),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_878),
.B(n_846),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_878),
.B(n_851),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_906),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_879),
.B(n_845),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_879),
.B(n_848),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_881),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_877),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_888),
.B(n_881),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_891),
.B(n_847),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_894),
.B(n_852),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_906),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_899),
.B(n_844),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_905),
.B(n_850),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_893),
.B(n_862),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_905),
.B(n_870),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_897),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_890),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_900),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_910),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_916),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_911),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_913),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_920),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_910),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_912),
.Y(n_938)
);

AND2x6_ASAP7_75t_L g939 ( 
.A(n_911),
.B(n_894),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_915),
.A2(n_886),
.B(n_902),
.C(n_892),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_913),
.B(n_907),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_927),
.B(n_901),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_916),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_926),
.A2(n_916),
.B(n_925),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_931),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_927),
.B(n_901),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_915),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_936),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_941),
.B(n_929),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_945),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_941),
.B(n_929),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_932),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_932),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_947),
.B(n_921),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_935),
.B(n_930),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_942),
.B(n_914),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_935),
.B(n_930),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_946),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_934),
.B(n_917),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_934),
.B(n_917),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_959),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_953),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_953),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_952),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_949),
.B(n_934),
.Y(n_965)
);

NAND4xp25_ASAP7_75t_L g966 ( 
.A(n_949),
.B(n_940),
.C(n_884),
.D(n_873),
.Y(n_966)
);

INVxp33_ASAP7_75t_SL g967 ( 
.A(n_948),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_951),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_962),
.Y(n_969)
);

CKINVDCx14_ASAP7_75t_R g970 ( 
.A(n_968),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_968),
.B(n_951),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_967),
.Y(n_972)
);

NAND4xp75_ASAP7_75t_L g973 ( 
.A(n_961),
.B(n_960),
.C(n_959),
.D(n_908),
.Y(n_973)
);

NAND4xp25_ASAP7_75t_SL g974 ( 
.A(n_961),
.B(n_960),
.C(n_903),
.D(n_956),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_963),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_969),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_972),
.B(n_954),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_975),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_971),
.B(n_954),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_970),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_973),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_975),
.B(n_967),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_974),
.A2(n_966),
.B(n_958),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_972),
.B(n_965),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_972),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_985),
.Y(n_986)
);

AOI222xp33_ASAP7_75t_L g987 ( 
.A1(n_981),
.A2(n_962),
.B1(n_964),
.B2(n_944),
.C1(n_950),
.C2(n_887),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_977),
.Y(n_988)
);

NAND4xp25_ASAP7_75t_L g989 ( 
.A(n_983),
.B(n_965),
.C(n_882),
.D(n_955),
.Y(n_989)
);

XOR2x2_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_928),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_982),
.B(n_876),
.C(n_950),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_979),
.B(n_955),
.Y(n_992)
);

AND2x4_ASAP7_75t_SL g993 ( 
.A(n_978),
.B(n_957),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_980),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_994),
.B(n_984),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_993),
.B(n_988),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_986),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_992),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_990),
.Y(n_999)
);

NOR2x1_ASAP7_75t_L g1000 ( 
.A(n_989),
.B(n_976),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_987),
.B(n_957),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_991),
.B(n_882),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_934),
.Y(n_1003)
);

OAI211xp5_ASAP7_75t_L g1004 ( 
.A1(n_1000),
.A2(n_885),
.B(n_855),
.C(n_854),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_1001),
.A2(n_883),
.B(n_944),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_995),
.A2(n_938),
.B(n_937),
.C(n_945),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_1003),
.B(n_883),
.Y(n_1007)
);

AOI211x1_ASAP7_75t_L g1008 ( 
.A1(n_996),
.A2(n_904),
.B(n_938),
.C(n_937),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_L g1009 ( 
.A(n_997),
.B(n_853),
.C(n_945),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_998),
.B(n_861),
.C(n_905),
.Y(n_1010)
);

OAI211xp5_ASAP7_75t_L g1011 ( 
.A1(n_1002),
.A2(n_885),
.B(n_925),
.C(n_922),
.Y(n_1011)
);

AOI221xp5_ASAP7_75t_L g1012 ( 
.A1(n_999),
.A2(n_905),
.B1(n_931),
.B2(n_928),
.C(n_914),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_1002),
.A2(n_905),
.B(n_918),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1008),
.B(n_939),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_L g1015 ( 
.A(n_1007),
.B(n_922),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_1005),
.A2(n_921),
.B1(n_931),
.B2(n_933),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_1010),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1006),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_1009),
.B(n_939),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_1004),
.A2(n_939),
.B(n_943),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1011),
.B(n_912),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1012),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1008),
.B(n_939),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_1011),
.A2(n_918),
.B(n_911),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1006),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_1018),
.A2(n_939),
.B(n_943),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_L g1028 ( 
.A(n_1017),
.B(n_889),
.C(n_933),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1014),
.A2(n_939),
.B1(n_911),
.B2(n_837),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_L g1030 ( 
.A(n_1026),
.B(n_52),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_L g1031 ( 
.A(n_1023),
.B(n_895),
.C(n_923),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_1022),
.A2(n_919),
.B(n_923),
.C(n_909),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_1024),
.B(n_898),
.C(n_900),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1016),
.A2(n_939),
.B1(n_919),
.B2(n_835),
.Y(n_1034)
);

AOI221xp5_ASAP7_75t_L g1035 ( 
.A1(n_1020),
.A2(n_924),
.B1(n_890),
.B2(n_909),
.C(n_896),
.Y(n_1035)
);

AOI211xp5_ASAP7_75t_L g1036 ( 
.A1(n_1021),
.A2(n_896),
.B(n_924),
.C(n_77),
.Y(n_1036)
);

OAI311xp33_ASAP7_75t_L g1037 ( 
.A1(n_1027),
.A2(n_1025),
.A3(n_1015),
.B1(n_1019),
.C1(n_80),
.Y(n_1037)
);

AOI331xp33_ASAP7_75t_L g1038 ( 
.A1(n_1030),
.A2(n_74),
.A3(n_75),
.B1(n_79),
.B2(n_83),
.B3(n_85),
.C1(n_87),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_1028),
.B(n_88),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_1032),
.B(n_89),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_1031),
.B(n_90),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_1036),
.B(n_93),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_1029),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_94),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_L g1045 ( 
.A(n_1033),
.B(n_1034),
.C(n_98),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1042),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1041),
.Y(n_1047)
);

XNOR2xp5_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_101),
.Y(n_1048)
);

NAND4xp75_ASAP7_75t_L g1049 ( 
.A(n_1040),
.B(n_1039),
.C(n_1044),
.D(n_1037),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1045),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_1038),
.B(n_103),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1041),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1042),
.B(n_104),
.Y(n_1053)
);

NAND4xp75_ASAP7_75t_L g1054 ( 
.A(n_1042),
.B(n_190),
.C(n_108),
.D(n_109),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1038),
.B(n_106),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_1039),
.Y(n_1056)
);

OAI221xp5_ASAP7_75t_L g1057 ( 
.A1(n_1050),
.A2(n_1051),
.B1(n_1055),
.B2(n_1046),
.C(n_1056),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1048),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1053),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_1047),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_SL g1061 ( 
.A1(n_1052),
.A2(n_1049),
.B(n_1054),
.C(n_113),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_1055),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1051),
.B(n_110),
.Y(n_1063)
);

NAND4xp25_ASAP7_75t_L g1064 ( 
.A(n_1050),
.B(n_112),
.C(n_114),
.D(n_115),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1051),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1051),
.B(n_117),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1060),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1059),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1063),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1066),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1058),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1062),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1057),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_1064),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1061),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1060),
.B(n_118),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1065),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1065),
.Y(n_1079)
);

OAI221xp5_ASAP7_75t_L g1080 ( 
.A1(n_1067),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.C(n_128),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_1077),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1068),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1076),
.A2(n_135),
.B(n_137),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_1069),
.B(n_138),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1074),
.B(n_139),
.Y(n_1086)
);

AOI221xp5_ASAP7_75t_L g1087 ( 
.A1(n_1073),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.C(n_144),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1070),
.B(n_145),
.Y(n_1088)
);

NOR2x1p5_ASAP7_75t_L g1089 ( 
.A(n_1083),
.B(n_1072),
.Y(n_1089)
);

OAI211xp5_ASAP7_75t_SL g1090 ( 
.A1(n_1086),
.A2(n_1071),
.B(n_1082),
.C(n_1075),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1088),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_1084),
.B(n_1078),
.C(n_148),
.Y(n_1092)
);

NOR3x2_ASAP7_75t_L g1093 ( 
.A(n_1085),
.B(n_1078),
.C(n_149),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_1080),
.B(n_1081),
.C(n_1087),
.Y(n_1094)
);

NOR2x1p5_ASAP7_75t_L g1095 ( 
.A(n_1083),
.B(n_147),
.Y(n_1095)
);

AOI211xp5_ASAP7_75t_L g1096 ( 
.A1(n_1090),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_SL g1097 ( 
.A1(n_1091),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1089),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_1098)
);

AOI22x1_ASAP7_75t_L g1099 ( 
.A1(n_1096),
.A2(n_1095),
.B1(n_1093),
.B2(n_1092),
.Y(n_1099)
);

AOI211xp5_ASAP7_75t_L g1100 ( 
.A1(n_1099),
.A2(n_1094),
.B(n_1097),
.C(n_1098),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_1100),
.B(n_161),
.C(n_162),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1101),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1101),
.B(n_189),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_1101),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_L g1105 ( 
.A(n_1104),
.B(n_163),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1102),
.A2(n_164),
.B(n_166),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_1103),
.B(n_167),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1106),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.C(n_172),
.Y(n_1108)
);

AOI211xp5_ASAP7_75t_L g1109 ( 
.A1(n_1108),
.A2(n_1107),
.B(n_1105),
.C(n_175),
.Y(n_1109)
);


endmodule