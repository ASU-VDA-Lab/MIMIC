module fake_ariane_1125_n_652 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_652);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_652;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_617;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_93),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_0),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_39),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_1),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_26),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_32),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_0),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_52),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_83),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_53),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_104),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_50),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_8),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_80),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_58),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_15),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_34),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_68),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_10),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_19),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_24),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

BUFx2_ASAP7_75t_SL g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_103),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_18),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_46),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_44),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_12),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_1),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_29),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_47),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_125),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_5),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_61),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_98),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_107),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_123),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_89),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_101),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_65),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_2),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

BUFx8_ASAP7_75t_SL g210 ( 
.A(n_196),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_2),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_3),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_3),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_165),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_196),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_152),
.B(n_4),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_152),
.B(n_154),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_6),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_140),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_150),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_6),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_7),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_9),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_154),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_11),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_194),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_12),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_170),
.B(n_13),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_13),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_139),
.B(n_14),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_143),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_151),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_189),
.B1(n_193),
.B2(n_201),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_155),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_156),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_213),
.A2(n_189),
.B1(n_193),
.B2(n_201),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_153),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_247),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_207),
.B1(n_206),
.B2(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

AO22x2_ASAP7_75t_L g264 ( 
.A1(n_211),
.A2(n_159),
.B1(n_200),
.B2(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_213),
.A2(n_227),
.B1(n_225),
.B2(n_208),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_221),
.A2(n_204),
.B1(n_192),
.B2(n_190),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_244),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

OR2x6_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_157),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_220),
.B(n_250),
.Y(n_271)
);

BUFx6f_ASAP7_75t_SL g272 ( 
.A(n_221),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_211),
.A2(n_188),
.B1(n_184),
.B2(n_181),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_160),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_162),
.Y(n_276)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_221),
.A2(n_180),
.B1(n_178),
.B2(n_173),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_240),
.A2(n_168),
.B1(n_166),
.B2(n_21),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_220),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_210),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_243),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_217),
.B1(n_214),
.B2(n_230),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_23),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_L g290 ( 
.A1(n_224),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_137),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_211),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_292)
);

AO22x2_ASAP7_75t_L g293 ( 
.A1(n_220),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_48),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_209),
.B(n_136),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_209),
.B(n_49),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_253),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_250),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_298)
);

OA22x2_ASAP7_75t_L g299 ( 
.A1(n_237),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_212),
.B(n_135),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_251),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_237),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_212),
.B(n_134),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_210),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_237),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_245),
.B(n_228),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_255),
.B(n_232),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_232),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_245),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_261),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_253),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_218),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_300),
.A2(n_245),
.B(n_228),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_291),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_268),
.B(n_234),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_289),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_260),
.B(n_234),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_253),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g337 ( 
.A(n_266),
.B(n_242),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_215),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_279),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_270),
.B(n_215),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_270),
.B(n_241),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_241),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_256),
.B(n_218),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_264),
.Y(n_348)
);

XNOR2x2_ASAP7_75t_L g349 ( 
.A(n_264),
.B(n_293),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_236),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_262),
.B(n_236),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_304),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_286),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_303),
.B(n_248),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_285),
.B(n_248),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_292),
.B(n_235),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_280),
.B(n_222),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_263),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_261),
.B(n_248),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_283),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_263),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_283),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_261),
.B(n_248),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_258),
.B(n_222),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_311),
.A2(n_252),
.B(n_231),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_235),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_235),
.B1(n_219),
.B2(n_223),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_371),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_322),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_308),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_235),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_311),
.B(n_316),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_223),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_345),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_318),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_333),
.B(n_76),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_326),
.A2(n_231),
.B(n_223),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_231),
.B(n_223),
.Y(n_391)
);

BUFx4f_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_77),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_307),
.B(n_231),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_216),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_320),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_321),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_78),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_323),
.B(n_216),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_321),
.B(n_216),
.Y(n_402)
);

OR2x2_ASAP7_75t_SL g403 ( 
.A(n_358),
.B(n_79),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_324),
.B(n_216),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_346),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_312),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_82),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_313),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_84),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_339),
.B(n_85),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_346),
.B(n_335),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_314),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_86),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_360),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_350),
.B(n_88),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_90),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_351),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_350),
.B(n_353),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_354),
.B(n_91),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_361),
.A2(n_92),
.B(n_95),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_338),
.Y(n_431)
);

BUFx4f_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_351),
.B(n_355),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_381),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_356),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_434),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_432),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_363),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_385),
.B(n_349),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_437),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_398),
.B(n_361),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_405),
.B(n_97),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_424),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_325),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_378),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_392),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g465 ( 
.A1(n_373),
.A2(n_99),
.B(n_100),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_383),
.B(n_435),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_421),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_414),
.B(n_105),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_387),
.B(n_377),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_380),
.B(n_108),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_418),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_377),
.B(n_109),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_427),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_384),
.B(n_113),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_114),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_388),
.B(n_115),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_394),
.B(n_117),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_119),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_120),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_456),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_446),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_475),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_475),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_448),
.Y(n_489)
);

INVx5_ASAP7_75t_SL g490 ( 
.A(n_442),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_456),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

INVx3_ASAP7_75t_SL g500 ( 
.A(n_438),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_443),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_478),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_453),
.A2(n_384),
.B1(n_431),
.B2(n_416),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_478),
.B(n_426),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_473),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_462),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_473),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_502),
.A2(n_481),
.B1(n_478),
.B2(n_433),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_507),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

BUFx2_ASAP7_75t_SL g515 ( 
.A(n_487),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_501),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_503),
.A2(n_453),
.B(n_481),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_492),
.Y(n_520)
);

INVx6_ASAP7_75t_L g521 ( 
.A(n_483),
.Y(n_521)
);

BUFx8_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_505),
.A2(n_481),
.B1(n_433),
.B2(n_457),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_492),
.B(n_445),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_494),
.Y(n_526)
);

BUFx4f_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_500),
.Y(n_528)
);

CKINVDCx11_ASAP7_75t_R g529 ( 
.A(n_500),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_494),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_491),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_505),
.A2(n_461),
.B1(n_449),
.B2(n_454),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_480),
.Y(n_535)
);

INVx11_ASAP7_75t_L g536 ( 
.A(n_483),
.Y(n_536)
);

BUFx4_ASAP7_75t_SL g537 ( 
.A(n_501),
.Y(n_537)
);

CKINVDCx6p67_ASAP7_75t_R g538 ( 
.A(n_483),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_512),
.A2(n_505),
.B1(n_454),
.B2(n_449),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_523),
.A2(n_449),
.B1(n_455),
.B2(n_459),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_533),
.A2(n_449),
.B1(n_455),
.B2(n_459),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_518),
.A2(n_452),
.B1(n_373),
.B2(n_479),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_479),
.B1(n_441),
.B2(n_468),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_519),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_441),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_516),
.A2(n_403),
.B1(n_392),
.B2(n_400),
.Y(n_546)
);

BUFx4f_ASAP7_75t_SL g547 ( 
.A(n_522),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_524),
.A2(n_468),
.B(n_389),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g550 ( 
.A1(n_526),
.A2(n_417),
.B(n_451),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_469),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_515),
.B(n_469),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_530),
.A2(n_389),
.B(n_426),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_531),
.A2(n_430),
.B(n_476),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_532),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_534),
.A2(n_450),
.B1(n_463),
.B2(n_467),
.Y(n_556)
);

CKINVDCx11_ASAP7_75t_R g557 ( 
.A(n_529),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_521),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_521),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_525),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_527),
.A2(n_465),
.B1(n_458),
.B2(n_430),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_417),
.B(n_440),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_477),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_538),
.A2(n_460),
.B1(n_466),
.B2(n_429),
.Y(n_564)
);

OAI222xp33_ASAP7_75t_L g565 ( 
.A1(n_537),
.A2(n_429),
.B1(n_482),
.B2(n_485),
.C1(n_484),
.C2(n_495),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_514),
.A2(n_429),
.B1(n_458),
.B2(n_465),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_536),
.A2(n_486),
.B1(n_489),
.B2(n_497),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_525),
.A2(n_458),
.B1(n_407),
.B2(n_422),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_514),
.A2(n_485),
.B1(n_495),
.B2(n_482),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_546),
.A2(n_410),
.B1(n_444),
.B2(n_519),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_543),
.A2(n_484),
.B1(n_496),
.B2(n_412),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_555),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_517),
.Y(n_573)
);

OAI222xp33_ASAP7_75t_L g574 ( 
.A1(n_543),
.A2(n_496),
.B1(n_413),
.B2(n_474),
.C1(n_472),
.C2(n_471),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_545),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_561),
.A2(n_470),
.B1(n_375),
.B2(n_473),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_542),
.A2(n_375),
.B1(n_447),
.B2(n_410),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_542),
.A2(n_447),
.B1(n_374),
.B2(n_408),
.Y(n_578)
);

NOR3xp33_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_425),
.C(n_413),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_568),
.A2(n_489),
.B1(n_486),
.B2(n_497),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_552),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_566),
.A2(n_447),
.B1(n_374),
.B2(n_408),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_564),
.A2(n_522),
.B1(n_517),
.B2(n_490),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_504),
.C(n_498),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_562),
.B(n_504),
.C(n_498),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_553),
.B(n_504),
.C(n_498),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_566),
.A2(n_444),
.B1(n_471),
.B2(n_401),
.Y(n_587)
);

OAI222xp33_ASAP7_75t_L g588 ( 
.A1(n_539),
.A2(n_376),
.B1(n_404),
.B2(n_386),
.C1(n_499),
.C2(n_506),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_541),
.A2(n_386),
.B1(n_404),
.B2(n_418),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_549),
.A2(n_486),
.B1(n_489),
.B2(n_497),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_544),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_541),
.A2(n_539),
.B1(n_540),
.B2(n_563),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_548),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_581),
.B(n_559),
.Y(n_594)
);

AOI21xp33_ASAP7_75t_SL g595 ( 
.A1(n_591),
.A2(n_547),
.B(n_557),
.Y(n_595)
);

AOI221xp5_ASAP7_75t_L g596 ( 
.A1(n_579),
.A2(n_556),
.B1(n_565),
.B2(n_540),
.C(n_558),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_560),
.Y(n_597)
);

NAND2x1_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_560),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_572),
.B(n_567),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_592),
.A2(n_569),
.B1(n_556),
.B2(n_508),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_506),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_570),
.A2(n_391),
.B(n_390),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_585),
.B(n_584),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_590),
.B(n_576),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_506),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_574),
.A2(n_390),
.B(n_391),
.Y(n_606)
);

NAND4xp25_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_395),
.C(n_402),
.D(n_508),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_597),
.B(n_571),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_596),
.B(n_589),
.C(n_580),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_582),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_593),
.B(n_498),
.Y(n_611)
);

NAND4xp25_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_587),
.C(n_499),
.D(n_402),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_604),
.A2(n_493),
.B1(n_511),
.B2(n_499),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_594),
.Y(n_614)
);

NOR2x1p5_ASAP7_75t_L g615 ( 
.A(n_598),
.B(n_607),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_595),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_614),
.B(n_599),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_606),
.C(n_602),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_608),
.Y(n_619)
);

XOR2x2_ASAP7_75t_L g620 ( 
.A(n_609),
.B(n_605),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_601),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_610),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_619),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_620),
.B(n_612),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_619),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_618),
.A2(n_613),
.B1(n_600),
.B2(n_493),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_616),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_623),
.Y(n_628)
);

OA22x2_ASAP7_75t_L g629 ( 
.A1(n_624),
.A2(n_621),
.B1(n_622),
.B2(n_617),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_626),
.A2(n_618),
.B1(n_627),
.B2(n_625),
.Y(n_630)
);

OA22x2_ASAP7_75t_L g631 ( 
.A1(n_624),
.A2(n_574),
.B1(n_588),
.B2(n_490),
.Y(n_631)
);

XNOR2x1_ASAP7_75t_L g632 ( 
.A(n_624),
.B(n_121),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_628),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_632),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_630),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_634),
.A2(n_631),
.B1(n_629),
.B2(n_493),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_633),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_637),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_638),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_639),
.Y(n_640)
);

AO22x2_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_635),
.B1(n_633),
.B2(n_636),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_641),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_642),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_643),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_490),
.B1(n_511),
.B2(n_493),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_645),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_490),
.B1(n_511),
.B2(n_504),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_646),
.A2(n_511),
.B1(n_504),
.B2(n_498),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_648),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_647),
.Y(n_650)
);

AOI221xp5_ASAP7_75t_L g651 ( 
.A1(n_649),
.A2(n_588),
.B1(n_510),
.B2(n_128),
.C(n_129),
.Y(n_651)
);

AOI211xp5_ASAP7_75t_L g652 ( 
.A1(n_651),
.A2(n_650),
.B(n_510),
.C(n_132),
.Y(n_652)
);


endmodule