module fake_jpeg_425_n_694 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_694);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_694;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_538;
wire n_358;
wire n_47;
wire n_625;
wire n_312;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_10),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_5),
.B(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_60),
.B(n_63),
.Y(n_180)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_62),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_8),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_109),
.Y(n_148)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g166 ( 
.A(n_70),
.Y(n_166)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_74),
.B(n_76),
.Y(n_186)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_75),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_23),
.B(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_85),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_86),
.B(n_87),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_10),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g177 ( 
.A(n_89),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_90),
.B(n_92),
.Y(n_201)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_39),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_91),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_36),
.B(n_6),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_98),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_102),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_103),
.B(n_104),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_6),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_11),
.Y(n_109)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_110),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_118),
.B(n_55),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_19),
.Y(n_119)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_121),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_19),
.Y(n_128)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_23),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_31),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_134),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_55),
.B1(n_35),
.B2(n_56),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_147),
.A2(n_100),
.B1(n_61),
.B2(n_105),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_158),
.A2(n_162),
.B1(n_49),
.B2(n_41),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_71),
.A2(n_55),
.B1(n_34),
.B2(n_54),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_164),
.B(n_165),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_172),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_174),
.B(n_184),
.Y(n_258)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_91),
.B(n_56),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g300 ( 
.A(n_185),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_96),
.A2(n_56),
.B1(n_57),
.B2(n_35),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_188),
.A2(n_224),
.B(n_0),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_192),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_194),
.B(n_210),
.Y(n_267)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_67),
.Y(n_210)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_108),
.Y(n_213)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_77),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_5),
.Y(n_276)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_26),
.Y(n_230)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_106),
.Y(n_223)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

HAxp5_ASAP7_75t_SL g224 ( 
.A(n_74),
.B(n_57),
.CON(n_224),
.SN(n_224)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_79),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_230),
.B(n_237),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g236 ( 
.A1(n_186),
.A2(n_93),
.A3(n_85),
.B1(n_113),
.B2(n_131),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_236),
.B(n_239),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_54),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_94),
.B1(n_81),
.B2(n_111),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_240),
.A2(n_275),
.B1(n_281),
.B2(n_295),
.Y(n_328)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

INVx3_ASAP7_75t_SL g352 ( 
.A(n_241),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_157),
.A2(n_57),
.B1(n_128),
.B2(n_119),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_242),
.A2(n_261),
.B1(n_170),
.B2(n_151),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_41),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_243),
.B(n_245),
.Y(n_347)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx4_ASAP7_75t_SL g340 ( 
.A(n_244),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_148),
.B(n_32),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_32),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_247),
.B(n_248),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_175),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_180),
.B(n_30),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_250),
.B(n_251),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_171),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_139),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_186),
.A2(n_95),
.B1(n_97),
.B2(n_99),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_253),
.A2(n_265),
.B1(n_297),
.B2(n_259),
.Y(n_309)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_254),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_132),
.Y(n_255)
);

INVx11_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_180),
.B(n_49),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_256),
.B(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_257),
.Y(n_345)
);

OA22x2_ASAP7_75t_L g335 ( 
.A1(n_259),
.A2(n_163),
.B1(n_203),
.B2(n_198),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_168),
.A2(n_57),
.B1(n_110),
.B2(n_88),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_195),
.B(n_14),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_264),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_192),
.A2(n_64),
.B1(n_85),
.B2(n_125),
.Y(n_265)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_176),
.Y(n_270)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_270),
.Y(n_351)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_271),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_147),
.A2(n_38),
.B1(n_46),
.B2(n_12),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_272),
.Y(n_332)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_146),
.Y(n_274)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_195),
.A2(n_38),
.B1(n_12),
.B2(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_276),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

CKINVDCx12_ASAP7_75t_R g279 ( 
.A(n_166),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_171),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_289),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_188),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_281)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_137),
.Y(n_285)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_184),
.A2(n_13),
.B(n_15),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_286),
.Y(n_366)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_144),
.B(n_183),
.Y(n_289)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_190),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_140),
.B(n_4),
.C(n_14),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_156),
.C(n_181),
.Y(n_337)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_191),
.A2(n_4),
.B1(n_18),
.B2(n_3),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_181),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_301),
.Y(n_343)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_152),
.B(n_199),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_134),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_302),
.B(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_154),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_138),
.Y(n_304)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_169),
.Y(n_305)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_143),
.B(n_3),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_189),
.Y(n_307)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_309),
.B(n_335),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_258),
.B(n_224),
.CI(n_160),
.CON(n_311),
.SN(n_311)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_153),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_179),
.B1(n_225),
.B2(n_216),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_314),
.A2(n_323),
.B1(n_244),
.B2(n_274),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_173),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_317),
.B(n_360),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_238),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_318),
.B(n_334),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_267),
.A2(n_305),
.B1(n_179),
.B2(n_216),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g329 ( 
.A(n_231),
.B(n_178),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_SL g394 ( 
.A(n_329),
.B(n_249),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_242),
.A2(n_145),
.B1(n_225),
.B2(n_163),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_309),
.B1(n_357),
.B2(n_328),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_268),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_261),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_227),
.B(n_228),
.C(n_235),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_344),
.B(n_367),
.C(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_234),
.Y(n_346)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_346),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_354),
.A2(n_283),
.B1(n_249),
.B2(n_260),
.Y(n_400)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_234),
.Y(n_355)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_232),
.A2(n_145),
.B1(n_167),
.B2(n_203),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_241),
.B1(n_294),
.B2(n_252),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_268),
.B(n_161),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_285),
.A2(n_135),
.B1(n_151),
.B2(n_211),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_290),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_235),
.B(n_166),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_266),
.B(n_159),
.C(n_149),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_266),
.B(n_296),
.C(n_291),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_317),
.B(n_300),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_370),
.B(n_335),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_177),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_372),
.B(n_375),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_292),
.Y(n_375)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_300),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_378),
.B(n_380),
.Y(n_438)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_232),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_381),
.A2(n_330),
.B1(n_319),
.B2(n_356),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_382),
.B(n_387),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_298),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_385),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_299),
.Y(n_385)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g439 ( 
.A(n_386),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_329),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_394),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_417),
.Y(n_426)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_329),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_402),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_393),
.A2(n_415),
.B1(n_418),
.B2(n_352),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_320),
.A2(n_193),
.B1(n_198),
.B2(n_167),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_321),
.B1(n_363),
.B2(n_352),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_288),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_401),
.Y(n_456)
);

O2A1O1Ixp33_ASAP7_75t_L g397 ( 
.A1(n_332),
.A2(n_290),
.B(n_215),
.C(n_233),
.Y(n_397)
);

AO21x1_ASAP7_75t_L g435 ( 
.A1(n_397),
.A2(n_413),
.B(n_389),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_311),
.B(n_233),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_398),
.A2(n_308),
.B(n_361),
.Y(n_458)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_399),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_345),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_319),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_403),
.Y(n_421)
);

INVx13_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_404),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_320),
.B(n_254),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_406),
.B(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_333),
.B(n_296),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_316),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_414),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_291),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_416),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_366),
.A2(n_260),
.B1(n_136),
.B2(n_282),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_347),
.B(n_282),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_310),
.B(n_277),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_367),
.C(n_364),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_422),
.B(n_432),
.C(n_443),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_381),
.A2(n_366),
.B1(n_335),
.B2(n_311),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_427),
.A2(n_428),
.B1(n_450),
.B2(n_452),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_374),
.B(n_325),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_377),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_433),
.B(n_440),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_442),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_377),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_344),
.C(n_324),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_401),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_420),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_398),
.A2(n_308),
.B(n_361),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g489 ( 
.A1(n_448),
.A2(n_397),
.B(n_385),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_411),
.A2(n_406),
.B1(n_395),
.B2(n_410),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_324),
.C(n_326),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_443),
.C(n_422),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_410),
.A2(n_374),
.B1(n_399),
.B2(n_370),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_410),
.A2(n_335),
.B1(n_331),
.B2(n_321),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_453),
.A2(n_457),
.B1(n_459),
.B2(n_393),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_387),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_388),
.A2(n_348),
.B1(n_356),
.B2(n_313),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_454),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_469),
.Y(n_499)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_462),
.Y(n_506)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_436),
.B(n_414),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_465),
.B(n_485),
.Y(n_503)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_373),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_468),
.B(n_474),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_440),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_473),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_472),
.A2(n_453),
.B1(n_459),
.B2(n_420),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_454),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_378),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_375),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_475),
.B(n_480),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_372),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_481),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_482),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g479 ( 
.A(n_421),
.B(n_322),
.C(n_384),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_479),
.B(n_484),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_380),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_435),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_454),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_486),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_436),
.B(n_416),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_370),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_445),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_425),
.C(n_456),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_423),
.A2(n_370),
.B1(n_398),
.B2(n_389),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_488),
.A2(n_452),
.B1(n_426),
.B2(n_458),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_489),
.A2(n_448),
.B(n_435),
.Y(n_524)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_491),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_382),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_493),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_438),
.B(n_417),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_497),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_438),
.B(n_340),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_496),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_456),
.B(n_327),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_430),
.B(n_372),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_515),
.C(n_519),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_480),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_501),
.B(n_522),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_504),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_425),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_505),
.B(n_507),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_425),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_470),
.A2(n_450),
.B1(n_427),
.B2(n_426),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_470),
.A2(n_426),
.B1(n_428),
.B2(n_447),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_472),
.A2(n_449),
.B1(n_434),
.B2(n_447),
.Y(n_513)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_513),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_485),
.C(n_465),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_469),
.B(n_394),
.C(n_429),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_461),
.B(n_449),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_383),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_491),
.Y(n_522)
);

XNOR2x2_ASAP7_75t_SL g537 ( 
.A(n_524),
.B(n_488),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_460),
.A2(n_429),
.B1(n_442),
.B2(n_431),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_526),
.A2(n_464),
.B1(n_490),
.B2(n_486),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_461),
.B(n_408),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_527),
.B(n_521),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_473),
.A2(n_431),
.B1(n_413),
.B2(n_424),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_528),
.A2(n_463),
.B1(n_402),
.B2(n_412),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_478),
.B(n_407),
.C(n_392),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_494),
.C(n_492),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_371),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_532),
.B(n_533),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_477),
.B(n_371),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_477),
.B(n_482),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_390),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_493),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_535),
.B(n_466),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_483),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_536),
.B(n_543),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_537),
.B(n_540),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_482),
.B(n_478),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_539),
.A2(n_548),
.B(n_511),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_520),
.Y(n_541)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_481),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_455),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_544),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_545),
.A2(n_500),
.B1(n_528),
.B2(n_532),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_499),
.A2(n_476),
.B(n_497),
.Y(n_548)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_549),
.Y(n_586)
);

OA22x2_ASAP7_75t_L g550 ( 
.A1(n_526),
.A2(n_508),
.B1(n_510),
.B2(n_509),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_559),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g581 ( 
.A(n_551),
.B(n_564),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_515),
.B(n_409),
.C(n_392),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_554),
.C(n_562),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_498),
.B(n_424),
.C(n_418),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_555),
.A2(n_557),
.B1(n_561),
.B2(n_530),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_499),
.B(n_379),
.Y(n_556)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_556),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_529),
.A2(n_383),
.B1(n_462),
.B2(n_390),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_558),
.Y(n_577)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_516),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_560),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_326),
.C(n_327),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_519),
.B(n_376),
.C(n_386),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_565),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_397),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_503),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_516),
.Y(n_565)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_512),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_567),
.Y(n_584)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_523),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_568),
.B(n_523),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_505),
.B(n_339),
.C(n_338),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_525),
.C(n_502),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_548),
.A2(n_539),
.B(n_542),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_572),
.B(n_579),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_576),
.A2(n_592),
.B(n_596),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_580),
.B(n_581),
.Y(n_616)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_582),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_583),
.A2(n_587),
.B1(n_560),
.B2(n_534),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_566),
.A2(n_511),
.B1(n_529),
.B2(n_500),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_547),
.B(n_551),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_588),
.B(n_591),
.Y(n_599)
);

CKINVDCx14_ASAP7_75t_R g589 ( 
.A(n_540),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_595),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_553),
.B(n_531),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_546),
.A2(n_531),
.B(n_533),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_554),
.B(n_531),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_594),
.B(n_597),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_546),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_546),
.A2(n_533),
.B(n_532),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_538),
.C(n_562),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_598),
.B(n_600),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_SL g600 ( 
.A(n_593),
.B(n_552),
.C(n_559),
.Y(n_600)
);

A2O1A1O1Ixp25_ASAP7_75t_L g604 ( 
.A1(n_573),
.A2(n_537),
.B(n_534),
.C(n_550),
.D(n_538),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_604),
.B(n_606),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_586),
.A2(n_545),
.B1(n_556),
.B2(n_555),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_605),
.A2(n_587),
.B1(n_583),
.B2(n_577),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_547),
.C(n_569),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_506),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_607),
.B(n_608),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_594),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_597),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_609),
.A2(n_619),
.B1(n_439),
.B2(n_386),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_502),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_611),
.B(n_612),
.Y(n_628)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_582),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_576),
.B(n_550),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_613),
.B(n_617),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_574),
.B(n_557),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_614),
.B(n_580),
.Y(n_624)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_584),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_550),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_618),
.B(n_603),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_574),
.B(n_560),
.C(n_339),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_620),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_588),
.B(n_338),
.C(n_362),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_621),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_622),
.A2(n_630),
.B1(n_404),
.B2(n_193),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_604),
.A2(n_572),
.B(n_573),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g656 ( 
.A1(n_623),
.A2(n_625),
.B(n_358),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_624),
.B(n_637),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_610),
.A2(n_590),
.B(n_592),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_596),
.C(n_581),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_627),
.B(n_633),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_SL g629 ( 
.A(n_616),
.B(n_577),
.Y(n_629)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_629),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_610),
.A2(n_570),
.B1(n_584),
.B2(n_312),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_602),
.A2(n_570),
.B1(n_313),
.B2(n_312),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_635),
.A2(n_621),
.B1(n_616),
.B2(n_353),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_600),
.A2(n_615),
.B1(n_609),
.B2(n_614),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_639),
.B(n_640),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_601),
.B(n_598),
.C(n_606),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_608),
.B(n_177),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_641),
.B(n_599),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_625),
.A2(n_620),
.B(n_599),
.Y(n_644)
);

MAJx2_ASAP7_75t_L g659 ( 
.A(n_644),
.B(n_656),
.C(n_637),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_645),
.Y(n_660)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_647),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_631),
.A2(n_376),
.B(n_439),
.Y(n_648)
);

XNOR2x1_ASAP7_75t_L g661 ( 
.A(n_648),
.B(n_641),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_626),
.A2(n_353),
.B1(n_246),
.B2(n_404),
.Y(n_649)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_649),
.Y(n_663)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_630),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_651),
.B(n_656),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_652),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_638),
.A2(n_155),
.B1(n_161),
.B2(n_255),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_653),
.B(n_654),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_640),
.B(n_362),
.C(n_358),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_628),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_655),
.B(n_350),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_632),
.B(n_351),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_657),
.B(n_636),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_L g679 ( 
.A(n_659),
.B(n_661),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_661),
.B(n_644),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_650),
.A2(n_623),
.B(n_629),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_665),
.A2(n_642),
.B(n_646),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_667),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_634),
.C(n_627),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_668),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_655),
.B(n_624),
.Y(n_669)
);

AOI31xp33_ASAP7_75t_L g676 ( 
.A1(n_669),
.A2(n_670),
.A3(n_654),
.B(n_648),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_672),
.B(n_673),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_667),
.B(n_660),
.C(n_651),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_674),
.A2(n_676),
.B(n_677),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_662),
.A2(n_642),
.B(n_646),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_663),
.B(n_652),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_678),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_679),
.B(n_653),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_675),
.B(n_658),
.C(n_664),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_680),
.B(n_683),
.C(n_671),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_671),
.A2(n_658),
.B(n_659),
.Y(n_683)
);

XOR2xp5_ASAP7_75t_L g686 ( 
.A(n_685),
.B(n_679),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_686),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_SL g689 ( 
.A1(n_687),
.A2(n_688),
.B1(n_277),
.B2(n_262),
.Y(n_689)
);

AOI322xp5_ASAP7_75t_L g688 ( 
.A1(n_681),
.A2(n_673),
.A3(n_255),
.B1(n_155),
.B2(n_172),
.C1(n_222),
.C2(n_262),
.Y(n_688)
);

AOI322xp5_ASAP7_75t_L g691 ( 
.A1(n_689),
.A2(n_682),
.A3(n_684),
.B1(n_686),
.B2(n_350),
.C1(n_351),
.C2(n_3),
.Y(n_691)
);

OAI21xp33_ASAP7_75t_SL g692 ( 
.A1(n_691),
.A2(n_690),
.B(n_2),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_692),
.A2(n_1),
.B(n_3),
.C(n_431),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_693),
.A2(n_1),
.B(n_431),
.Y(n_694)
);


endmodule