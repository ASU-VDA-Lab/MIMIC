module fake_jpeg_14308_n_595 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_595);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_595;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_59),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_71),
.Y(n_130)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_68),
.B(n_78),
.Y(n_167)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_76),
.B(n_82),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_21),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_102),
.Y(n_147)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_88),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_93),
.B(n_106),
.Y(n_175)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_25),
.Y(n_103)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_17),
.B(n_1),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_30),
.Y(n_108)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_116),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_56),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_121),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g121 ( 
.A(n_56),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_30),
.B1(n_45),
.B2(n_42),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_126),
.A2(n_140),
.B1(n_160),
.B2(n_186),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_132),
.B(n_137),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_45),
.B1(n_42),
.B2(n_34),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_55),
.B(n_49),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_144),
.B(n_180),
.C(n_46),
.Y(n_238)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_108),
.A2(n_45),
.B1(n_34),
.B2(n_54),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_58),
.B(n_27),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_164),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_75),
.B(n_27),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_21),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_182),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_32),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_173),
.B(n_178),
.Y(n_246)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_57),
.Y(n_176)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_79),
.B(n_32),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_66),
.A2(n_34),
.B(n_3),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_81),
.A2(n_55),
.B1(n_49),
.B2(n_48),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_36),
.B1(n_47),
.B2(n_44),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_53),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_61),
.A2(n_44),
.B1(n_48),
.B2(n_47),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_105),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_191),
.B(n_99),
.Y(n_251)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_62),
.Y(n_197)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_19),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_200),
.B(n_204),
.Y(n_292)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_202),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_203),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_123),
.A2(n_74),
.B1(n_104),
.B2(n_101),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_207),
.A2(n_198),
.B1(n_196),
.B2(n_185),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_208),
.Y(n_319)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_209),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_114),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_210),
.B(n_214),
.Y(n_297)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_133),
.Y(n_211)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_111),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_215),
.B(n_221),
.Y(n_306)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_217),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_142),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_156),
.B(n_53),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_147),
.B(n_111),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_222),
.B(n_230),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_138),
.A2(n_67),
.B1(n_69),
.B2(n_59),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_223),
.A2(n_252),
.B1(n_261),
.B2(n_262),
.Y(n_273)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_225),
.A2(n_238),
.B1(n_265),
.B2(n_267),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_66),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_226),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_134),
.B(n_63),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_227),
.B(n_159),
.C(n_127),
.Y(n_304)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_229),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_145),
.B(n_36),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_135),
.A2(n_91),
.B1(n_89),
.B2(n_85),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_234),
.A2(n_196),
.B1(n_169),
.B2(n_185),
.Y(n_294)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_37),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_243),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_37),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_237),
.B(n_242),
.Y(n_322)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_239),
.Y(n_326)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_240),
.Y(n_276)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_151),
.Y(n_241)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_171),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_244),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_128),
.B(n_46),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_249),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_184),
.B(n_79),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_97),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_128),
.B(n_39),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_136),
.B(n_39),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_251),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_138),
.A2(n_86),
.B1(n_77),
.B2(n_80),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_189),
.B(n_2),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_253),
.B(n_255),
.Y(n_321)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_254),
.Y(n_311)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_186),
.B(n_3),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_269),
.Y(n_312)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_158),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_155),
.B(n_3),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_260),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_127),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_263),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_160),
.A2(n_4),
.B(n_5),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_122),
.B(n_8),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_162),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_155),
.B(n_6),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_162),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_268),
.Y(n_323)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_153),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_219),
.A2(n_176),
.B1(n_197),
.B2(n_83),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g367 ( 
.A1(n_282),
.A2(n_288),
.B1(n_308),
.B2(n_314),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_236),
.A2(n_166),
.B1(n_148),
.B2(n_198),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_263),
.B1(n_259),
.B2(n_205),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_238),
.B(n_127),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_206),
.B(n_159),
.Y(n_286)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_212),
.A2(n_140),
.B(n_126),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_293),
.A2(n_229),
.B1(n_258),
.B2(n_224),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_294),
.A2(n_213),
.B1(n_208),
.B2(n_203),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_227),
.B(n_142),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_296),
.B(n_298),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_227),
.B(n_141),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_304),
.B(n_152),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_219),
.A2(n_188),
.B(n_122),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_207),
.A2(n_73),
.B1(n_183),
.B2(n_169),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_246),
.A2(n_152),
.B1(n_150),
.B2(n_124),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_226),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_305),
.C(n_303),
.Y(n_363)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_307),
.A2(n_264),
.B1(n_234),
.B2(n_252),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_328),
.A2(n_331),
.B1(n_338),
.B2(n_343),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_299),
.B(n_220),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_329),
.B(n_333),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_330),
.B(n_344),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_307),
.A2(n_223),
.B1(n_183),
.B2(n_202),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_332),
.A2(n_309),
.B(n_311),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_244),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_362),
.B1(n_320),
.B2(n_295),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_211),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_339),
.B(n_347),
.Y(n_404)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_340),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_199),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_342),
.B(n_345),
.Y(n_374)
);

OAI22x1_ASAP7_75t_SL g343 ( 
.A1(n_273),
.A2(n_257),
.B1(n_269),
.B2(n_261),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_322),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_349),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_254),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_348),
.A2(n_368),
.B1(n_281),
.B2(n_280),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_241),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_232),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_232),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_355),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_369),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_288),
.A2(n_216),
.B1(n_205),
.B2(n_267),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_354),
.A2(n_358),
.B1(n_294),
.B2(n_295),
.Y(n_384)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_360),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_231),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_357),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_316),
.A2(n_216),
.B1(n_265),
.B2(n_262),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_286),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_364),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_363),
.A2(n_284),
.B(n_315),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_7),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_7),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_366),
.Y(n_406)
);

AO22x1_ASAP7_75t_SL g366 ( 
.A1(n_286),
.A2(n_152),
.B1(n_150),
.B2(n_124),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_286),
.B(n_7),
.Y(n_369)
);

OAI31xp33_ASAP7_75t_L g370 ( 
.A1(n_361),
.A2(n_336),
.A3(n_367),
.B(n_366),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_370),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_372),
.B(n_345),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_332),
.A2(n_308),
.B(n_367),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_373),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_284),
.C(n_298),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_401),
.C(n_402),
.Y(n_431)
);

OAI32xp33_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_275),
.A3(n_290),
.B1(n_310),
.B2(n_301),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_366),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_380),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_SL g383 ( 
.A(n_364),
.B(n_304),
.C(n_296),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g423 ( 
.A(n_383),
.B(n_338),
.CI(n_270),
.CON(n_423),
.SN(n_423)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_384),
.A2(n_397),
.B1(n_405),
.B2(n_335),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_389),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_359),
.A2(n_282),
.B1(n_291),
.B2(n_314),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_399),
.B1(n_343),
.B2(n_406),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_336),
.A2(n_291),
.B(n_287),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_330),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_391),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_340),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_340),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_403),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_328),
.A2(n_282),
.B1(n_287),
.B2(n_275),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_282),
.B1(n_314),
.B2(n_279),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_400),
.B(n_276),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_344),
.C(n_336),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_302),
.C(n_274),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_340),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_331),
.A2(n_314),
.B1(n_300),
.B2(n_285),
.Y(n_405)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_407),
.Y(n_410)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_410),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_411),
.A2(n_432),
.B1(n_386),
.B2(n_399),
.Y(n_452)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_412),
.A2(n_404),
.B(n_380),
.Y(n_464)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_365),
.C(n_369),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_425),
.C(n_427),
.Y(n_446)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_415),
.Y(n_465)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_341),
.Y(n_418)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_358),
.Y(n_419)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_406),
.A2(n_329),
.A3(n_367),
.B1(n_356),
.B2(n_354),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_377),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_376),
.B1(n_384),
.B2(n_405),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_422),
.B(n_424),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_372),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_390),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_368),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_360),
.Y(n_426)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_355),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_398),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_428),
.B(n_379),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_397),
.A2(n_285),
.B1(n_346),
.B2(n_348),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_434),
.B1(n_442),
.B2(n_403),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_433),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_373),
.A2(n_280),
.B1(n_319),
.B2(n_289),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_342),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_439),
.C(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_395),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_440),
.Y(n_467)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_376),
.A2(n_319),
.B1(n_337),
.B2(n_320),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_444),
.A2(n_449),
.B1(n_452),
.B2(n_464),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_453),
.B1(n_411),
.B2(n_437),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_383),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_448),
.B(n_412),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_417),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_458),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_421),
.A2(n_395),
.B1(n_402),
.B2(n_370),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_387),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_455),
.B(n_459),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_387),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_409),
.A2(n_400),
.B(n_404),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_472),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_374),
.Y(n_463)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_466),
.B(n_431),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_468),
.A2(n_326),
.B1(n_276),
.B2(n_270),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_409),
.A2(n_391),
.B(n_396),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_473),
.Y(n_480)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_474),
.B(n_407),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_456),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_485),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_494),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_482),
.A2(n_489),
.B1(n_491),
.B2(n_496),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_431),
.C(n_427),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_493),
.C(n_465),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_463),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_473),
.B(n_379),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_467),
.Y(n_523)
);

BUFx5_ASAP7_75t_L g487 ( 
.A(n_462),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_487),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_466),
.B(n_439),
.Y(n_488)
);

XNOR2x1_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_450),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_453),
.A2(n_435),
.B1(n_442),
.B2(n_440),
.Y(n_489)
);

HAxp5_ASAP7_75t_SL g490 ( 
.A(n_460),
.B(n_420),
.CON(n_490),
.SN(n_490)
);

NOR3xp33_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_447),
.C(n_467),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_454),
.A2(n_415),
.B1(n_416),
.B2(n_429),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_446),
.B(n_436),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_497),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_414),
.C(n_418),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_495),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_454),
.A2(n_434),
.B1(n_419),
.B2(n_408),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_394),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_452),
.A2(n_441),
.B1(n_393),
.B2(n_334),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_500),
.B1(n_443),
.B2(n_469),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_302),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_468),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_461),
.A2(n_327),
.B1(n_281),
.B2(n_274),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_501),
.A2(n_462),
.B1(n_458),
.B2(n_457),
.Y(n_507)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_502),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_503),
.B(n_513),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_470),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_505),
.B(n_519),
.Y(n_542)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_506),
.B(n_512),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_507),
.A2(n_508),
.B1(n_523),
.B2(n_496),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_510),
.Y(n_537)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_478),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_476),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_514),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_521),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_493),
.A2(n_471),
.B(n_447),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_518),
.B(n_524),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_450),
.Y(n_519)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_522),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_461),
.C(n_469),
.Y(n_524)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_515),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_526),
.B(n_528),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_504),
.A2(n_480),
.B(n_483),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_527),
.A2(n_519),
.B(n_474),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_497),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_514),
.A2(n_520),
.B1(n_498),
.B2(n_501),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_531),
.B(n_532),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_481),
.C(n_494),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_489),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_533),
.B(n_535),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_482),
.Y(n_535)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_539),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_499),
.C(n_443),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_541),
.B(n_505),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_544),
.B(n_547),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_527),
.A2(n_490),
.B1(n_507),
.B2(n_520),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_546),
.A2(n_540),
.B1(n_530),
.B2(n_538),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_511),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_537),
.A2(n_516),
.B(n_521),
.Y(n_548)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_548),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_511),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_553),
.Y(n_562)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_540),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_550),
.A2(n_546),
.B1(n_545),
.B2(n_554),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_551),
.A2(n_150),
.B1(n_11),
.B2(n_14),
.Y(n_569)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_525),
.B(n_500),
.Y(n_552)
);

CKINVDCx14_ASAP7_75t_R g565 ( 
.A(n_552),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_457),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_326),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_556),
.B(n_529),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_537),
.A2(n_218),
.B(n_231),
.Y(n_557)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_557),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_542),
.C(n_529),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_559),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_549),
.B(n_542),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_569),
.Y(n_574)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_564),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_552),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_124),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_567),
.B(n_557),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_573),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_561),
.A2(n_551),
.B(n_553),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_571),
.A2(n_558),
.B(n_569),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_562),
.B(n_564),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_576),
.B(n_577),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_562),
.B(n_556),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_560),
.B(n_552),
.C(n_548),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_578),
.B(n_8),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_572),
.A2(n_565),
.B1(n_563),
.B2(n_568),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_582),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_580),
.A2(n_575),
.B(n_574),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_578),
.A2(n_16),
.B1(n_11),
.B2(n_14),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_584),
.B(n_574),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_585),
.B(n_583),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_586),
.A2(n_588),
.B(n_583),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_581),
.A2(n_8),
.B(n_11),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_589),
.A2(n_590),
.B(n_587),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_591),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_14),
.C(n_15),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_15),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_16),
.Y(n_595)
);


endmodule