module fake_jpeg_31676_n_523 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_523);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_523;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_51),
.B(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_63),
.Y(n_114)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_16),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_68),
.B(n_74),
.Y(n_148)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx2_ASAP7_75t_R g73 ( 
.A(n_38),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_24),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_32),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_81),
.B(n_85),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_24),
.Y(n_83)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_1),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_28),
.B(n_1),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_1),
.Y(n_109)
);

BUFx3_ASAP7_75t_SL g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_25),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_123),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_110),
.B(n_124),
.Y(n_167)
);

BUFx4f_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_26),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_131),
.B(n_40),
.Y(n_200)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_94),
.Y(n_138)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_83),
.A2(n_73),
.B1(n_82),
.B2(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_142),
.A2(n_79),
.B1(n_76),
.B2(n_66),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_90),
.B(n_45),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_26),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_60),
.B(n_27),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_69),
.Y(n_178)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_75),
.Y(n_198)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_165),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_71),
.C(n_67),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_189),
.C(n_195),
.Y(n_225)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_173),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_64),
.B1(n_53),
.B2(n_61),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_174),
.A2(n_199),
.B1(n_210),
.B2(n_220),
.Y(n_238)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_178),
.B(n_192),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_78),
.B1(n_62),
.B2(n_55),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_179),
.A2(n_43),
.B1(n_58),
.B2(n_49),
.Y(n_270)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_117),
.A2(n_52),
.B1(n_88),
.B2(n_84),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_139),
.B1(n_159),
.B2(n_112),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_194),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx6_ASAP7_75t_SL g247 ( 
.A(n_183),
.Y(n_247)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_94),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_217),
.Y(n_237)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_96),
.C(n_86),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_150),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_102),
.B(n_45),
.C(n_27),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_47),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_197),
.B(n_200),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_202),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_104),
.A2(n_89),
.B1(n_77),
.B2(n_49),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_40),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_213),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_207),
.A2(n_69),
.B1(n_37),
.B2(n_44),
.Y(n_271)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_152),
.A2(n_89),
.B1(n_77),
.B2(n_49),
.Y(n_210)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_211),
.Y(n_246)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_19),
.Y(n_213)
);

AO22x2_ASAP7_75t_L g214 ( 
.A1(n_142),
.A2(n_69),
.B1(n_43),
.B2(n_42),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_215),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_103),
.A2(n_19),
.B1(n_48),
.B2(n_47),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_114),
.B(n_48),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_219),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_121),
.B(n_35),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_111),
.B(n_35),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_113),
.A2(n_108),
.B1(n_141),
.B2(n_160),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_143),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_226),
.B(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_191),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_228),
.B(n_240),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_149),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_187),
.A2(n_166),
.B(n_169),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_210),
.B(n_199),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_217),
.B1(n_112),
.B2(n_159),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_258),
.B1(n_270),
.B2(n_208),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_111),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_202),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_181),
.A2(n_147),
.B1(n_139),
.B2(n_160),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_250),
.A2(n_254),
.B1(n_255),
.B2(n_194),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_111),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_261),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_141),
.B1(n_136),
.B2(n_113),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_108),
.B1(n_144),
.B2(n_130),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_179),
.A2(n_163),
.B1(n_158),
.B2(n_42),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_174),
.A2(n_43),
.B1(n_136),
.B2(n_143),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_125),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_186),
.A2(n_125),
.B1(n_115),
.B2(n_49),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_194),
.B(n_211),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_168),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_272),
.B(n_304),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_223),
.B(n_220),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_238),
.A2(n_203),
.B1(n_173),
.B2(n_165),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_278),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_288),
.B1(n_289),
.B2(n_293),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_242),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_281),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_221),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_284),
.A2(n_291),
.B1(n_230),
.B2(n_236),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_290),
.Y(n_332)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_286),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_256),
.A2(n_204),
.B1(n_196),
.B2(n_183),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_250),
.B1(n_226),
.B2(n_228),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_244),
.A2(n_171),
.B(n_168),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_237),
.A2(n_170),
.B1(n_175),
.B2(n_164),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_227),
.B(n_170),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_292),
.B(n_300),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_180),
.B1(n_176),
.B2(n_184),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_235),
.B(n_184),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_306),
.Y(n_315)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_227),
.B(n_171),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_301),
.B(n_302),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_46),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_46),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_303),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_237),
.B(n_46),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_255),
.A2(n_46),
.B1(n_37),
.B2(n_5),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_230),
.B1(n_236),
.B2(n_229),
.Y(n_338)
);

INVx4_ASAP7_75t_SL g306 ( 
.A(n_263),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_240),
.B(n_46),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_309),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_225),
.B(n_37),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_310),
.Y(n_346)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

INVx13_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_312),
.Y(n_351)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_314),
.A2(n_229),
.B1(n_233),
.B2(n_239),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_245),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_320),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_313),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_272),
.B(n_225),
.C(n_237),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_304),
.C(n_259),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_341),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_284),
.A2(n_257),
.B1(n_253),
.B2(n_234),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_333),
.A2(n_336),
.B1(n_337),
.B2(n_343),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_293),
.A2(n_247),
.B1(n_253),
.B2(n_257),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_336),
.B1(n_306),
.B2(n_333),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_274),
.A2(n_234),
.B1(n_270),
.B2(n_229),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_338),
.A2(n_306),
.B1(n_286),
.B2(n_307),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_265),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_274),
.A2(n_288),
.B1(n_289),
.B2(n_294),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_295),
.A2(n_231),
.B1(n_224),
.B2(n_269),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_344),
.A2(n_349),
.B1(n_3),
.B2(n_4),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_224),
.Y(n_345)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_231),
.Y(n_348)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_279),
.A2(n_273),
.B1(n_298),
.B2(n_294),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_341),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_320),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_322),
.B(n_280),
.Y(n_355)
);

NAND3xp33_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_340),
.C(n_342),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_317),
.A2(n_276),
.B(n_290),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_356),
.B(n_358),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_325),
.A2(n_298),
.B1(n_291),
.B2(n_305),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_365),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_285),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_332),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_323),
.Y(n_361)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_269),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_364),
.B(n_367),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_325),
.A2(n_298),
.B1(n_300),
.B2(n_307),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_366),
.A2(n_338),
.B1(n_319),
.B2(n_334),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_315),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_384),
.C(n_350),
.Y(n_397)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_304),
.B(n_312),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_381),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_321),
.A2(n_282),
.B(n_267),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_378),
.B(n_380),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_308),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_372),
.B(n_374),
.Y(n_411)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_345),
.Y(n_373)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_348),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_375),
.A2(n_351),
.B1(n_323),
.B2(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_315),
.B(n_312),
.Y(n_378)
);

OAI22x1_ASAP7_75t_L g379 ( 
.A1(n_328),
.A2(n_248),
.B1(n_314),
.B2(n_296),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_383),
.B1(n_324),
.B2(n_340),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_319),
.A2(n_311),
.B(n_248),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_327),
.A2(n_267),
.B1(n_37),
.B2(n_5),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_37),
.Y(n_382)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_382),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_3),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_326),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_396),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_387),
.A2(n_400),
.B1(n_401),
.B2(n_414),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_318),
.Y(n_391)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_378),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_412),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_393),
.A2(n_376),
.B1(n_379),
.B2(n_370),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_401),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_363),
.A2(n_334),
.B1(n_329),
.B2(n_346),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_363),
.A2(n_329),
.B1(n_346),
.B2(n_330),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_318),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_371),
.B(n_330),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_413),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_351),
.Y(n_407)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_339),
.B(n_352),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_409),
.A2(n_357),
.B(n_342),
.Y(n_438)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_352),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_360),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_415),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_389),
.A2(n_373),
.B1(n_362),
.B2(n_383),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_422),
.B1(n_440),
.B2(n_387),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_426),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_368),
.C(n_359),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_424),
.C(n_431),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_376),
.B1(n_359),
.B2(n_362),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_436),
.B1(n_394),
.B2(n_399),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_384),
.C(n_378),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_394),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_430),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_356),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_381),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_433),
.Y(n_458)
);

OAI211xp5_ASAP7_75t_L g435 ( 
.A1(n_406),
.A2(n_380),
.B(n_382),
.C(n_365),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_435),
.B(n_409),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_390),
.B1(n_411),
.B2(n_408),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_382),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_395),
.C(n_412),
.Y(n_450)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_438),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_408),
.A2(n_390),
.B1(n_388),
.B2(n_415),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_441),
.A2(n_434),
.B1(n_404),
.B2(n_6),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_409),
.Y(n_443)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_444),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_427),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_454),
.Y(n_476)
);

NAND2x1_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_392),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_448),
.B(n_426),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_432),
.A2(n_388),
.B1(n_405),
.B2(n_392),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_456),
.B1(n_417),
.B2(n_420),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_450),
.B(n_452),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_395),
.C(n_410),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_453),
.C(n_459),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_428),
.C(n_421),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_438),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_418),
.B(n_404),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_457),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_399),
.C(n_385),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_431),
.B(n_361),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_460),
.B(n_6),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_459),
.B(n_453),
.C(n_452),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_463),
.Y(n_484)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_440),
.C(n_437),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_466),
.B(n_469),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_467),
.Y(n_485)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_442),
.A2(n_429),
.B(n_419),
.C(n_427),
.Y(n_468)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_468),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_432),
.C(n_420),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_471),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_473),
.A2(n_458),
.B1(n_442),
.B2(n_449),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_3),
.C(n_5),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_7),
.Y(n_491)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_447),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_451),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_489),
.C(n_463),
.Y(n_494)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_480),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_472),
.A2(n_455),
.B1(n_441),
.B2(n_461),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_465),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_474),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_488),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_470),
.A2(n_455),
.B1(n_461),
.B2(n_447),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_450),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_7),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_491),
.B(n_7),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_467),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_494),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_482),
.A2(n_476),
.B1(n_468),
.B2(n_477),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_496),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_481),
.A2(n_475),
.B1(n_465),
.B2(n_462),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_462),
.C(n_478),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_501),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_499),
.A2(n_500),
.B1(n_481),
.B2(n_490),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_486),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_502),
.B(n_491),
.Y(n_505)
);

AOI21xp33_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_479),
.B(n_485),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_504),
.B(n_505),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_480),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_483),
.Y(n_509)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_498),
.A3(n_501),
.B1(n_497),
.B2(n_494),
.C1(n_8),
.C2(n_12),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_512),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_10),
.C(n_11),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_513),
.B(n_509),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_515),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_503),
.C(n_510),
.Y(n_516)
);

AOI322xp5_ASAP7_75t_L g518 ( 
.A1(n_516),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_508),
.C2(n_514),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_12),
.C(n_10),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_517),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_520),
.A2(n_11),
.B(n_12),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_11),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_522),
.Y(n_523)
);


endmodule