module real_jpeg_24260_n_16 (n_350, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_350;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_65),
.B1(n_68),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_29),
.B1(n_32),
.B2(n_76),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_76),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_1),
.A2(n_76),
.B1(n_82),
.B2(n_93),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_48),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_2),
.A2(n_48),
.B1(n_65),
.B2(n_68),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_2),
.A2(n_48),
.B1(n_80),
.B2(n_93),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_4),
.A2(n_60),
.B1(n_65),
.B2(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_4),
.A2(n_29),
.B1(n_32),
.B2(n_60),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_4),
.A2(n_60),
.B1(n_82),
.B2(n_93),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_38),
.B1(n_65),
.B2(n_68),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_L g283 ( 
.A1(n_6),
.A2(n_38),
.B1(n_85),
.B2(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_SL g89 ( 
.A(n_7),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_8),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_8),
.A2(n_33),
.B1(n_65),
.B2(n_68),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_8),
.A2(n_33),
.B1(n_82),
.B2(n_92),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_67),
.B1(n_82),
.B2(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_9),
.A2(n_29),
.B1(n_32),
.B2(n_67),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_11),
.B(n_94),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_11),
.B(n_29),
.C(n_42),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_74),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_28),
.B1(n_115),
.B2(n_172),
.Y(n_171)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_13),
.A2(n_79),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_65),
.B1(n_68),
.B2(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_13),
.A2(n_29),
.B1(n_32),
.B2(n_98),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_342),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_329),
.B(n_341),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_296),
.A3(n_322),
.B1(n_327),
.B2(n_328),
.C(n_350),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_270),
.B(n_295),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_246),
.B(n_269),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_136),
.B(n_220),
.C(n_245),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_120),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_23),
.B(n_120),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_99),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_25),
.B(n_55),
.C(n_99),
.Y(n_221)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_39),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_27),
.B(n_39),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_34),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_28),
.A2(n_31),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_28),
.B(n_37),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_28),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_28),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_28),
.A2(n_36),
.B1(n_165),
.B2(n_172),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_28),
.A2(n_30),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_30),
.Y(n_134)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_32),
.B(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_35),
.A2(n_159),
.B(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_49),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_40),
.A2(n_52),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_40),
.A2(n_52),
.B1(n_148),
.B2(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_40),
.B(n_83),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_40),
.A2(n_44),
.B1(n_52),
.B2(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_40),
.A2(n_52),
.B(n_58),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_46),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_45),
.B(n_65),
.C(n_72),
.Y(n_188)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_46),
.B(n_144),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_46),
.A2(n_71),
.B(n_187),
.C(n_188),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_49),
.B(n_210),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_51),
.A2(n_62),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_58),
.B(n_61),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_52),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_52),
.A2(n_61),
.B(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.C(n_77),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_56),
.A2(n_57),
.B1(n_63),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_59),
.B(n_62),
.Y(n_210)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_64),
.Y(n_129)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_65),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_68),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_84),
.B(n_88),
.C(n_118),
.Y(n_117)
);

HAxp5_ASAP7_75t_SL g187 ( 
.A(n_65),
.B(n_83),
.CON(n_187),
.SN(n_187)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_89),
.C(n_93),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_69),
.A2(n_74),
.B1(n_128),
.B2(n_187),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_69),
.B(n_234),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_69),
.A2(n_74),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_69),
.A2(n_74),
.B(n_110),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_70),
.A2(n_108),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_70),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_74),
.B(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_86),
.B1(n_94),
.B2(n_95),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B(n_84),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_83),
.B(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_85),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_86),
.A2(n_94),
.B1(n_105),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_86),
.B(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_86),
.A2(n_94),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_86),
.A2(n_320),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_96),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_87),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_94),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_94),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_111),
.B2(n_119),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_102),
.B(n_106),
.C(n_119),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_103),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_103),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_108),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_108),
.A2(n_233),
.B(n_292),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_109),
.B(n_265),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_110),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_117),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_124),
.B(n_125),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.C(n_132),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_135),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_219),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_214),
.B(n_218),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_199),
.B(n_213),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_183),
.B(n_198),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_160),
.B(n_182),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_157),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_169),
.B(n_181),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_167),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_177),
.B(n_180),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_197),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_197),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_193),
.C(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_201),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_208),
.C(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_222),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_244),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_235),
.B1(n_242),
.B2(n_243),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_228),
.C(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_242),
.C(n_244),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_248),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_268),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_256),
.C(n_268),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_252),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_251),
.A2(n_276),
.B(n_280),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_254),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_254),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_266),
.B2(n_267),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_263),
.C(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_261),
.B(n_302),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_262),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_271),
.B(n_272),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_294),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_286),
.B2(n_287),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_286),
.C(n_294),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_285),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_282),
.Y(n_336)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B(n_293),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_293),
.A2(n_298),
.B1(n_309),
.B2(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_311),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_311),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_309),
.C(n_310),
.Y(n_297)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_308),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_300),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_304),
.C(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_314),
.C(n_321),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_306),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_307),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_316),
.C(n_318),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_321),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_331),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_339),
.B2(n_340),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_334),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_335),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_337),
.C(n_339),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_344),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_348),
.Y(n_347)
);


endmodule