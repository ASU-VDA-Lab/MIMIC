module fake_jpeg_22468_n_282 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_18),
.B1(n_20),
.B2(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_40),
.B1(n_35),
.B2(n_28),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_37),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_49),
.B1(n_50),
.B2(n_35),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_28),
.B1(n_32),
.B2(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_39),
.B1(n_37),
.B2(n_28),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_39),
.B1(n_37),
.B2(n_46),
.Y(n_95)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_66),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_69),
.B1(n_81),
.B2(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_62),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_52),
.B(n_53),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_73),
.C(n_74),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_36),
.C(n_33),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_36),
.C(n_33),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_35),
.B1(n_36),
.B2(n_24),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_48),
.B1(n_46),
.B2(n_31),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_83),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_27),
.B1(n_29),
.B2(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_19),
.B1(n_16),
.B2(n_24),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_19),
.B1(n_16),
.B2(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_31),
.Y(n_85)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_111),
.B1(n_64),
.B2(n_78),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_99),
.B1(n_83),
.B2(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_95),
.B1(n_59),
.B2(n_76),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_96),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_103),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_27),
.B1(n_29),
.B2(n_46),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_25),
.C(n_27),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_88),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_25),
.B1(n_22),
.B2(n_3),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_77),
.B1(n_71),
.B2(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_117),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_68),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_95),
.B(n_91),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_59),
.Y(n_116)
);

OA21x2_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_95),
.B(n_89),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_119),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_120),
.A2(n_130),
.B(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_84),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_84),
.B1(n_74),
.B2(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_126),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_110),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_127),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_135),
.B(n_2),
.Y(n_168)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_134),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_59),
.B1(n_25),
.B2(n_22),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_1),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_87),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_149),
.B(n_162),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_122),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_147),
.C(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_88),
.C(n_94),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_103),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_159),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_94),
.A3(n_102),
.B1(n_95),
.B2(n_104),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_126),
.B(n_118),
.C(n_115),
.D(n_129),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_111),
.C(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_2),
.C(n_4),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_5),
.C(n_6),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_101),
.C(n_5),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_138),
.C(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_118),
.B1(n_126),
.B2(n_163),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_167),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_180),
.C(n_189),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_127),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_183),
.B(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_181),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_194),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_182),
.B(n_172),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_195),
.B(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_117),
.C(n_7),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_159),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_6),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_179),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_153),
.B1(n_143),
.B2(n_154),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_214),
.B1(n_211),
.B2(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_147),
.C(n_143),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_174),
.C(n_180),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_153),
.B1(n_169),
.B2(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_173),
.B1(n_182),
.B2(n_190),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_143),
.B(n_157),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_214),
.B(n_212),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_221),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_227),
.B1(n_218),
.B2(n_198),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_227),
.B(n_230),
.Y(n_242)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_201),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_204),
.B(n_177),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

XOR2x2_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_189),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_203),
.B(n_202),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g235 ( 
.A(n_231),
.B(n_210),
.C(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_206),
.CI(n_199),
.CON(n_244),
.SN(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_228),
.C(n_215),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_233),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_249),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_201),
.C(n_226),
.Y(n_250)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_242),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_244),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_254),
.B1(n_255),
.B2(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_208),
.B1(n_217),
.B2(n_219),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_R g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_244),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_245),
.B1(n_253),
.B2(n_255),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_266),
.B1(n_197),
.B2(n_155),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_248),
.C(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_234),
.C(n_148),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_224),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_269),
.B(n_270),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_241),
.A3(n_262),
.B1(n_237),
.B2(n_204),
.C1(n_219),
.C2(n_155),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_148),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_175),
.B1(n_213),
.B2(n_166),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_7),
.Y(n_277)
);

AOI321xp33_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_267),
.A3(n_166),
.B1(n_8),
.B2(n_11),
.C(n_6),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_271),
.C(n_8),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_275),
.B1(n_11),
.B2(n_12),
.Y(n_280)
);

NAND4xp25_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_278),
.C(n_12),
.D(n_14),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_281),
.Y(n_282)
);


endmodule