module real_jpeg_9399_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_315, n_6, n_314, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_315;
input n_6;
input n_314;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_16),
.B(n_28),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_2),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_78),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_97),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_97),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_97),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_43),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_4),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_5),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_102),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_102),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_102),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_31),
.B(n_63),
.C(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_31),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_11),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_109),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_109),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_12),
.A2(n_35),
.B1(n_65),
.B2(n_66),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_13),
.A2(n_50),
.B1(n_65),
.B2(n_66),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_50),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_15),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_138),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_138),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_138),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_16),
.A2(n_31),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_16),
.B(n_31),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_16),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_16),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_16),
.A2(n_27),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_27),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_16),
.B(n_51),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_16),
.A2(n_40),
.B1(n_41),
.B2(n_122),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_17),
.A2(n_40),
.B1(n_41),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_17),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_60),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_60),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_85),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_83),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_70),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_52),
.B1(n_53),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_25),
.A2(n_30),
.B1(n_56),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_25),
.A2(n_30),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_25),
.A2(n_30),
.B1(n_147),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_25),
.A2(n_30),
.B1(n_163),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_25),
.A2(n_30),
.B1(n_203),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_25),
.A2(n_30),
.B1(n_214),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_25),
.A2(n_30),
.B1(n_240),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_25),
.A2(n_30),
.B1(n_82),
.B2(n_258),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_29),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_30),
.B(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_31),
.B(n_33),
.Y(n_151)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_32),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_45),
.B1(n_48),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_46),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_41),
.A2(n_46),
.B(n_122),
.C(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_44),
.A2(n_51),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_48),
.B1(n_59),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_45),
.A2(n_48),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_45),
.A2(n_48),
.B1(n_218),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_45),
.A2(n_48),
.B1(n_243),
.B2(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_45),
.A2(n_48),
.B1(n_77),
.B2(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.C(n_61),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_61),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_64),
.B(n_68),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_64),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_64),
.B1(n_108),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_64),
.B1(n_135),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_62),
.A2(n_64),
.B1(n_143),
.B2(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_62),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_62),
.A2(n_64),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_62),
.A2(n_64),
.B1(n_226),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_62),
.A2(n_64),
.B1(n_235),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_62),
.A2(n_64),
.B1(n_68),
.B2(n_267),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_64),
.B(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_64),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_65),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_65),
.B(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.C(n_79),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_301),
.Y(n_306)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_76),
.C(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_76),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_76),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_79),
.B(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_298),
.A3(n_307),
.B1(n_310),
.B2(n_311),
.C(n_314),
.Y(n_85)
);

AOI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_251),
.A3(n_286),
.B1(n_292),
.B2(n_297),
.C(n_315),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_208),
.C(n_247),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_178),
.B(n_207),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_157),
.B(n_177),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_140),
.B(n_156),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_129),
.B(n_139),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_115),
.B(n_128),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_98),
.A2(n_99),
.B1(n_155),
.B2(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_119),
.B1(n_120),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_110),
.B2(n_114),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_123),
.B(n_127),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_121),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_120),
.B1(n_137),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_119),
.A2(n_120),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_119),
.A2(n_120),
.B1(n_189),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_119),
.A2(n_120),
.B1(n_223),
.B2(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_119),
.A2(n_120),
.B(n_233),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_141),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.CI(n_136),
.CON(n_132),
.SN(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.CI(n_148),
.CON(n_141),
.SN(n_141)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_170),
.B2(n_171),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_173),
.C(n_175),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_169),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_180),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_192),
.C(n_193),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_187),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_201),
.C(n_204),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_209),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_228),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_210),
.B(n_228),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_221),
.C(n_227),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_219),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_SL g245 ( 
.A(n_215),
.B(n_219),
.C(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_227),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_245),
.B2(n_246),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_231),
.B(n_236),
.C(n_246),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_234),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_241),
.C(n_244),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_239),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_270),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_252),
.B(n_270),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.C(n_269),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_254),
.B1(n_263),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_259),
.C(n_262),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_257),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_263),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_265),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_280),
.B(n_282),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_266),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_284),
.B2(n_285),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_277),
.C(n_285),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B(n_276),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_300),
.C(n_304),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_276),
.B(n_300),
.CI(n_304),
.CON(n_309),
.SN(n_309)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_282),
.B2(n_283),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_305),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_309),
.Y(n_313)
);


endmodule