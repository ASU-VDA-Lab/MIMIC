module real_jpeg_13222_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_271, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_271;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_255;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_267;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_2),
.A2(n_60),
.B1(n_62),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_107)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_4),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_97),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_4),
.A2(n_60),
.B1(n_62),
.B2(n_97),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_4),
.A2(n_31),
.B1(n_33),
.B2(n_97),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_6),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_60),
.B1(n_62),
.B2(n_78),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_31),
.B1(n_33),
.B2(n_78),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_41),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_41),
.B1(n_60),
.B2(n_62),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g233 ( 
.A(n_11),
.B(n_31),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_60),
.C(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_12),
.B(n_34),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_12),
.A2(n_63),
.B(n_151),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_12),
.A2(n_32),
.B(n_33),
.C(n_178),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_12),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_12),
.B(n_44),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_13),
.A2(n_31),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_13),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_13),
.A2(n_38),
.B1(n_60),
.B2(n_62),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_54),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_54),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_54),
.B1(n_60),
.B2(n_62),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_15),
.A2(n_46),
.B1(n_60),
.B2(n_62),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_15),
.A2(n_31),
.B1(n_33),
.B2(n_46),
.Y(n_224)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_21),
.B(n_101),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_89),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_22),
.A2(n_23),
.B1(n_81),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_80),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_42),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_26),
.B(n_42),
.C(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_27),
.A2(n_39),
.B1(n_40),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_27),
.A2(n_183),
.B(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_27),
.A2(n_39),
.B1(n_197),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_27),
.A2(n_184),
.B(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_28),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_35),
.B(n_136),
.Y(n_178)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_33),
.A2(n_45),
.A3(n_49),
.B1(n_221),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_34),
.B(n_100),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_35),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_36),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_37),
.A2(n_39),
.B(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_39),
.A2(n_99),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B(n_51),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_47),
.B1(n_48),
.B2(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_45),
.A2(n_47),
.B(n_136),
.C(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_48),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_48),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_48),
.A2(n_96),
.B(n_118),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_52),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_56),
.A2(n_69),
.B1(n_70),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_56),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_62),
.B(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_63),
.A2(n_68),
.B1(n_180),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_63),
.A2(n_68),
.B1(n_204),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_65),
.B(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_64),
.A2(n_65),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_65),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_68),
.A2(n_157),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_68),
.B(n_136),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_68),
.A2(n_165),
.B(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_77),
.B2(n_79),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_72),
.B1(n_79),
.B2(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_77),
.B1(n_79),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_72),
.B(n_138),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_72),
.A2(n_79),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_87),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_76),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_76),
.B(n_136),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_76),
.A2(n_148),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_81),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_88),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_83),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_88),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_89),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_98),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_90),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_91),
.B(n_93),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_92),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_94),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_95),
.B(n_98),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_123),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_111),
.B2(n_112),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_110),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_108),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_106),
.A2(n_137),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_121),
.B2(n_122),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_264),
.B(n_269),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_238),
.A3(n_257),
.B1(n_262),
.B2(n_263),
.C(n_271),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_213),
.B(n_237),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_191),
.B(n_212),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_173),
.B(n_190),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_153),
.B(n_172),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_134),
.B1(n_139),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_146),
.C(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_161),
.B(n_171),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_166),
.B(n_170),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_175),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_185),
.C(n_189),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_179),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_205),
.B2(n_206),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_208),
.C(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_199),
.C(n_203),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_215),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_228),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_229),
.C(n_230),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_222),
.B2(n_227),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_223),
.C(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_250),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_250),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_248),
.C(n_249),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_241),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_247),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_254),
.C(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_268),
.Y(n_269)
);


endmodule