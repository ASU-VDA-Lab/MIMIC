module fake_jpeg_12505_n_352 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_51),
.Y(n_86)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_51),
.B1(n_45),
.B2(n_36),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_59),
.A2(n_80),
.B1(n_35),
.B2(n_20),
.Y(n_108)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_17),
.B1(n_19),
.B2(n_33),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_46),
.B1(n_54),
.B2(n_29),
.Y(n_90)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_76),
.Y(n_94)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_37),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_71),
.A2(n_77),
.B1(n_81),
.B2(n_34),
.Y(n_119)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_17),
.B1(n_18),
.B2(n_31),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_41),
.A2(n_18),
.B1(n_34),
.B2(n_35),
.Y(n_81)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_16),
.Y(n_98)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_108),
.B1(n_121),
.B2(n_47),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_107),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_97),
.B(n_98),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_39),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_124),
.C(n_43),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_38),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_41),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_109),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_20),
.B(n_33),
.C(n_32),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_110),
.B(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_49),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_24),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_24),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_32),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_125),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_35),
.B1(n_47),
.B2(n_43),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_61),
.B(n_29),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_34),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_50),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_129),
.B(n_2),
.Y(n_185)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_72),
.B1(n_84),
.B2(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_136),
.B1(n_137),
.B2(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_72),
.B1(n_43),
.B2(n_74),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_78),
.B1(n_70),
.B2(n_55),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_90),
.A2(n_70),
.B1(n_56),
.B2(n_55),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_149),
.B1(n_102),
.B2(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_143),
.Y(n_170)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_56),
.B1(n_82),
.B2(n_34),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_34),
.B1(n_50),
.B2(n_28),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_102),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_50),
.B(n_9),
.C(n_10),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_10),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_125),
.B1(n_94),
.B2(n_106),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_124),
.B1(n_96),
.B2(n_95),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_104),
.B(n_103),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_176),
.B(n_180),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_160),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_99),
.B1(n_110),
.B2(n_97),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_174),
.B1(n_183),
.B2(n_136),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_162),
.B(n_177),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_163),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_93),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_166),
.B(n_175),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_112),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_93),
.B(n_114),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_104),
.B(n_103),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_99),
.B1(n_96),
.B2(n_126),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_95),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_149),
.B(n_124),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_96),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_145),
.B1(n_131),
.B2(n_146),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_133),
.B1(n_142),
.B2(n_151),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_128),
.A2(n_50),
.B1(n_9),
.B2(n_11),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_135),
.C(n_147),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_2),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_2),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_138),
.B(n_15),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_3),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_129),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_220),
.C(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_197),
.B(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_217),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_219),
.B1(n_165),
.B2(n_194),
.Y(n_235)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_223),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_174),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_211),
.B(n_213),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_158),
.B(n_143),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_169),
.B(n_176),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_144),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_171),
.A2(n_137),
.B1(n_132),
.B2(n_130),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_218),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g216 ( 
.A1(n_172),
.A2(n_158),
.B(n_7),
.C(n_11),
.D(n_12),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_167),
.C(n_184),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_3),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_7),
.C(n_11),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_189),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_173),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_228),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_4),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_226),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_12),
.B1(n_14),
.B2(n_6),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_4),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_164),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_188),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_234),
.C(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_188),
.C(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_244),
.B1(n_210),
.B2(n_196),
.Y(n_259)
);

OAI211xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_180),
.B(n_191),
.C(n_178),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_241),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_186),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_239),
.A2(n_256),
.B(n_223),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_184),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_196),
.A2(n_207),
.B1(n_224),
.B2(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_167),
.B1(n_165),
.B2(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_179),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_251),
.C(n_227),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_250),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_170),
.C(n_160),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_183),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_271),
.B1(n_273),
.B2(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_240),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_205),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_264),
.C(n_267),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_200),
.C(n_198),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_214),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_208),
.C(n_215),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_208),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_272),
.C(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_226),
.B1(n_223),
.B2(n_209),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_220),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_216),
.B1(n_14),
.B2(n_5),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_255),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_4),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_279),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_239),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_232),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_234),
.B(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_285),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_243),
.B1(n_251),
.B2(n_256),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_267),
.B(n_249),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_289),
.A2(n_243),
.B1(n_256),
.B2(n_261),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_277),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_253),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_253),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_261),
.C(n_262),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_302),
.Y(n_323)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_263),
.C(n_268),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_281),
.B(n_294),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_281),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_310),
.Y(n_314)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_272),
.C(n_257),
.Y(n_310)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_266),
.C(n_275),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_308),
.B(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_282),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_320),
.B(n_322),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_305),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_307),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_301),
.Y(n_333)
);

XOR2x2_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_285),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_318),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_286),
.B1(n_289),
.B2(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_329),
.Y(n_338)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_298),
.B(n_297),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_332),
.B(n_319),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_287),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_330),
.B(n_334),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_299),
.C(n_311),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_304),
.C(n_295),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_314),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_337),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_340),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_316),
.B(n_313),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_333),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_317),
.C(n_306),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_341),
.B(n_334),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_344),
.B(n_338),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_346),
.A2(n_347),
.B(n_284),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_342),
.A2(n_280),
.B(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_345),
.C(n_252),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_252),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_273),
.C(n_5),
.Y(n_352)
);


endmodule