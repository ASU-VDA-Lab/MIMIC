module fake_jpeg_9227_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_7),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_23),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_16),
.B1(n_27),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_53),
.B1(n_57),
.B2(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_20),
.B1(n_27),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_36),
.B1(n_45),
.B2(n_20),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_71),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_72),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_0),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_24),
.B1(n_44),
.B2(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_94),
.B1(n_112),
.B2(n_63),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_81),
.B(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_92),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_44),
.B1(n_41),
.B2(n_46),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_105),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_46),
.C(n_48),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_106),
.C(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_54),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_35),
.B1(n_19),
.B2(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_31),
.C(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_111),
.B1(n_25),
.B2(n_1),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_58),
.B1(n_54),
.B2(n_74),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_43),
.C(n_31),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_58),
.A2(n_31),
.A3(n_34),
.B1(n_33),
.B2(n_26),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_35),
.A3(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_117),
.A2(n_25),
.B1(n_9),
.B2(n_13),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_137),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_99),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_35),
.C(n_28),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_132),
.C(n_113),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_133),
.B1(n_127),
.B2(n_122),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_35),
.C(n_28),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_114),
.B1(n_104),
.B2(n_98),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_105),
.B(n_98),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_84),
.B(n_82),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_159),
.B(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_152),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_149),
.A2(n_160),
.B1(n_171),
.B2(n_91),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_135),
.Y(n_184)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_158),
.B(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_111),
.B1(n_110),
.B2(n_108),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_84),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_85),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_82),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_165),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_99),
.B(n_95),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_101),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_11),
.B1(n_128),
.B2(n_4),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_115),
.B(n_99),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_174),
.B(n_129),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_92),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_81),
.B1(n_107),
.B2(n_83),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_180),
.B1(n_139),
.B2(n_140),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_8),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_135),
.C(n_120),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_0),
.B(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_97),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_2),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_96),
.B1(n_91),
.B2(n_8),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_146),
.B1(n_124),
.B2(n_10),
.Y(n_194)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_182),
.A2(n_191),
.B(n_195),
.Y(n_238)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_206),
.C(n_193),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_187),
.A2(n_205),
.B1(n_195),
.B2(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_197),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_156),
.B(n_154),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_199),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_198),
.B1(n_171),
.B2(n_152),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_8),
.B1(n_13),
.B2(n_11),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_148),
.B(n_13),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_140),
.B1(n_91),
.B2(n_128),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_163),
.A3(n_175),
.B1(n_149),
.B2(n_155),
.C1(n_160),
.C2(n_168),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_1),
.B(n_2),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_158),
.B(n_178),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_3),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_2),
.C(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_153),
.B(n_6),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_216),
.A2(n_224),
.B(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_219),
.B(n_229),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_178),
.B1(n_179),
.B2(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_178),
.B1(n_157),
.B2(n_5),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_185),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_203),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_233),
.B(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_5),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_5),
.B(n_6),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_236),
.C(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_190),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_6),
.C(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_212),
.C(n_191),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_186),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_182),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_261),
.C(n_238),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_257),
.B1(n_258),
.B2(n_218),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_214),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_186),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_231),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_260),
.B(n_233),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_223),
.B1(n_222),
.B2(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_201),
.B1(n_199),
.B2(n_203),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_196),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_206),
.Y(n_261)
);

AOI22x1_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_194),
.B1(n_184),
.B2(n_209),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_264),
.B1(n_224),
.B2(n_215),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_184),
.B1(n_189),
.B2(n_211),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_234),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_273),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_267),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_276),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_236),
.C(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_271),
.C(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_253),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_215),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_218),
.C(n_228),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_220),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_232),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_247),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_281),
.B1(n_256),
.B2(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_235),
.C(n_221),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_251),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_200),
.B1(n_244),
.B2(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_248),
.B(n_200),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_260),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_254),
.C(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_242),
.Y(n_291)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_294),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_283),
.Y(n_294)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_259),
.B(n_250),
.Y(n_301)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

NOR2x1_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_249),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_301),
.B(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_270),
.C(n_273),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_311),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_250),
.B(n_245),
.Y(n_304)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_299),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_266),
.CI(n_271),
.CON(n_306),
.SN(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_296),
.C(n_285),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_285),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_317),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_321),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_316),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_296),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_289),
.B1(n_297),
.B2(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_289),
.C(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_302),
.C(n_312),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_288),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_308),
.Y(n_327)
);

NOR4xp25_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_316),
.C(n_320),
.D(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_310),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_332),
.C(n_301),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_325),
.B(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_334),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_325),
.C(n_328),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_306),
.Y(n_339)
);


endmodule