module fake_netlist_1_152_n_701 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_701);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_701;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_305;
wire n_100;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_472;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_132;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_75), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_21), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_62), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_12), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_42), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_77), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_48), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_54), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_1), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_24), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_59), .Y(n_92) );
NOR2xp67_ASAP7_75t_L g93 ( .A(n_28), .B(n_36), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_0), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_71), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_15), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_61), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_64), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_16), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_19), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_23), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_56), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_37), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_66), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_12), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_26), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_22), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_24), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_22), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_73), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_32), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_19), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_53), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_31), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_29), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_1), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_45), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_57), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_44), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_39), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_7), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_3), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_40), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_129), .B(n_0), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_103), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_129), .B(n_2), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_103), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_103), .B(n_4), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_102), .B(n_4), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_84), .B(n_5), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_102), .B(n_5), .Y(n_144) );
NAND2xp33_ASAP7_75t_L g145 ( .A(n_89), .B(n_80), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_119), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_118), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_84), .B(n_6), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_92), .B(n_38), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_92), .B(n_35), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_114), .Y(n_158) );
NAND2xp33_ASAP7_75t_R g159 ( .A(n_104), .B(n_41), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_121), .Y(n_161) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_81), .B(n_79), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_81), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_110), .Y(n_164) );
INVxp67_ASAP7_75t_L g165 ( .A(n_91), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_85), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_86), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_125), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_121), .B(n_6), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_89), .Y(n_171) );
OR2x6_ASAP7_75t_L g172 ( .A(n_95), .B(n_8), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_121), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_114), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_86), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_135), .B(n_107), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_146), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_170), .B(n_95), .Y(n_183) );
XOR2xp5_ASAP7_75t_L g184 ( .A(n_169), .B(n_110), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_173), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_165), .B(n_112), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_163), .B(n_108), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_164), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_163), .B(n_128), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_166), .B(n_101), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_170), .B(n_128), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_172), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
BUFx4f_ASAP7_75t_L g198 ( .A(n_172), .Y(n_198) );
AND2x4_ASAP7_75t_SL g199 ( .A(n_172), .B(n_96), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_173), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_155), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_166), .B(n_90), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_167), .B(n_105), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_173), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_156), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_170), .B(n_96), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_167), .B(n_122), .Y(n_209) );
INVx4_ASAP7_75t_SL g210 ( .A(n_150), .Y(n_210) );
INVx5_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_130), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_162), .B(n_88), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_173), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_156), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_168), .B(n_127), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_168), .B(n_126), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_130), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_143), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_175), .B(n_126), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_143), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_130), .Y(n_225) );
INVx4_ASAP7_75t_SL g226 ( .A(n_150), .Y(n_226) );
NAND3x1_ASAP7_75t_L g227 ( .A(n_141), .B(n_98), .C(n_111), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g231 ( .A1(n_162), .A2(n_82), .B1(n_98), .B2(n_111), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_149), .B(n_113), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_158), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_153), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_153), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_188), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_195), .B(n_172), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_186), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_178), .B(n_131), .Y(n_239) );
OR2x6_ASAP7_75t_L g240 ( .A(n_195), .B(n_138), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_192), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_196), .B(n_138), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_199), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_232), .A2(n_138), .B(n_144), .C(n_134), .Y(n_244) );
INVx1_ASAP7_75t_SL g245 ( .A(n_180), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_187), .B(n_175), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_192), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_196), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_213), .B(n_138), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_193), .B(n_175), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_199), .Y(n_254) );
NAND2x2_ASAP7_75t_L g255 ( .A(n_232), .B(n_162), .Y(n_255) );
NAND3xp33_ASAP7_75t_SL g256 ( .A(n_180), .B(n_97), .C(n_113), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_214), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
AND2x6_ASAP7_75t_L g260 ( .A(n_183), .B(n_170), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_214), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_198), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_209), .B(n_137), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_177), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_192), .Y(n_265) );
OR2x4_ASAP7_75t_L g266 ( .A(n_216), .B(n_114), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_179), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_183), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_203), .B(n_137), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_221), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_197), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_185), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_213), .A2(n_137), .B1(n_144), .B2(n_133), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_183), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_228), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_185), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_184), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_191), .B(n_137), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_190), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_231), .A2(n_144), .B1(n_150), .B2(n_152), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_198), .B(n_144), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_213), .A2(n_150), .B1(n_152), .B2(n_136), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_201), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_194), .A2(n_150), .B1(n_152), .B2(n_136), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_184), .Y(n_291) );
OR2x2_ASAP7_75t_SL g292 ( .A(n_227), .B(n_114), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_194), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_228), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_191), .B(n_152), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_194), .A2(n_152), .B1(n_133), .B2(n_161), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_201), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_205), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_205), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_194), .A2(n_152), .B1(n_161), .B2(n_114), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_200), .Y(n_303) );
AOI222xp33_ASAP7_75t_L g304 ( .A1(n_282), .A2(n_208), .B1(n_217), .B2(n_147), .C1(n_148), .C2(n_160), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_236), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_269), .Y(n_310) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_253), .B(n_208), .Y(n_311) );
BUFx6f_ASAP7_75t_SL g312 ( .A(n_254), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_254), .B(n_211), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_278), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_236), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_238), .Y(n_317) );
CKINVDCx16_ASAP7_75t_R g318 ( .A(n_291), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_244), .A2(n_220), .B(n_208), .C(n_204), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_255), .A2(n_208), .B1(n_227), .B2(n_159), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_278), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_237), .B(n_114), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_245), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_251), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
OR2x6_ASAP7_75t_SL g327 ( .A(n_282), .B(n_207), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_251), .Y(n_328) );
BUFx5_ASAP7_75t_L g329 ( .A(n_241), .Y(n_329) );
NOR2xp67_ASAP7_75t_L g330 ( .A(n_256), .B(n_219), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_255), .A2(n_215), .B1(n_207), .B2(n_152), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_239), .B(n_215), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_259), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_250), .A2(n_152), .B1(n_234), .B2(n_230), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_263), .A2(n_235), .B(n_234), .C(n_230), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_249), .B(n_182), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_293), .B(n_219), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_237), .A2(n_211), .B1(n_224), .B2(n_223), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_259), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_258), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_250), .B(n_223), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_249), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_266), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g344 ( .A1(n_237), .A2(n_235), .B1(n_224), .B2(n_160), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_253), .B(n_211), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_237), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_262), .B(n_182), .Y(n_347) );
OR2x6_ASAP7_75t_L g348 ( .A(n_262), .B(n_87), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_240), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_250), .B(n_189), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_240), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_260), .A2(n_211), .B1(n_115), .B2(n_124), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_240), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_250), .B(n_189), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_240), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_264), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_242), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_247), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_247), .B(n_211), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_317), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_335), .A2(n_270), .B(n_297), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_307), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_307), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_335), .A2(n_275), .B(n_301), .C(n_300), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_332), .A2(n_286), .B(n_246), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_322), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_344), .A2(n_260), .B1(n_277), .B2(n_242), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_316), .B(n_242), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_311), .A2(n_242), .B1(n_260), .B2(n_285), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_311), .A2(n_260), .B1(n_283), .B2(n_301), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_349), .A2(n_260), .B1(n_289), .B2(n_300), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_308), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_308), .B(n_267), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_354), .A2(n_358), .B1(n_304), .B2(n_356), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_319), .A2(n_148), .B1(n_139), .B2(n_147), .C(n_252), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_306), .A2(n_260), .B1(n_267), .B2(n_299), .C1(n_268), .C2(n_271), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_323), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_344), .A2(n_260), .B1(n_273), .B2(n_299), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_356), .A2(n_273), .B1(n_279), .B2(n_275), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_326), .B(n_292), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_318), .B(n_292), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_333), .Y(n_385) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_322), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_339), .A2(n_287), .B(n_290), .Y(n_387) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_331), .A2(n_302), .B(n_298), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_339), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_322), .B(n_289), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_139), .B(n_145), .C(n_87), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_346), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_351), .A2(n_348), .B1(n_346), .B2(n_336), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_348), .A2(n_294), .B1(n_241), .B2(n_247), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_378), .A2(n_343), .B(n_320), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_378), .A2(n_330), .B1(n_331), .B2(n_336), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_369), .A2(n_327), .B1(n_266), .B2(n_341), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_340), .B1(n_352), .B2(n_337), .C(n_313), .Y(n_399) );
AO22x1_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_357), .B1(n_338), .B2(n_328), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_371), .A2(n_324), .B1(n_328), .B2(n_312), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_377), .B(n_334), .C(n_350), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_384), .A2(n_334), .B1(n_124), .B2(n_123), .C(n_99), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_384), .A2(n_369), .B1(n_383), .B2(n_372), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_324), .B1(n_266), .B2(n_355), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_366), .A2(n_93), .B(n_88), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_361), .A2(n_305), .B1(n_309), .B2(n_315), .C(n_321), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
NOR2xp67_ASAP7_75t_L g411 ( .A(n_386), .B(n_310), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_395), .A2(n_312), .B1(n_353), .B2(n_347), .Y(n_413) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_370), .A2(n_347), .B(n_359), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_386), .A2(n_345), .B1(n_359), .B2(n_325), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_376), .A2(n_329), .B1(n_325), .B2(n_359), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_380), .A2(n_377), .B(n_362), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_379), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_385), .B(n_325), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_375), .B(n_345), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_385), .B(n_329), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_375), .B(n_314), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_419), .B(n_393), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_401), .B(n_389), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_421), .B(n_389), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_417), .A2(n_362), .B(n_387), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_419), .B(n_363), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_399), .B(n_363), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_417), .A2(n_387), .B(n_367), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_398), .A2(n_368), .B1(n_392), .B2(n_365), .Y(n_432) );
AOI222xp33_ASAP7_75t_L g433 ( .A1(n_405), .A2(n_390), .B1(n_363), .B2(n_365), .C1(n_381), .C2(n_373), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_397), .A2(n_367), .B1(n_394), .B2(n_388), .C(n_365), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_407), .A2(n_391), .B(n_93), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_406), .B(n_391), .C(n_390), .Y(n_436) );
OAI33xp33_ASAP7_75t_L g437 ( .A1(n_401), .A2(n_120), .A3(n_99), .B1(n_100), .B2(n_106), .B3(n_123), .Y(n_437) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_409), .A2(n_157), .B(n_117), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_404), .A2(n_390), .B1(n_388), .B2(n_120), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_421), .B(n_388), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_396), .A2(n_117), .B(n_106), .Y(n_441) );
XNOR2xp5_ASAP7_75t_L g442 ( .A(n_412), .B(n_388), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_412), .A2(n_116), .B1(n_109), .B2(n_100), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_402), .B(n_109), .C(n_116), .D(n_158), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_408), .A2(n_174), .B1(n_157), .B2(n_202), .C(n_200), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_403), .A2(n_329), .B1(n_202), .B2(n_274), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_411), .A2(n_314), .B1(n_247), .B2(n_295), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_410), .A2(n_157), .B(n_206), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_418), .B(n_9), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_418), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
AO31x2_ASAP7_75t_L g454 ( .A1(n_422), .A2(n_284), .A3(n_296), .B(n_281), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_422), .A2(n_360), .B1(n_294), .B2(n_261), .Y(n_455) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_413), .A2(n_174), .B(n_132), .C(n_140), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_424), .A2(n_329), .B1(n_257), .B2(n_261), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_423), .B(n_274), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_450), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_450), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_450), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_440), .B(n_407), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_443), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_440), .B(n_407), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_427), .B(n_411), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_427), .B(n_423), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_443), .B(n_420), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_454), .Y(n_469) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_426), .B(n_416), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_452), .B(n_420), .Y(n_471) );
NOR3xp33_ASAP7_75t_SL g472 ( .A(n_444), .B(n_415), .C(n_414), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_444), .B(n_400), .C(n_222), .Y(n_473) );
OAI31xp33_ASAP7_75t_SL g474 ( .A1(n_432), .A2(n_400), .A3(n_10), .B(n_11), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_453), .Y(n_476) );
OAI33xp33_ASAP7_75t_L g477 ( .A1(n_425), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_13), .B3(n_14), .Y(n_477) );
INVx6_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_454), .Y(n_479) );
OAI31xp33_ASAP7_75t_L g480 ( .A1(n_439), .A2(n_13), .A3(n_14), .B(n_15), .Y(n_480) );
OAI211xp5_ASAP7_75t_SL g481 ( .A1(n_441), .A2(n_233), .B(n_222), .C(n_229), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_441), .A2(n_174), .B1(n_132), .B2(n_140), .C(n_171), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g483 ( .A(n_456), .B(n_76), .Y(n_483) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_442), .A2(n_16), .B1(n_17), .B2(n_18), .C(n_20), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_451), .B(n_17), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_433), .A2(n_329), .B1(n_174), .B2(n_130), .Y(n_488) );
AND3x1_ASAP7_75t_L g489 ( .A(n_451), .B(n_18), .C(n_20), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_430), .B(n_21), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_433), .B(n_23), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_436), .A2(n_174), .B1(n_130), .B2(n_132), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_458), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_454), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_442), .B(n_130), .Y(n_495) );
OAI221xp5_ASAP7_75t_SL g496 ( .A1(n_445), .A2(n_257), .B1(n_272), .B2(n_284), .C(n_281), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_458), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_428), .B(n_171), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_428), .B(n_171), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_454), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_454), .B(n_171), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_431), .B(n_171), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_436), .A2(n_272), .B1(n_140), .B2(n_132), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_431), .B(n_171), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_489), .B(n_448), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_462), .B(n_435), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_476), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_467), .B(n_431), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_474), .A2(n_445), .B(n_458), .C(n_434), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_461), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_462), .B(n_431), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_475), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_438), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_459), .B(n_438), .Y(n_518) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_489), .B(n_438), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_463), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_462), .B(n_435), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_484), .A2(n_437), .B1(n_446), .B2(n_435), .C(n_140), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_449), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_487), .B(n_457), .Y(n_525) );
OAI211xp5_ASAP7_75t_SL g526 ( .A1(n_472), .A2(n_447), .B(n_455), .C(n_229), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_463), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_463), .Y(n_528) );
AOI33xp33_ASAP7_75t_L g529 ( .A1(n_488), .A2(n_233), .A3(n_296), .B1(n_276), .B2(n_303), .B3(n_140), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_464), .B(n_449), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_471), .B(n_449), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_477), .B(n_303), .C(n_276), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_460), .Y(n_533) );
AND4x1_ASAP7_75t_L g534 ( .A(n_480), .B(n_25), .C(n_27), .D(n_30), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_464), .B(n_140), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_471), .B(n_132), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_460), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_464), .B(n_132), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_460), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_485), .B(n_33), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_494), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_464), .B(n_34), .Y(n_542) );
OAI211xp5_ASAP7_75t_SL g543 ( .A1(n_491), .A2(n_43), .B(n_46), .C(n_47), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_500), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_500), .B(n_49), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_468), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_468), .B(n_50), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_465), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_502), .B(n_51), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_469), .B(n_52), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_495), .B(n_55), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_478), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_495), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_486), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_493), .B(n_58), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_479), .B(n_60), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_490), .A2(n_288), .B(n_68), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_493), .B(n_67), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_478), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_466), .B(n_69), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_546), .B(n_470), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
NOR2x1p5_ASAP7_75t_L g565 ( .A(n_554), .B(n_502), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_553), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
NOR4xp25_ASAP7_75t_L g569 ( .A(n_506), .B(n_496), .C(n_504), .D(n_497), .Y(n_569) );
OAI32xp33_ASAP7_75t_L g570 ( .A1(n_552), .A2(n_473), .A3(n_497), .B1(n_481), .B2(n_486), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_550), .B(n_483), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_546), .B(n_470), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_512), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_555), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_549), .B(n_479), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_541), .Y(n_576) );
OAI21xp33_ASAP7_75t_L g577 ( .A1(n_522), .A2(n_492), .B(n_502), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_525), .B(n_502), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_541), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_510), .B(n_501), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_511), .B(n_478), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_517), .Y(n_583) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_517), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_510), .B(n_486), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_519), .A2(n_480), .B(n_482), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_544), .B(n_501), .Y(n_587) );
AOI32xp33_ASAP7_75t_L g588 ( .A1(n_543), .A2(n_499), .A3(n_498), .B1(n_505), .B2(n_503), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_544), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_521), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_522), .B(n_505), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_521), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_555), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_550), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_536), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_531), .B(n_499), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_548), .B(n_498), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_548), .B(n_503), .Y(n_598) );
OA211x2_ASAP7_75t_L g599 ( .A1(n_523), .A2(n_72), .B(n_74), .C(n_78), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_513), .B(n_225), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_527), .B(n_225), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_513), .B(n_225), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_528), .B(n_225), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_539), .B(n_225), .Y(n_604) );
OAI31xp33_ASAP7_75t_L g605 ( .A1(n_550), .A2(n_210), .A3(n_226), .B(n_218), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_508), .B(n_212), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_520), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_520), .B(n_212), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_533), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_533), .B(n_212), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_537), .Y(n_611) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_542), .B(n_265), .Y(n_612) );
XNOR2x1_ASAP7_75t_L g613 ( .A(n_565), .B(n_552), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_573), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_567), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_583), .B(n_537), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_568), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_563), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_564), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_584), .B(n_535), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_591), .B(n_535), .Y(n_621) );
AND2x2_ASAP7_75t_SL g622 ( .A(n_612), .B(n_519), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_582), .B(n_540), .Y(n_623) );
XNOR2xp5_ASAP7_75t_L g624 ( .A(n_612), .B(n_534), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_566), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_576), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_580), .B(n_538), .Y(n_627) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_578), .Y(n_628) );
AOI211x1_ASAP7_75t_L g629 ( .A1(n_586), .A2(n_558), .B(n_557), .C(n_551), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_562), .A2(n_538), .B1(n_561), .B2(n_507), .Y(n_630) );
AO22x2_ASAP7_75t_L g631 ( .A1(n_575), .A2(n_507), .B1(n_530), .B2(n_524), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_589), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_578), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_590), .B(n_507), .Y(n_634) );
XNOR2xp5_ASAP7_75t_L g635 ( .A(n_572), .B(n_560), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_592), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_577), .A2(n_551), .B1(n_542), .B2(n_524), .C1(n_530), .C2(n_545), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_575), .B(n_514), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_569), .A2(n_514), .B(n_559), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_579), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_581), .Y(n_641) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_594), .B(n_559), .Y(n_642) );
XNOR2xp5_ASAP7_75t_L g643 ( .A(n_591), .B(n_547), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_570), .A2(n_532), .B1(n_526), .B2(n_556), .C(n_518), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_587), .Y(n_645) );
AOI32xp33_ASAP7_75t_L g646 ( .A1(n_594), .A2(n_556), .A3(n_518), .B1(n_529), .B2(n_288), .Y(n_646) );
XOR2x2_ASAP7_75t_L g647 ( .A(n_571), .B(n_288), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_607), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_581), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_571), .A2(n_212), .B1(n_218), .B2(n_265), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_611), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_595), .B(n_218), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_585), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_574), .Y(n_654) );
OAI21xp33_ASAP7_75t_SL g655 ( .A1(n_588), .A2(n_210), .B(n_226), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_598), .B(n_265), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_598), .B(n_280), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_600), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_593), .B(n_210), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_597), .A2(n_280), .B(n_295), .C(n_226), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_602), .A2(n_295), .B(n_280), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_605), .A2(n_226), .B(n_599), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_596), .A2(n_593), .B(n_609), .C(n_604), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_609), .B(n_606), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_608), .B(n_610), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_601), .A2(n_563), .B1(n_549), .B2(n_509), .C(n_582), .Y(n_666) );
XOR2x2_ASAP7_75t_L g667 ( .A(n_603), .B(n_184), .Y(n_667) );
XNOR2xp5_ASAP7_75t_L g668 ( .A(n_643), .B(n_667), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_639), .A2(n_615), .B(n_618), .C(n_614), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g670 ( .A1(n_623), .A2(n_666), .A3(n_641), .B1(n_640), .B2(n_649), .C1(n_653), .C2(n_622), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_624), .A2(n_637), .B(n_663), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_650), .B(n_613), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_631), .A2(n_637), .B1(n_638), .B2(n_635), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_629), .A2(n_655), .B(n_644), .C(n_630), .Y(n_674) );
XNOR2x1_ASAP7_75t_L g675 ( .A(n_631), .B(n_647), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_650), .A2(n_628), .B(n_642), .Y(n_676) );
NOR4xp25_ASAP7_75t_L g677 ( .A(n_641), .B(n_617), .C(n_646), .D(n_645), .Y(n_677) );
NOR3xp33_ASAP7_75t_SL g678 ( .A(n_662), .B(n_657), .C(n_656), .Y(n_678) );
AOI22x1_ASAP7_75t_L g679 ( .A1(n_633), .A2(n_621), .B1(n_658), .B2(n_665), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_616), .A2(n_620), .B(n_634), .Y(n_680) );
NAND5xp2_ASAP7_75t_L g681 ( .A(n_670), .B(n_660), .C(n_657), .D(n_656), .E(n_661), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_679), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_677), .B(n_652), .C(n_636), .Y(n_683) );
AOI211x1_ASAP7_75t_L g684 ( .A1(n_671), .A2(n_616), .B(n_627), .C(n_625), .Y(n_684) );
AO22x2_ASAP7_75t_L g685 ( .A1(n_675), .A2(n_619), .B1(n_626), .B2(n_632), .Y(n_685) );
XOR2xp5_ASAP7_75t_L g686 ( .A(n_668), .B(n_627), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_680), .B(n_648), .Y(n_687) );
NAND4xp75_ASAP7_75t_L g688 ( .A(n_672), .B(n_664), .C(n_651), .D(n_659), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_682), .A2(n_673), .B1(n_676), .B2(n_687), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_685), .B(n_676), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_684), .B(n_683), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_685), .A2(n_669), .B1(n_674), .B2(n_678), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_689), .A2(n_688), .B1(n_686), .B2(n_681), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_690), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_691), .B(n_654), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_695), .Y(n_696) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_693), .B(n_692), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_696), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_698), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_699), .B(n_697), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_697), .B(n_694), .Y(n_701) );
endmodule