module fake_jpeg_31000_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_27),
.B(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_96),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_17),
.B(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_97),
.Y(n_126)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_74),
.Y(n_161)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_101),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_102),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_105),
.Y(n_129)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_106),
.Y(n_143)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_107),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_114),
.A2(n_26),
.B1(n_34),
.B2(n_49),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_24),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_115),
.B(n_136),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_36),
.B1(n_38),
.B2(n_24),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_116),
.A2(n_33),
.B1(n_22),
.B2(n_41),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_19),
.B1(n_51),
.B2(n_35),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_120),
.A2(n_121),
.B1(n_34),
.B2(n_49),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_54),
.A2(n_19),
.B1(n_51),
.B2(n_35),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_38),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_31),
.B(n_50),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_137),
.B(n_166),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_55),
.A2(n_36),
.B1(n_51),
.B2(n_44),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_149),
.B1(n_42),
.B2(n_22),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_80),
.B(n_46),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_57),
.A2(n_37),
.B1(n_46),
.B2(n_45),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_81),
.B(n_17),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_92),
.B(n_45),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_44),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_93),
.A2(n_26),
.B1(n_19),
.B2(n_39),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_59),
.B(n_39),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_94),
.B(n_37),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_173),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_189),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_112),
.A2(n_42),
.B(n_35),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_175),
.A2(n_210),
.B(n_15),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_176),
.B(n_184),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_178),
.B1(n_133),
.B2(n_156),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_126),
.B(n_42),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_179),
.B(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_183),
.A2(n_187),
.B1(n_216),
.B2(n_221),
.Y(n_258)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_161),
.Y(n_185)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_53),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_194),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_73),
.B1(n_65),
.B2(n_67),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_130),
.B(n_33),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_191),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_192),
.B(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_113),
.B(n_41),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_111),
.A2(n_124),
.B1(n_163),
.B2(n_117),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_198),
.A2(n_199),
.B1(n_215),
.B2(n_217),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_117),
.A2(n_33),
.B1(n_22),
.B2(n_83),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_53),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_209),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_144),
.B(n_108),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_5),
.B(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_34),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_49),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_152),
.B(n_154),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_213),
.B(n_220),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_109),
.Y(n_214)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_125),
.A2(n_86),
.B1(n_77),
.B2(n_78),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_120),
.A2(n_106),
.B1(n_102),
.B2(n_99),
.Y(n_216)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_114),
.A2(n_79),
.B1(n_63),
.B2(n_97),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_110),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_205),
.B(n_221),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_186),
.A2(n_146),
.B1(n_165),
.B2(n_95),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_236),
.A2(n_240),
.B1(n_244),
.B2(n_251),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_248),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_146),
.B1(n_165),
.B2(n_133),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_191),
.A2(n_139),
.B1(n_131),
.B2(n_160),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_213),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_179),
.A2(n_139),
.B1(n_160),
.B2(n_148),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_185),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_201),
.A2(n_168),
.B1(n_119),
.B2(n_123),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_217),
.B1(n_223),
.B2(n_190),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_182),
.B(n_181),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_181),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_182),
.A2(n_201),
.B(n_205),
.C(n_193),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_175),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_263),
.B(n_289),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_264),
.A2(n_268),
.B(n_254),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_216),
.B1(n_205),
.B2(n_187),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_265),
.A2(n_274),
.B1(n_293),
.B2(n_225),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_224),
.A2(n_192),
.B1(n_196),
.B2(n_204),
.Y(n_268)
);

XOR2x2_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_194),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_286),
.C(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_272),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_224),
.A2(n_209),
.B1(n_183),
.B2(n_172),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_279),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_231),
.B(n_193),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_276),
.B(n_231),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_188),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_278),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_282),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_230),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_228),
.A2(n_178),
.B(n_210),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_239),
.B(n_246),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_202),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_284),
.B(n_152),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_212),
.B1(n_127),
.B2(n_123),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_285),
.A2(n_287),
.B1(n_236),
.B2(n_255),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_180),
.C(n_208),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_119),
.B1(n_127),
.B2(n_142),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_226),
.B(n_176),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_291),
.B(n_292),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_195),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_233),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_281),
.B1(n_264),
.B2(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_302),
.B1(n_315),
.B2(n_285),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_300),
.A2(n_304),
.B(n_314),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_303),
.B(n_277),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_227),
.B1(n_243),
.B2(n_259),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_305),
.A2(n_290),
.B1(n_268),
.B2(n_293),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_246),
.B(n_237),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_307),
.A2(n_324),
.B(n_266),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_310),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_248),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_262),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_317),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_321),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_265),
.A2(n_240),
.B1(n_243),
.B2(n_245),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_245),
.Y(n_317)
);

AO21x2_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_227),
.B(n_253),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_291),
.B1(n_278),
.B2(n_272),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_288),
.B(n_249),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_323),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_269),
.A2(n_261),
.B(n_232),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_325),
.A2(n_333),
.B1(n_342),
.B2(n_354),
.Y(n_362)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_331),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_270),
.C(n_286),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_332),
.C(n_337),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_330),
.A2(n_300),
.B(n_295),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_322),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_270),
.C(n_286),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_265),
.B1(n_290),
.B2(n_274),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_273),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_310),
.C(n_317),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_322),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_338),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_263),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_339),
.B(n_351),
.Y(n_367)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_346),
.B1(n_318),
.B2(n_298),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_341),
.A2(n_345),
.B1(n_347),
.B2(n_320),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_296),
.A2(n_267),
.B1(n_271),
.B2(n_294),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_297),
.B(n_276),
.Y(n_343)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_318),
.Y(n_381)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_305),
.A2(n_292),
.B1(n_280),
.B2(n_252),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_261),
.C(n_238),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_324),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_242),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_184),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_309),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_315),
.A2(n_280),
.B1(n_252),
.B2(n_241),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_341),
.A2(n_312),
.B1(n_301),
.B2(n_314),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_358),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_356),
.A2(n_366),
.B1(n_379),
.B2(n_382),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_360),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_297),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g411 ( 
.A(n_363),
.B(n_380),
.CI(n_256),
.CON(n_411),
.SN(n_411)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_330),
.A2(n_295),
.B(n_312),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_369),
.B(n_370),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_345),
.A2(n_323),
.B1(n_320),
.B2(n_305),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_320),
.B(n_308),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_349),
.A2(n_304),
.B(n_308),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_336),
.A2(n_347),
.B(n_327),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_371),
.B(n_375),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_374),
.A2(n_346),
.B1(n_335),
.B2(n_333),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_336),
.A2(n_320),
.B(n_303),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_316),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_384),
.C(n_385),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_325),
.A2(n_320),
.B1(n_299),
.B2(n_298),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_377),
.A2(n_369),
.B1(n_368),
.B2(n_338),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_320),
.B1(n_299),
.B2(n_298),
.Y(n_379)
);

XOR2x1_ASAP7_75t_SL g380 ( 
.A(n_352),
.B(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_331),
.A2(n_241),
.B1(n_223),
.B2(n_214),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_343),
.A2(n_232),
.B(n_238),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_354),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_197),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_218),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_386),
.A2(n_393),
.B1(n_395),
.B2(n_404),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_389),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_348),
.Y(n_388)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_348),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_392),
.A2(n_409),
.B1(n_385),
.B2(n_365),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_362),
.A2(n_353),
.B1(n_342),
.B2(n_326),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_377),
.B1(n_368),
.B2(n_357),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_371),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_401),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_364),
.B(n_344),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_334),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_256),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_350),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_403),
.B(n_405),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_380),
.A2(n_337),
.B1(n_214),
.B2(n_219),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_242),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_356),
.A2(n_366),
.B1(n_355),
.B2(n_379),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_408),
.B1(n_413),
.B2(n_414),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_358),
.A2(n_370),
.B1(n_382),
.B2(n_378),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_411),
.B(n_256),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_360),
.A2(n_219),
.B1(n_260),
.B2(n_189),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_383),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_376),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_424),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_417),
.A2(n_419),
.B1(n_393),
.B2(n_404),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_378),
.C(n_234),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_423),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_260),
.B1(n_204),
.B2(n_222),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_397),
.Y(n_420)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_234),
.C(n_260),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_220),
.B(n_206),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_426),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_409),
.C(n_390),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_207),
.C(n_135),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_429),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_135),
.C(n_151),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_431),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_118),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_406),
.A2(n_142),
.B1(n_168),
.B2(n_173),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_435),
.A2(n_422),
.B1(n_437),
.B2(n_431),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_413),
.Y(n_442)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_421),
.Y(n_441)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_442),
.B(n_151),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_454),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_415),
.A2(n_394),
.B1(n_400),
.B2(n_398),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_447),
.B1(n_452),
.B2(n_457),
.Y(n_474)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_428),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_451),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_398),
.B1(n_410),
.B2(n_407),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_427),
.A2(n_386),
.B1(n_388),
.B2(n_396),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_448),
.A2(n_450),
.B1(n_11),
.B2(n_15),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_417),
.A2(n_399),
.B1(n_402),
.B2(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_434),
.A2(n_411),
.B1(n_173),
.B2(n_217),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_411),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_456),
.Y(n_465)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_418),
.C(n_423),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_459),
.B(n_464),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_455),
.Y(n_460)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_460),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_416),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_466),
.Y(n_489)
);

OAI321xp33_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_424),
.A3(n_419),
.B1(n_425),
.B2(n_430),
.C(n_429),
.Y(n_463)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_436),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_467),
.A2(n_473),
.B1(n_7),
.B2(n_13),
.Y(n_483)
);

AOI21xp33_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_148),
.B(n_12),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_468),
.A2(n_10),
.B(n_14),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_470),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_162),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_444),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_440),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_452),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_50),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_440),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_472),
.Y(n_476)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_483),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_467),
.A2(n_453),
.B(n_442),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_479),
.A2(n_2),
.B(n_3),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_487),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_439),
.C(n_50),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_30),
.C(n_50),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_488),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_473),
.A2(n_5),
.B1(n_12),
.B2(n_7),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_486),
.A2(n_474),
.B1(n_461),
.B2(n_4),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_4),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_498),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_477),
.B1(n_479),
.B2(n_483),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_494),
.B(n_495),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_490),
.A2(n_462),
.B(n_470),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_484),
.A2(n_30),
.B(n_50),
.Y(n_496)
);

MAJx2_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_486),
.C(n_50),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_477),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_2),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_2),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_30),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_489),
.C(n_481),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_503),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_510),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_493),
.A2(n_497),
.B(n_500),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_508),
.Y(n_512)
);

AOI21xp33_ASAP7_75t_L g509 ( 
.A1(n_494),
.A2(n_489),
.B(n_43),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_509),
.A2(n_501),
.B(n_504),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_514),
.B(n_515),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_491),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_506),
.C(n_491),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_517),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_513),
.A2(n_502),
.B(n_498),
.Y(n_518)
);

NOR3xp33_ASAP7_75t_SL g520 ( 
.A(n_518),
.B(n_511),
.C(n_30),
.Y(n_520)
);

AOI322xp5_ASAP7_75t_L g521 ( 
.A1(n_520),
.A2(n_2),
.A3(n_3),
.B1(n_30),
.B2(n_43),
.C1(n_516),
.C2(n_519),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_3),
.Y(n_522)
);

AOI21x1_ASAP7_75t_SL g523 ( 
.A1(n_522),
.A2(n_30),
.B(n_43),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_43),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_43),
.Y(n_525)
);


endmodule