module fake_jpeg_80_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_53),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_47),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_37),
.C(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_62),
.B(n_87),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_20),
.B1(n_21),
.B2(n_36),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_64),
.A2(n_71),
.B1(n_91),
.B2(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_20),
.B1(n_21),
.B2(n_36),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_36),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_6),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_35),
.B1(n_29),
.B2(n_27),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_75),
.A2(n_82),
.B1(n_12),
.B2(n_68),
.Y(n_135)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_35),
.B1(n_27),
.B2(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_97),
.B1(n_64),
.B2(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_35),
.B1(n_29),
.B2(n_17),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_2),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_30),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_42),
.A2(n_30),
.B1(n_15),
.B2(n_33),
.Y(n_91)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_37),
.B1(n_34),
.B2(n_33),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_101),
.Y(n_114)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_105),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_10),
.C(n_12),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_43),
.A2(n_15),
.B1(n_31),
.B2(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_31),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_8),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_15),
.B1(n_3),
.B2(n_5),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_135),
.B1(n_92),
.B2(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_14),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_117),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_63),
.B1(n_88),
.B2(n_93),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_2),
.C(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_136),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_14),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_129),
.B(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_87),
.B(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_98),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_104),
.B1(n_78),
.B2(n_76),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_147),
.B1(n_149),
.B2(n_161),
.Y(n_181)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_73),
.B(n_81),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_129),
.B(n_124),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_146),
.A2(n_138),
.B1(n_121),
.B2(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_69),
.B1(n_106),
.B2(n_61),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_61),
.B1(n_106),
.B2(n_88),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_164),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_96),
.A3(n_100),
.B1(n_81),
.B2(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_86),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_86),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.Y(n_183)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_114),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_123),
.B1(n_121),
.B2(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_110),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_133),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_160),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_185),
.B1(n_147),
.B2(n_140),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_187),
.B(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_120),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_121),
.B1(n_139),
.B2(n_132),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_121),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_191),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_139),
.B(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_118),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_118),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_151),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_144),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_177),
.B(n_158),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_197),
.B(n_213),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_143),
.B(n_171),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_148),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_207),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_205),
.B1(n_212),
.B2(n_178),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_141),
.B1(n_162),
.B2(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_174),
.B(n_187),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_149),
.B1(n_168),
.B2(n_154),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_142),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_191),
.C(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_220),
.C(n_225),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_204),
.B1(n_212),
.B2(n_206),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_223),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_181),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_194),
.B(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_200),
.C(n_197),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_194),
.C(n_193),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_180),
.C(n_175),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_180),
.B(n_188),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_207),
.B(n_206),
.Y(n_236)
);

BUFx12f_ASAP7_75t_SL g230 ( 
.A(n_229),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_236),
.B(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_221),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_205),
.B1(n_202),
.B2(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_228),
.C(n_225),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_229),
.B1(n_224),
.B2(n_216),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_231),
.B1(n_233),
.B2(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_219),
.C(n_214),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_235),
.C(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_234),
.C(n_239),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_241),
.B(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_236),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_261),
.B(n_205),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_241),
.B(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_248),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

A2O1A1O1Ixp25_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_251),
.B(n_255),
.C(n_246),
.D(n_205),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_203),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_203),
.Y(n_270)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.C(n_268),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_258),
.Y(n_272)
);


endmodule