module fake_ariane_2867_n_1858 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1858);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1858;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1759;
wire n_1557;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_99),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_36),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_40),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_34),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_90),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_87),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_70),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_138),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_22),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_177),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_115),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_116),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_96),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_34),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_67),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_54),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_104),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_9),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_23),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_91),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_98),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_88),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_4),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_10),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_38),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_66),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_56),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_65),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_78),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_16),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_22),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_95),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_113),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_39),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_101),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_64),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_106),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_62),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_62),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_9),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_137),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_14),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_134),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_21),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_136),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_160),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_125),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_49),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_85),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_167),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_111),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_144),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_123),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_79),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_151),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_121),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_66),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_83),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_14),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_122),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_126),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_77),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_139),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_158),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_46),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_71),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_19),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_39),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_49),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_174),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_156),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_26),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_112),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_127),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_119),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_76),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_37),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_114),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_75),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_154),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_5),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_53),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_135),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_3),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_20),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_86),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_19),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_124),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_18),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_29),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_170),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_93),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_27),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_41),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_163),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_25),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_142),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_7),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_100),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_2),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_43),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_57),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_44),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_58),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_110),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_152),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_146),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_44),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_68),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_74),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_60),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_27),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_54),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_21),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_63),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_65),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_33),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_153),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_52),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_118),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_59),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_3),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_131),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_58),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_171),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_37),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_73),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_81),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_145),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_150),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_108),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_157),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_42),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_45),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_109),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_159),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_191),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_341),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_227),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_185),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_265),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_185),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_186),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_186),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_182),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_188),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_188),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_189),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_225),
.B(n_0),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_320),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_199),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_248),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_190),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_203),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_204),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_192),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_213),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_193),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_209),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_183),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_192),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_194),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_194),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_207),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_279),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_216),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_292),
.B(n_0),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_210),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_217),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_210),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_215),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_215),
.Y(n_401)
);

BUFx2_ASAP7_75t_SL g402 ( 
.A(n_353),
.Y(n_402)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_234),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_222),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_222),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_236),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_238),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_228),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_227),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_243),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_244),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_315),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_247),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_225),
.B(n_1),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_253),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_257),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_262),
.B(n_1),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_262),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_270),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_228),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_214),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_245),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_304),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_245),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_275),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_323),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_250),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_260),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_267),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_227),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_362),
.B(n_181),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_283),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_267),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_288),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_353),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_289),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_291),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_269),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_213),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_353),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_269),
.B(n_2),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_319),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_319),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_293),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_227),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_296),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_319),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_272),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_308),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_272),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_277),
.B(n_5),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_313),
.Y(n_453)
);

INVx4_ASAP7_75t_R g454 ( 
.A(n_205),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_364),
.B(n_221),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_387),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_380),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_372),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_368),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_389),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_409),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_365),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_379),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_381),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_366),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_369),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_369),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_370),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_378),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_370),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_371),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_402),
.B(n_255),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_371),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_373),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_373),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_402),
.B(n_310),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_R g489 ( 
.A(n_383),
.B(n_187),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_384),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_375),
.A2(n_294),
.B(n_277),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_375),
.B(n_211),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_377),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_377),
.B(n_211),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_453),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_367),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_395),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_385),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_385),
.B(n_218),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_398),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_406),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_R g504 ( 
.A(n_407),
.B(n_316),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_390),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_391),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_391),
.B(n_218),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_410),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_411),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_367),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_393),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_392),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_397),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_442),
.A2(n_298),
.B(n_294),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_399),
.B(n_233),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_432),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_400),
.B(n_298),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_401),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_401),
.B(n_292),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_394),
.A2(n_360),
.B1(n_223),
.B2(n_226),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_412),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_376),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_415),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_408),
.B(n_233),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_491),
.A2(n_420),
.B1(n_422),
.B2(n_408),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_467),
.B(n_403),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_473),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_467),
.B(n_470),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_482),
.B(n_414),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_470),
.B(n_420),
.Y(n_540)
);

INVx4_ASAP7_75t_SL g541 ( 
.A(n_476),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_440),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_475),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_529),
.B(n_416),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_482),
.B(n_417),
.C(n_425),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_382),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_471),
.B(n_422),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_529),
.B(n_433),
.Y(n_549)
);

NAND3xp33_ASAP7_75t_L g550 ( 
.A(n_487),
.B(n_437),
.C(n_435),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_484),
.B(n_424),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_483),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_484),
.B(n_445),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_466),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_484),
.B(n_447),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_529),
.B(n_312),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_472),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_489),
.B(n_429),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_496),
.B(n_388),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_522),
.B(n_424),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_487),
.A2(n_452),
.B1(n_305),
.B2(n_451),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_522),
.B(n_427),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_522),
.B(n_427),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_472),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_522),
.B(n_428),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_485),
.B(n_428),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_486),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_526),
.B(n_396),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_488),
.B(n_430),
.Y(n_578)
);

BUFx4f_ASAP7_75t_L g579 ( 
.A(n_476),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_493),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_529),
.B(n_312),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_476),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_493),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_477),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_491),
.A2(n_451),
.B1(n_449),
.B2(n_430),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_512),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_477),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_513),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_529),
.B(n_314),
.Y(n_595)
);

INVx4_ASAP7_75t_SL g596 ( 
.A(n_477),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_504),
.A2(n_419),
.B1(n_438),
.B2(n_421),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_477),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_457),
.B(n_311),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_515),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_515),
.B(n_434),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_497),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_518),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_480),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_518),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_480),
.B(n_314),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_500),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_524),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_524),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_525),
.B(n_434),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_480),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_501),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

BUFx4f_ASAP7_75t_L g615 ( 
.A(n_480),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_523),
.B(n_331),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_528),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_480),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_528),
.B(n_439),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_491),
.A2(n_449),
.B1(n_439),
.B2(n_386),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_531),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_531),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_480),
.B(n_331),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_457),
.A2(n_223),
.B1(n_226),
.B2(n_230),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_475),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_460),
.A2(n_423),
.B1(n_426),
.B2(n_441),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_475),
.B(n_333),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_491),
.A2(n_311),
.B1(n_326),
.B2(n_327),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_511),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_510),
.B(n_436),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_498),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_498),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_478),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_523),
.B(n_198),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_523),
.B(n_202),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_489),
.B(n_443),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_498),
.B(n_503),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_498),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_498),
.B(n_333),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_527),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_498),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_491),
.A2(n_286),
.B1(n_280),
.B2(n_276),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_510),
.B(n_444),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_523),
.B(n_230),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_523),
.B(n_335),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_502),
.A2(n_448),
.B1(n_337),
.B2(n_322),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_502),
.B(n_232),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_498),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_481),
.B(n_335),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_481),
.B(n_346),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_503),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_514),
.B(n_354),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_533),
.A2(n_307),
.B1(n_276),
.B2(n_360),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_514),
.B(n_521),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_509),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_458),
.B(n_231),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_521),
.B(n_354),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_L g659 ( 
.A(n_530),
.B(n_231),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_503),
.B(n_357),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_503),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_503),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_468),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_533),
.A2(n_301),
.B1(n_261),
.B2(n_306),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_468),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_503),
.B(n_357),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_503),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_532),
.B(n_227),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_505),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_505),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_505),
.B(n_506),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_505),
.Y(n_672)
);

AND2x6_ASAP7_75t_L g673 ( 
.A(n_492),
.B(n_184),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_492),
.B(n_184),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_505),
.Y(n_675)
);

NOR2x1p5_ASAP7_75t_L g676 ( 
.A(n_463),
.B(n_251),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_504),
.A2(n_479),
.B1(n_458),
.B2(n_464),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_505),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_520),
.B(n_240),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_505),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_555),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_544),
.B(n_464),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_554),
.B(n_479),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_544),
.B(n_549),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_554),
.B(n_557),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_SL g687 ( 
.A(n_613),
.B(n_549),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_557),
.B(n_492),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_539),
.B(n_519),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_539),
.B(n_520),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_566),
.B(n_494),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_566),
.B(n_568),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_534),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_559),
.B(n_506),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_559),
.A2(n_533),
.B1(n_517),
.B2(n_507),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_537),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_581),
.B(n_506),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_550),
.B(n_519),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_643),
.A2(n_533),
.B1(n_516),
.B2(n_506),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_555),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_568),
.B(n_494),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_553),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_677),
.B(n_519),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_672),
.A2(n_516),
.B(n_519),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_679),
.B(n_494),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_599),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_643),
.A2(n_533),
.B1(n_516),
.B2(n_506),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_581),
.B(n_506),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_602),
.B(n_469),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_564),
.B(n_461),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_563),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_679),
.B(n_499),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_629),
.A2(n_506),
.B1(n_517),
.B2(n_507),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_573),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_595),
.B(n_536),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_555),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_599),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_542),
.B(n_461),
.Y(n_719)
);

INVx8_ASAP7_75t_L g720 ( 
.A(n_673),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_545),
.B(n_499),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_556),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_595),
.A2(n_517),
.B1(n_507),
.B2(n_499),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_519),
.B(n_456),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_546),
.B(n_338),
.C(n_334),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_536),
.B(n_567),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_572),
.A2(n_261),
.B(n_306),
.C(n_252),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_597),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_545),
.B(n_495),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_630),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_572),
.B(n_519),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_616),
.A2(n_646),
.B1(n_674),
.B2(n_673),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_574),
.A2(n_342),
.B1(n_345),
.B2(n_347),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_584),
.B(n_519),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_576),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_578),
.B(n_519),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_251),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_654),
.A2(n_239),
.B1(n_235),
.B2(n_328),
.C(n_327),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_580),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_558),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_538),
.B(n_350),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_585),
.B(n_252),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_673),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_543),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_588),
.B(n_280),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_555),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_628),
.A2(n_650),
.B(n_653),
.C(n_651),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_641),
.B(n_495),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_569),
.A2(n_328),
.B(n_348),
.C(n_343),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_591),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_607),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_614),
.B(n_286),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_656),
.B(n_352),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_593),
.B(n_301),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_594),
.B(n_307),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_600),
.B(n_324),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_648),
.B(n_324),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_638),
.A2(n_297),
.B(n_462),
.Y(n_758)
);

BUFx10_ASAP7_75t_L g759 ( 
.A(n_659),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_625),
.B(n_329),
.C(n_343),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_625),
.B(n_196),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_673),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_558),
.B(n_197),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_635),
.B(n_636),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_603),
.B(n_326),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_644),
.B(n_329),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_633),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_645),
.B(n_200),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_605),
.B(n_330),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_608),
.B(n_330),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_570),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_673),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_629),
.A2(n_664),
.B1(n_654),
.B2(n_542),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_645),
.B(n_201),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_582),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_609),
.A2(n_340),
.B1(n_348),
.B2(n_359),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_610),
.B(n_456),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_617),
.B(n_456),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_664),
.A2(n_340),
.B1(n_205),
.B2(n_336),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_622),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_623),
.B(n_206),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_540),
.B(n_456),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_655),
.A2(n_456),
.B(n_462),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_676),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_621),
.B(n_208),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_582),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_626),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_616),
.A2(n_336),
.B1(n_361),
.B2(n_281),
.Y(n_788)
);

BUFx5_ASAP7_75t_L g789 ( 
.A(n_674),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_SL g790 ( 
.A(n_647),
.B(n_219),
.C(n_212),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_633),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_583),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_631),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_548),
.B(n_551),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_542),
.A2(n_237),
.B1(n_249),
.B2(n_359),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_657),
.B(n_561),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_583),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_562),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_601),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_611),
.B(n_454),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_577),
.B(n_627),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_590),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_220),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_SL g804 ( 
.A1(n_577),
.A2(n_359),
.B1(n_249),
.B2(n_237),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_562),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_634),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_620),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_616),
.B(n_359),
.Y(n_808)
);

OAI221xp5_ASAP7_75t_L g809 ( 
.A1(n_577),
.A2(n_359),
.B1(n_224),
.B2(n_295),
.C(n_229),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_637),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_646),
.B(n_241),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_571),
.B(n_6),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_661),
.B(n_6),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_646),
.B(n_674),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_661),
.B(n_10),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_674),
.A2(n_468),
.B1(n_193),
.B2(n_273),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_646),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_590),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_674),
.B(n_242),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_612),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_628),
.A2(n_193),
.B1(n_273),
.B2(n_356),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_565),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_565),
.B(n_618),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_535),
.B(n_246),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_668),
.A2(n_299),
.B1(n_254),
.B2(n_256),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_535),
.B(n_258),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_619),
.B(n_11),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_650),
.A2(n_653),
.B(n_658),
.C(n_651),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_587),
.B(n_468),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_587),
.A2(n_300),
.B1(n_259),
.B2(n_263),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_658),
.B(n_264),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_619),
.B(n_266),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_666),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_606),
.B(n_468),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_579),
.B(n_268),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_606),
.A2(n_317),
.B1(n_271),
.B2(n_274),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_579),
.B(n_278),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_686),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_716),
.A2(n_638),
.B(n_678),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_716),
.B(n_592),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_690),
.B(n_633),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_773),
.A2(n_615),
.B1(n_598),
.B2(n_639),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_705),
.A2(n_649),
.B(n_652),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_692),
.A2(n_615),
.B(n_598),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_729),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_SL g846 ( 
.A(n_710),
.B(n_282),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_731),
.A2(n_680),
.B(n_667),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_748),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_720),
.B(n_624),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_689),
.A2(n_670),
.B(n_652),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_720),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_682),
.B(n_660),
.C(n_640),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_736),
.A2(n_649),
.B(n_642),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_693),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_747),
.A2(n_592),
.B(n_632),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_688),
.B(n_632),
.Y(n_856)
);

AO21x1_ASAP7_75t_L g857 ( 
.A1(n_684),
.A2(n_665),
.B(n_663),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_828),
.A2(n_639),
.B(n_586),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_829),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_685),
.A2(n_455),
.B(n_462),
.C(n_15),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_730),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_720),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_696),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_SL g864 ( 
.A1(n_684),
.A2(n_455),
.B(n_596),
.C(n_541),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_690),
.A2(n_675),
.B(n_669),
.C(n_662),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_698),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_764),
.B(n_633),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_764),
.B(n_662),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_703),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_772),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_724),
.A2(n_455),
.B(n_596),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_711),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_728),
.B(n_662),
.Y(n_873)
);

BUFx4f_ASAP7_75t_L g874 ( 
.A(n_719),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_794),
.A2(n_823),
.B(n_713),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_712),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_760),
.A2(n_675),
.B(n_669),
.C(n_662),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_715),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_694),
.A2(n_575),
.B(n_604),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_741),
.B(n_706),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_741),
.B(n_669),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_794),
.A2(n_675),
.B(n_669),
.Y(n_882)
);

BUFx12f_ASAP7_75t_L g883 ( 
.A(n_740),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_812),
.A2(n_675),
.B(n_604),
.C(n_589),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_762),
.B(n_575),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_691),
.A2(n_604),
.B1(n_589),
.B2(n_586),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_735),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_812),
.A2(n_604),
.B(n_589),
.C(n_586),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_759),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_823),
.A2(n_702),
.B(n_782),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_L g891 ( 
.A1(n_752),
.A2(n_287),
.B(n_285),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_732),
.A2(n_589),
.B1(n_586),
.B2(n_575),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_760),
.A2(n_596),
.B1(n_541),
.B2(n_575),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_799),
.B(n_541),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_817),
.A2(n_325),
.B1(n_284),
.B2(n_290),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_807),
.B(n_302),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_722),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_762),
.B(n_468),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_699),
.A2(n_465),
.B(n_459),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_683),
.B(n_358),
.C(n_355),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_782),
.A2(n_321),
.B(n_303),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_707),
.B(n_718),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_SL g903 ( 
.A(n_751),
.B(n_351),
.C(n_349),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_783),
.A2(n_318),
.B(n_309),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_832),
.A2(n_344),
.B(n_332),
.Y(n_905)
);

AO22x1_ASAP7_75t_L g906 ( 
.A1(n_801),
.A2(n_273),
.B1(n_193),
.B2(n_17),
.Y(n_906)
);

BUFx12f_ASAP7_75t_L g907 ( 
.A(n_759),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_694),
.A2(n_465),
.B(n_459),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_697),
.A2(n_465),
.B(n_459),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_721),
.B(n_12),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_727),
.A2(n_13),
.B(n_17),
.C(n_20),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_810),
.B(n_24),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_709),
.A2(n_778),
.B(n_777),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_777),
.A2(n_465),
.B(n_459),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_817),
.A2(n_465),
.B1(n_26),
.B2(n_28),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_778),
.A2(n_179),
.B(n_176),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_835),
.A2(n_175),
.B(n_172),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_837),
.A2(n_166),
.B(n_164),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_739),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_726),
.B(n_25),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_772),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_804),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_793),
.B(n_751),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_719),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_719),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_723),
.B(n_31),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_737),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_798),
.A2(n_162),
.B(n_161),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_795),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_750),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_795),
.B(n_35),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_798),
.A2(n_155),
.B(n_143),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_805),
.A2(n_133),
.B(n_132),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_780),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_L g935 ( 
.A(n_762),
.B(n_789),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_787),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_806),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_833),
.A2(n_128),
.B(n_117),
.Y(n_938)
);

O2A1O1Ixp5_ASAP7_75t_L g939 ( 
.A1(n_831),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_796),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_805),
.A2(n_97),
.B(n_84),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_768),
.B(n_47),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_822),
.A2(n_48),
.B(n_50),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_695),
.B(n_50),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_775),
.A2(n_51),
.B(n_52),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_743),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_714),
.B(n_59),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_786),
.A2(n_61),
.B(n_63),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_774),
.B(n_64),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_792),
.A2(n_797),
.B(n_802),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_813),
.A2(n_815),
.B(n_827),
.C(n_809),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_704),
.A2(n_814),
.B(n_824),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_818),
.A2(n_820),
.B(n_700),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_781),
.A2(n_734),
.B(n_808),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_700),
.A2(n_708),
.B(n_758),
.Y(n_955)
);

AOI33xp33_ASAP7_75t_L g956 ( 
.A1(n_784),
.A2(n_779),
.A3(n_749),
.B1(n_821),
.B2(n_714),
.B3(n_757),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_687),
.B(n_753),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_827),
.A2(n_815),
.B(n_813),
.C(n_765),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_762),
.B(n_789),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_725),
.A2(n_779),
.B(n_788),
.C(n_761),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_708),
.A2(n_826),
.B(n_834),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_742),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_771),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_745),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_681),
.A2(n_701),
.B(n_717),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_754),
.B(n_769),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_681),
.A2(n_701),
.B(n_717),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_738),
.A2(n_725),
.B(n_790),
.C(n_821),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_743),
.A2(n_772),
.B1(n_785),
.B2(n_803),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_762),
.B(n_789),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_755),
.A2(n_756),
.B(n_770),
.C(n_776),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_800),
.B(n_744),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_681),
.A2(n_701),
.B(n_717),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_744),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_811),
.A2(n_819),
.B(n_766),
.C(n_763),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_681),
.A2(n_701),
.B(n_717),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_767),
.A2(n_816),
.B1(n_746),
.B2(n_791),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_830),
.B(n_789),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_733),
.B(n_825),
.C(n_836),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_816),
.A2(n_789),
.B(n_746),
.C(n_791),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_767),
.B(n_746),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_791),
.A2(n_828),
.B(n_747),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_767),
.A2(n_692),
.B(n_731),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_693),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_689),
.A2(n_705),
.B(n_638),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_693),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_716),
.A2(n_773),
.B1(n_692),
.B2(n_685),
.Y(n_987)
);

NOR2xp67_ASAP7_75t_L g988 ( 
.A(n_751),
.B(n_613),
.Y(n_988)
);

CKINVDCx10_ASAP7_75t_R g989 ( 
.A(n_719),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_716),
.A2(n_685),
.B(n_581),
.C(n_595),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_730),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_747),
.A2(n_828),
.B(n_692),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_692),
.A2(n_736),
.B(n_731),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_692),
.A2(n_736),
.B(n_731),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_692),
.A2(n_736),
.B(n_731),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_716),
.B(n_688),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_716),
.B(n_688),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_720),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_716),
.B(n_688),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_L g1000 ( 
.A1(n_685),
.A2(n_684),
.B(n_581),
.C(n_595),
.Y(n_1000)
);

BUFx2_ASAP7_75t_SL g1001 ( 
.A(n_710),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_716),
.A2(n_773),
.B1(n_692),
.B2(n_685),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_716),
.B(n_688),
.Y(n_1003)
);

O2A1O1Ixp5_ASAP7_75t_L g1004 ( 
.A1(n_685),
.A2(n_684),
.B(n_581),
.C(n_595),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_690),
.B(n_684),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_716),
.B(n_688),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_716),
.A2(n_685),
.B(n_581),
.C(n_595),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_716),
.B(n_688),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_693),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_716),
.B(n_688),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_748),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_716),
.B(n_685),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_689),
.A2(n_705),
.B(n_638),
.Y(n_1013)
);

OAI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_716),
.A2(n_738),
.B1(n_577),
.B2(n_482),
.Y(n_1014)
);

AO22x1_ASAP7_75t_L g1015 ( 
.A1(n_760),
.A2(n_380),
.B1(n_460),
.B2(n_602),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_1012),
.A2(n_990),
.B(n_1007),
.C(n_920),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_875),
.A2(n_997),
.B(n_996),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_848),
.B(n_1011),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_1012),
.A2(n_920),
.B(n_987),
.C(n_1002),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_SL g1020 ( 
.A1(n_980),
.A2(n_955),
.B(n_999),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_992),
.A2(n_958),
.B(n_890),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_958),
.A2(n_951),
.B(n_982),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_993),
.A2(n_995),
.B(n_994),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_922),
.B(n_968),
.C(n_979),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1003),
.A2(n_1008),
.B(n_1006),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_862),
.B(n_870),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_845),
.B(n_988),
.Y(n_1028)
);

OA22x2_ASAP7_75t_L g1029 ( 
.A1(n_872),
.A2(n_845),
.B1(n_912),
.B2(n_924),
.Y(n_1029)
);

AND3x2_ASAP7_75t_L g1030 ( 
.A(n_872),
.B(n_861),
.C(n_846),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1000),
.A2(n_1004),
.B(n_880),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_871),
.A2(n_853),
.B(n_899),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1010),
.A2(n_913),
.B(n_881),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_850),
.A2(n_952),
.B(n_855),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_840),
.A2(n_868),
.B(n_867),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_882),
.A2(n_858),
.B(n_844),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_847),
.A2(n_909),
.B(n_908),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_897),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_857),
.A2(n_839),
.A3(n_969),
.B(n_865),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1005),
.A2(n_856),
.B(n_971),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_959),
.A2(n_970),
.B(n_953),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1005),
.A2(n_914),
.B(n_978),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_859),
.B(n_873),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_838),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_959),
.A2(n_967),
.B(n_973),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_965),
.A2(n_976),
.B(n_898),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1014),
.B(n_923),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_935),
.A2(n_966),
.B(n_884),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_971),
.A2(n_910),
.B(n_954),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_968),
.A2(n_960),
.B(n_942),
.C(n_949),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_862),
.B(n_870),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1014),
.A2(n_926),
.B1(n_944),
.B2(n_947),
.Y(n_1052)
);

AOI211x1_ASAP7_75t_L g1053 ( 
.A1(n_929),
.A2(n_878),
.B(n_887),
.C(n_1009),
.Y(n_1053)
);

CKINVDCx8_ASAP7_75t_R g1054 ( 
.A(n_989),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_874),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_870),
.B(n_998),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_859),
.B(n_962),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1015),
.B(n_940),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_841),
.A2(n_852),
.B(n_842),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_942),
.A2(n_949),
.B(n_979),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_977),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_854),
.A2(n_930),
.B1(n_984),
.B2(n_876),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_950),
.A2(n_879),
.B(n_885),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_912),
.B(n_874),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_964),
.B(n_902),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_991),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_885),
.A2(n_961),
.B(n_938),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_861),
.B(n_925),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_863),
.B(n_866),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_889),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_902),
.B(n_956),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_870),
.Y(n_1072)
);

BUFx8_ASAP7_75t_L g1073 ( 
.A(n_883),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_869),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_886),
.A2(n_981),
.B(n_916),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_919),
.A2(n_934),
.B1(n_986),
.B2(n_936),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_888),
.A2(n_937),
.B(n_975),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_877),
.A2(n_864),
.B(n_860),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_972),
.A2(n_892),
.B(n_906),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_907),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_957),
.A2(n_900),
.B1(n_940),
.B2(n_931),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_891),
.B(n_896),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_998),
.B(n_851),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_900),
.B(n_974),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_963),
.B(n_851),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_921),
.B(n_998),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_998),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_928),
.A2(n_941),
.B(n_932),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_911),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_921),
.B(n_894),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_849),
.B(n_893),
.Y(n_1091)
);

BUFx10_ASAP7_75t_L g1092 ( 
.A(n_849),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_901),
.A2(n_939),
.B(n_905),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_849),
.B(n_864),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_904),
.A2(n_917),
.B(n_918),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_903),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_943),
.A2(n_945),
.B(n_948),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_933),
.A2(n_915),
.B(n_946),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_895),
.B(n_927),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_996),
.B(n_997),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_872),
.B(n_728),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_862),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_983),
.A2(n_899),
.B(n_993),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1012),
.A2(n_716),
.B(n_690),
.C(n_990),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_SL g1108 ( 
.A1(n_987),
.A2(n_1002),
.B(n_982),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_996),
.B(n_997),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1111)
);

INVx8_ASAP7_75t_L g1112 ( 
.A(n_889),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1012),
.A2(n_716),
.B(n_690),
.C(n_990),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_838),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_996),
.B(n_997),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_838),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_870),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1000),
.A2(n_1004),
.B(n_716),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_845),
.B(n_677),
.Y(n_1122)
);

AND2x2_ASAP7_75t_SL g1123 ( 
.A(n_874),
.B(n_773),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_872),
.B(n_728),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_SL g1126 ( 
.A1(n_980),
.A2(n_743),
.B(n_955),
.Y(n_1126)
);

INVx3_ASAP7_75t_SL g1127 ( 
.A(n_897),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1012),
.A2(n_716),
.B(n_690),
.C(n_990),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_1001),
.B(n_584),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_874),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_983),
.A2(n_899),
.B(n_993),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_872),
.B(n_728),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_983),
.A2(n_899),
.B(n_993),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_992),
.A2(n_875),
.B(n_958),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_996),
.B(n_997),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_996),
.B(n_997),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_870),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_996),
.B(n_997),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_843),
.A2(n_1013),
.B(n_985),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_996),
.B(n_997),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1014),
.A2(n_542),
.B1(n_487),
.B2(n_482),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_SL g1144 ( 
.A1(n_987),
.A2(n_1002),
.B1(n_716),
.B2(n_1014),
.C(n_793),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_996),
.B(n_997),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_992),
.A2(n_875),
.B(n_958),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_992),
.A2(n_875),
.B(n_958),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_L g1148 ( 
.A1(n_951),
.A2(n_992),
.B(n_685),
.C(n_880),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1000),
.A2(n_1004),
.B(n_716),
.Y(n_1150)
);

OA22x2_ASAP7_75t_L g1151 ( 
.A1(n_872),
.A2(n_577),
.B1(n_542),
.B2(n_719),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_862),
.B(n_870),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_854),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_983),
.A2(n_899),
.B(n_993),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_996),
.B(n_997),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_992),
.A2(n_875),
.B(n_958),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_872),
.B(n_728),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_996),
.B(n_997),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_875),
.A2(n_692),
.B(n_996),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_883),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1055),
.B(n_1130),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1024),
.A2(n_1110),
.B(n_1100),
.Y(n_1166)
);

AO21x2_ASAP7_75t_L g1167 ( 
.A1(n_1036),
.A2(n_1049),
.B(n_1024),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1109),
.B(n_1116),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1111),
.A2(n_1149),
.B(n_1114),
.Y(n_1169)
);

CKINVDCx6p67_ASAP7_75t_R g1170 ( 
.A(n_1127),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1019),
.A2(n_1050),
.B1(n_1160),
.B2(n_1157),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1116),
.B(n_1135),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1153),
.A2(n_1161),
.B(n_1154),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1038),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1064),
.B(n_1151),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1087),
.B(n_1027),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1017),
.A2(n_1048),
.B(n_1033),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1069),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1143),
.B(n_1135),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1068),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1066),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1074),
.Y(n_1182)
);

OAI31xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1025),
.A2(n_1060),
.A3(n_1047),
.B(n_1052),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1123),
.A2(n_1151),
.B1(n_1029),
.B2(n_1108),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1054),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1021),
.A2(n_1158),
.B(n_1146),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_SL g1187 ( 
.A(n_1162),
.B(n_1080),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1136),
.B(n_1140),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1125),
.B(n_1132),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1122),
.A2(n_1159),
.B1(n_1029),
.B2(n_1052),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1072),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1028),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1155),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1062),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1044),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1112),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1072),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1136),
.B(n_1140),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1087),
.B(n_1051),
.Y(n_1199)
);

OR2x2_ASAP7_75t_SL g1200 ( 
.A(n_1096),
.B(n_1142),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1112),
.B(n_1057),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1093),
.A2(n_1031),
.B(n_1120),
.C(n_1150),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1030),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1148),
.A2(n_1016),
.B(n_1107),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1072),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1142),
.B(n_1145),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1145),
.B(n_1160),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1073),
.B(n_1112),
.Y(n_1208)
);

OR2x6_ASAP7_75t_SL g1209 ( 
.A(n_1157),
.B(n_1071),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1073),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1057),
.B(n_1043),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1076),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1070),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1096),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1058),
.B(n_1065),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1134),
.A2(n_1146),
.B(n_1147),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1113),
.B(n_1128),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1065),
.B(n_1144),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1048),
.A2(n_1022),
.B(n_1020),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1096),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1043),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1115),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1139),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1139),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1139),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1081),
.A2(n_1099),
.B(n_1022),
.C(n_1082),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1147),
.A2(n_1158),
.B(n_1126),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1036),
.A2(n_1095),
.B(n_1040),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1084),
.B(n_1071),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1129),
.B(n_1117),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1091),
.B(n_1087),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1092),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1042),
.A2(n_1035),
.B(n_1077),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1053),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1056),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_L g1236 ( 
.A(n_1056),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_1092),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1067),
.C(n_1078),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1091),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_SL g1240 ( 
.A1(n_1097),
.A2(n_1042),
.B(n_1078),
.C(n_1104),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1087),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1061),
.A2(n_1094),
.B1(n_1104),
.B2(n_1086),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1088),
.A2(n_1037),
.B(n_1098),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1085),
.B(n_1086),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1118),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1023),
.A2(n_1137),
.B(n_1141),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1085),
.B(n_1094),
.Y(n_1247)
);

NOR2x1_ASAP7_75t_SL g1248 ( 
.A(n_1118),
.B(n_1079),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1103),
.A2(n_1105),
.B(n_1138),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1090),
.B(n_1083),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1152),
.Y(n_1251)
);

AOI21xp33_ASAP7_75t_L g1252 ( 
.A1(n_1041),
.A2(n_1063),
.B(n_1034),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1152),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1039),
.B(n_1046),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1045),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1039),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1075),
.A2(n_1156),
.B1(n_1106),
.B2(n_1133),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1131),
.A2(n_1119),
.B1(n_1121),
.B2(n_1124),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1032),
.B(n_1026),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1060),
.B(n_602),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1019),
.A2(n_987),
.B1(n_1002),
.B2(n_997),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1018),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1060),
.B(n_602),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1073),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1019),
.A2(n_1050),
.B(n_1002),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1019),
.A2(n_1050),
.B(n_1060),
.C(n_1016),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1055),
.B(n_1130),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1072),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1019),
.A2(n_951),
.B(n_992),
.C(n_1022),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1069),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1273)
);

INVx5_ASAP7_75t_L g1274 ( 
.A(n_1072),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1060),
.B(n_602),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1019),
.A2(n_1050),
.B(n_1002),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1055),
.B(n_1130),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1069),
.Y(n_1278)
);

INVx3_ASAP7_75t_SL g1279 ( 
.A(n_1127),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1069),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1072),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1143),
.A2(n_599),
.B1(n_728),
.B2(n_1025),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1069),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1024),
.A2(n_992),
.B(n_1100),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1069),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1027),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1044),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1069),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1102),
.B(n_1125),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1019),
.A2(n_1050),
.B(n_1060),
.C(n_1016),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1044),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1055),
.B(n_1130),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1060),
.B(n_602),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_L g1294 ( 
.A(n_1050),
.B(n_1060),
.C(n_1019),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1112),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1024),
.A2(n_992),
.B(n_1100),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1073),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1027),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1044),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1026),
.B(n_1101),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1055),
.B(n_1130),
.Y(n_1303)
);

O2A1O1Ixp5_ASAP7_75t_L g1304 ( 
.A1(n_1019),
.A2(n_951),
.B(n_992),
.C(n_1022),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1245),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1211),
.B(n_1221),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1207),
.B(n_1206),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1194),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1274),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1286),
.B(n_1300),
.Y(n_1310)
);

CKINVDCx14_ASAP7_75t_R g1311 ( 
.A(n_1185),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1282),
.A2(n_1184),
.B1(n_1179),
.B2(n_1294),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1260),
.A2(n_1275),
.B1(n_1263),
.B2(n_1293),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1255),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1237),
.Y(n_1315)
);

BUFx4f_ASAP7_75t_SL g1316 ( 
.A(n_1264),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1250),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1243),
.A2(n_1228),
.B(n_1284),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1262),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1243),
.A2(n_1177),
.B(n_1166),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1178),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1231),
.B(n_1239),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1212),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1265),
.A2(n_1276),
.B1(n_1190),
.B2(n_1203),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1211),
.B(n_1265),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1256),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1261),
.A2(n_1276),
.B(n_1266),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1211),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1274),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1164),
.B(n_1168),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1183),
.B(n_1215),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1247),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1214),
.A2(n_1261),
.B1(n_1209),
.B2(n_1171),
.Y(n_1333)
);

BUFx4f_ASAP7_75t_SL g1334 ( 
.A(n_1299),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_1208),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1183),
.B(n_1229),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1171),
.A2(n_1290),
.B1(n_1217),
.B2(n_1188),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1254),
.Y(n_1338)
);

BUFx2_ASAP7_75t_R g1339 ( 
.A(n_1196),
.Y(n_1339)
);

AO21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1204),
.A2(n_1217),
.B(n_1163),
.Y(n_1340)
);

CKINVDCx11_ASAP7_75t_R g1341 ( 
.A(n_1279),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1175),
.A2(n_1291),
.B1(n_1287),
.B2(n_1195),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1201),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1272),
.Y(n_1344)
);

NOR2x1_ASAP7_75t_L g1345 ( 
.A(n_1201),
.B(n_1163),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1166),
.A2(n_1173),
.B(n_1169),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1180),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1234),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1278),
.Y(n_1349)
);

INVx4_ASAP7_75t_SL g1350 ( 
.A(n_1175),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1167),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1170),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1167),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1301),
.A2(n_1289),
.B1(n_1189),
.B2(n_1222),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1268),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1164),
.A2(n_1198),
.B1(n_1168),
.B2(n_1188),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1172),
.A2(n_1198),
.B1(n_1285),
.B2(n_1283),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1280),
.B(n_1288),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1268),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1182),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1271),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1193),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1270),
.A2(n_1304),
.B(n_1226),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1236),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1210),
.A2(n_1192),
.B1(n_1172),
.B2(n_1174),
.Y(n_1365)
);

INVx5_ASAP7_75t_L g1366 ( 
.A(n_1241),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1273),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1273),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1296),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1297),
.B(n_1302),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1297),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1181),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1230),
.A2(n_1220),
.B1(n_1218),
.B2(n_1204),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1259),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1259),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1244),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1233),
.B(n_1238),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1242),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1257),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1246),
.A2(n_1249),
.B(n_1169),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1173),
.A2(n_1252),
.B(n_1257),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1165),
.A2(n_1303),
.B1(n_1292),
.B2(n_1277),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1248),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1200),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1235),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1191),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1258),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1191),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1187),
.A2(n_1303),
.B1(n_1165),
.B2(n_1267),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1298),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1219),
.B(n_1269),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1213),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1191),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1186),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1224),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1216),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1267),
.A2(n_1277),
.B1(n_1292),
.B2(n_1232),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1295),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1227),
.A2(n_1253),
.B1(n_1176),
.B2(n_1199),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1202),
.A2(n_1240),
.B(n_1252),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1251),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1197),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1197),
.A2(n_1205),
.B(n_1223),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1176),
.A2(n_1199),
.B1(n_1225),
.B2(n_1205),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1281),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1281),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1281),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1197),
.A2(n_1205),
.B1(n_1223),
.B2(n_1269),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1223),
.A2(n_1243),
.B(n_1298),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1269),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1262),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1260),
.A2(n_1263),
.B1(n_1293),
.B2(n_1275),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1194),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1194),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1264),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1206),
.B(n_1211),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1185),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1241),
.Y(n_1419)
);

NOR2x1_ASAP7_75t_R g1420 ( 
.A(n_1185),
.B(n_602),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1255),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1194),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1340),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1308),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1417),
.B(n_1379),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1401),
.A2(n_1353),
.B(n_1351),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1319),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1323),
.B(n_1414),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1323),
.B(n_1414),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1338),
.B(n_1331),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1412),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_SL g1432 ( 
.A(n_1418),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1320),
.A2(n_1318),
.B(n_1381),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1415),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1360),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1362),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1325),
.B(n_1328),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1422),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1410),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1422),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1338),
.B(n_1331),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1320),
.A2(n_1318),
.B(n_1381),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1306),
.B(n_1370),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1336),
.B(n_1355),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1321),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1355),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1327),
.A2(n_1313),
.B1(n_1413),
.B2(n_1333),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1344),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1359),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1337),
.A2(n_1363),
.B(n_1312),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1305),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1392),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1359),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1392),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1324),
.A2(n_1345),
.B(n_1378),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1361),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1361),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1305),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1367),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1336),
.B(n_1367),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1325),
.B(n_1350),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1368),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1307),
.B(n_1330),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1306),
.B(n_1377),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1349),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1368),
.B(n_1369),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1369),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1382),
.A2(n_1380),
.B(n_1391),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1371),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1371),
.B(n_1377),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1325),
.B(n_1350),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1386),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1419),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1317),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1314),
.Y(n_1475)
);

NAND2x1_ASAP7_75t_L g1476 ( 
.A(n_1384),
.B(n_1314),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1326),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1373),
.A2(n_1356),
.B1(n_1399),
.B2(n_1390),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1326),
.Y(n_1479)
);

BUFx4f_ASAP7_75t_SL g1480 ( 
.A(n_1418),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1378),
.B(n_1317),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1317),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1347),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1374),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1375),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1358),
.B(n_1376),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1375),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1358),
.B(n_1376),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1335),
.A2(n_1354),
.B1(n_1357),
.B2(n_1383),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1332),
.B(n_1314),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1348),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1350),
.B(n_1421),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1365),
.B(n_1310),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1348),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1421),
.B(n_1388),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1397),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1384),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1346),
.Y(n_1499)
);

AOI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1346),
.A2(n_1404),
.B(n_1409),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1406),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1424),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1430),
.B(n_1346),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1466),
.B(n_1322),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1435),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1441),
.B(n_1444),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1441),
.B(n_1407),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1436),
.Y(n_1508)
);

OAI33xp33_ASAP7_75t_L g1509 ( 
.A1(n_1447),
.A2(n_1385),
.A3(n_1402),
.B1(n_1411),
.B2(n_1406),
.B3(n_1407),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1444),
.B(n_1408),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1460),
.B(n_1408),
.Y(n_1511)
);

OAI33xp33_ASAP7_75t_L g1512 ( 
.A1(n_1478),
.A2(n_1402),
.A3(n_1411),
.B1(n_1405),
.B2(n_1393),
.B3(n_1352),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1454),
.B(n_1452),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1423),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1460),
.B(n_1403),
.Y(n_1515)
);

INVxp67_ASAP7_75t_SL g1516 ( 
.A(n_1499),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1428),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1322),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1423),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1450),
.A2(n_1398),
.B1(n_1400),
.B2(n_1315),
.C(n_1342),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1454),
.B(n_1343),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1445),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1470),
.B(n_1343),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1481),
.B(n_1403),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1443),
.B(n_1428),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1429),
.B(n_1396),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1394),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1432),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1474),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1448),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1465),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1470),
.B(n_1343),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1454),
.B(n_1366),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1429),
.B(n_1464),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1427),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1425),
.B(n_1389),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1425),
.B(n_1389),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1476),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1492),
.B(n_1366),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1490),
.B(n_1495),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1490),
.B(n_1495),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1464),
.B(n_1396),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1482),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1486),
.B(n_1387),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1505),
.B(n_1431),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1535),
.B(n_1451),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1508),
.B(n_1472),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_SL g1548 ( 
.A(n_1528),
.B(n_1352),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1516),
.A2(n_1442),
.B(n_1433),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1522),
.B(n_1486),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1506),
.B(n_1497),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1530),
.B(n_1488),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1531),
.B(n_1455),
.C(n_1501),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1506),
.B(n_1488),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1520),
.A2(n_1489),
.B1(n_1458),
.B2(n_1493),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1540),
.B(n_1497),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1539),
.B(n_1483),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1517),
.B(n_1525),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1520),
.A2(n_1489),
.B1(n_1399),
.B2(n_1491),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1529),
.B(n_1477),
.C(n_1479),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1517),
.B(n_1463),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1426),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1529),
.B(n_1477),
.C(n_1479),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1541),
.B(n_1426),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1446),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1541),
.B(n_1426),
.Y(n_1566)
);

AND2x2_ASAP7_75t_SL g1567 ( 
.A(n_1521),
.B(n_1461),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1516),
.A2(n_1442),
.B(n_1433),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1534),
.B(n_1510),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1534),
.B(n_1446),
.Y(n_1570)
);

AND2x2_ASAP7_75t_SL g1571 ( 
.A(n_1521),
.B(n_1461),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1526),
.B(n_1480),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1510),
.B(n_1449),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1543),
.B(n_1372),
.C(n_1491),
.Y(n_1574)
);

NAND4xp25_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1494),
.C(n_1485),
.D(n_1487),
.Y(n_1575)
);

OAI221xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1542),
.A2(n_1503),
.B1(n_1532),
.B2(n_1523),
.C(n_1504),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1511),
.B(n_1475),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1504),
.B(n_1372),
.C(n_1494),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1512),
.A2(n_1471),
.B1(n_1461),
.B2(n_1437),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_1341),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1507),
.B(n_1434),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_1453),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1453),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1507),
.B(n_1438),
.Y(n_1584)
);

OAI221xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1542),
.A2(n_1456),
.B1(n_1457),
.B2(n_1459),
.C(n_1462),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1515),
.B(n_1456),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1518),
.A2(n_1440),
.B(n_1469),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1512),
.B(n_1315),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_SL g1589 ( 
.A(n_1519),
.B(n_1393),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1509),
.B(n_1500),
.C(n_1439),
.Y(n_1590)
);

NAND4xp25_ASAP7_75t_L g1591 ( 
.A(n_1514),
.B(n_1485),
.C(n_1487),
.D(n_1496),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1518),
.A2(n_1500),
.B(n_1498),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1502),
.B(n_1372),
.C(n_1467),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1524),
.B(n_1459),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1549),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1562),
.B(n_1564),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1588),
.B(n_1509),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1556),
.B(n_1527),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1560),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1527),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1551),
.B(n_1524),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1590),
.B(n_1467),
.C(n_1462),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1563),
.Y(n_1605)
);

AND2x2_ASAP7_75t_SL g1606 ( 
.A(n_1567),
.B(n_1471),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1502),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1549),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1549),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1549),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1558),
.B(n_1468),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1563),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1568),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1553),
.B(n_1538),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1570),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1565),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1581),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1581),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1568),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1562),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1568),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1584),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1567),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1553),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1564),
.B(n_1536),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1575),
.B(n_1468),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1566),
.B(n_1536),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1568),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1566),
.B(n_1537),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1533),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1575),
.B(n_1468),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1607),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1618),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1617),
.B(n_1569),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1550),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1624),
.B(n_1592),
.C(n_1559),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1600),
.B(n_1552),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1587),
.Y(n_1638)
);

INVxp33_ASAP7_75t_L g1639 ( 
.A(n_1598),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1607),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1617),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1618),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1618),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1622),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1598),
.B(n_1545),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1596),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1623),
.B(n_1630),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1622),
.Y(n_1648)
);

NOR2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1606),
.B(n_1339),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1596),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1554),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1623),
.B(n_1577),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1561),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1577),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1625),
.B(n_1546),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1547),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1603),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1603),
.B(n_1573),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1603),
.B(n_1582),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1605),
.B(n_1612),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1605),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1605),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1612),
.B(n_1583),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1612),
.B(n_1594),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1586),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1596),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1625),
.B(n_1567),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1659),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1663),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1635),
.B(n_1604),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1602),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1645),
.B(n_1616),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1669),
.B(n_1602),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1664),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1647),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1655),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1647),
.B(n_1602),
.Y(n_1681)
);

AOI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1639),
.A2(n_1620),
.A3(n_1626),
.B1(n_1631),
.B2(n_1555),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1658),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1667),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1667),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_SL g1687 ( 
.A(n_1639),
.B(n_1604),
.C(n_1626),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1646),
.Y(n_1688)
);

NAND2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1671),
.B(n_1606),
.Y(n_1689)
);

NAND2x1p5_ASAP7_75t_L g1690 ( 
.A(n_1649),
.B(n_1606),
.Y(n_1690)
);

NOR2x1_ASAP7_75t_R g1691 ( 
.A(n_1638),
.B(n_1416),
.Y(n_1691)
);

NAND2x1p5_ASAP7_75t_L g1692 ( 
.A(n_1651),
.B(n_1606),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1662),
.Y(n_1693)
);

AOI322xp5_ASAP7_75t_L g1694 ( 
.A1(n_1670),
.A2(n_1597),
.A3(n_1620),
.B1(n_1610),
.B2(n_1619),
.C1(n_1596),
.C2(n_1608),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1632),
.Y(n_1696)
);

XOR2x2_ASAP7_75t_L g1697 ( 
.A(n_1636),
.B(n_1574),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1640),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1652),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1660),
.B(n_1616),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1661),
.A2(n_1626),
.B(n_1631),
.C(n_1620),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1657),
.B(n_1616),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1661),
.Y(n_1706)
);

OR2x6_ASAP7_75t_L g1707 ( 
.A(n_1654),
.B(n_1593),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1666),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1637),
.B(n_1597),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1656),
.B(n_1599),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1665),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1656),
.B(n_1599),
.Y(n_1712)
);

OAI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1665),
.A2(n_1666),
.B(n_1631),
.Y(n_1713)
);

AOI322xp5_ASAP7_75t_L g1714 ( 
.A1(n_1657),
.A2(n_1597),
.A3(n_1610),
.B1(n_1619),
.B2(n_1609),
.C1(n_1613),
.C2(n_1608),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1672),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1697),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1673),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1706),
.B(n_1641),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1697),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1682),
.A2(n_1687),
.B1(n_1713),
.B2(n_1704),
.C(n_1694),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1687),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1690),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1711),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1691),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1693),
.Y(n_1725)
);

CKINVDCx16_ASAP7_75t_R g1726 ( 
.A(n_1707),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1699),
.B(n_1316),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1683),
.B(n_1625),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1688),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1676),
.B(n_1633),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1690),
.B(n_1599),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1625),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1678),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1708),
.B(n_1642),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1685),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1674),
.A2(n_1626),
.B1(n_1631),
.B2(n_1668),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1686),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1688),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1714),
.B(n_1609),
.C(n_1608),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1707),
.A2(n_1668),
.B1(n_1652),
.B2(n_1579),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1696),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1700),
.B(n_1608),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_1599),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1689),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1709),
.B(n_1643),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1698),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1701),
.B(n_1627),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1695),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1705),
.B(n_1627),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1675),
.B(n_1601),
.Y(n_1750)
);

OAI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1721),
.A2(n_1692),
.B1(n_1707),
.B2(n_1679),
.Y(n_1751)
);

AOI222xp33_ASAP7_75t_L g1752 ( 
.A1(n_1719),
.A2(n_1716),
.B1(n_1720),
.B2(n_1736),
.C1(n_1739),
.C2(n_1721),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1716),
.A2(n_1679),
.B(n_1681),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1741),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1334),
.Y(n_1755)
);

AOI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1719),
.A2(n_1702),
.B(n_1695),
.Y(n_1756)
);

OAI322xp33_ASAP7_75t_L g1757 ( 
.A1(n_1726),
.A2(n_1613),
.A3(n_1628),
.B1(n_1610),
.B2(n_1621),
.C1(n_1609),
.C2(n_1619),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1742),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1726),
.B(n_1710),
.Y(n_1759)
);

OR3x2_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1420),
.C(n_1591),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1731),
.B(n_1675),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1742),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1723),
.B(n_1710),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1740),
.A2(n_1684),
.B1(n_1702),
.B2(n_1692),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1715),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1723),
.A2(n_1700),
.B1(n_1679),
.B2(n_1684),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1731),
.B(n_1677),
.Y(n_1768)
);

AOI32xp33_ASAP7_75t_L g1769 ( 
.A1(n_1722),
.A2(n_1684),
.A3(n_1609),
.B1(n_1613),
.B2(n_1628),
.Y(n_1769)
);

OAI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1739),
.A2(n_1621),
.B1(n_1610),
.B2(n_1628),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1725),
.A2(n_1613),
.B1(n_1628),
.B2(n_1619),
.C(n_1621),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1724),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1715),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1725),
.B(n_1712),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1750),
.B(n_1677),
.Y(n_1775)
);

OAI322xp33_ASAP7_75t_L g1776 ( 
.A1(n_1746),
.A2(n_1621),
.A3(n_1703),
.B1(n_1611),
.B2(n_1650),
.C1(n_1648),
.C2(n_1644),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1717),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1758),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1755),
.B(n_1727),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1755),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1773),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1772),
.B(n_1746),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1763),
.B(n_1733),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1774),
.B(n_1733),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1759),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1758),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1754),
.B(n_1730),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1762),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1773),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1752),
.B(n_1735),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1765),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1775),
.B(n_1735),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1777),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1761),
.B(n_1750),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1762),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1775),
.B(n_1730),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1761),
.B(n_1737),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1766),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1780),
.A2(n_1751),
.B(n_1767),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1782),
.B(n_1722),
.C(n_1768),
.D(n_1769),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1790),
.A2(n_1753),
.B(n_1756),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1778),
.A2(n_1770),
.B1(n_1764),
.B2(n_1757),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1794),
.B(n_1768),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1794),
.B(n_1681),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1796),
.B(n_1737),
.Y(n_1805)
);

AND4x1_ASAP7_75t_L g1806 ( 
.A(n_1779),
.B(n_1760),
.C(n_1743),
.D(n_1311),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1796),
.B(n_1700),
.Y(n_1807)
);

OAI21xp33_ASAP7_75t_L g1808 ( 
.A1(n_1785),
.A2(n_1722),
.B(n_1744),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1783),
.B(n_1744),
.Y(n_1809)
);

AOI21xp33_ASAP7_75t_L g1810 ( 
.A1(n_1795),
.A2(n_1766),
.B(n_1738),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1784),
.A2(n_1760),
.B1(n_1743),
.B2(n_1732),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1778),
.A2(n_1771),
.B1(n_1718),
.B2(n_1729),
.C(n_1748),
.Y(n_1812)
);

NAND4xp75_ASAP7_75t_L g1813 ( 
.A(n_1801),
.B(n_1798),
.C(n_1788),
.D(n_1786),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1807),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1803),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1805),
.Y(n_1816)
);

NAND3xp33_ASAP7_75t_L g1817 ( 
.A(n_1801),
.B(n_1799),
.C(n_1808),
.Y(n_1817)
);

AOI211xp5_ASAP7_75t_L g1818 ( 
.A1(n_1811),
.A2(n_1776),
.B(n_1787),
.C(n_1797),
.Y(n_1818)
);

AND5x1_ASAP7_75t_L g1819 ( 
.A(n_1800),
.B(n_1802),
.C(n_1806),
.D(n_1812),
.E(n_1810),
.Y(n_1819)
);

NOR3x1_ASAP7_75t_L g1820 ( 
.A(n_1809),
.B(n_1787),
.C(n_1792),
.Y(n_1820)
);

NAND4xp25_ASAP7_75t_L g1821 ( 
.A(n_1804),
.B(n_1793),
.C(n_1791),
.D(n_1789),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1801),
.Y(n_1822)
);

OAI322xp33_ASAP7_75t_L g1823 ( 
.A1(n_1801),
.A2(n_1789),
.A3(n_1781),
.B1(n_1788),
.B2(n_1786),
.C1(n_1717),
.C2(n_1718),
.Y(n_1823)
);

NOR3xp33_ASAP7_75t_L g1824 ( 
.A(n_1801),
.B(n_1781),
.C(n_1738),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_L g1825 ( 
.A1(n_1822),
.A2(n_1742),
.B(n_1548),
.C(n_1734),
.Y(n_1825)
);

NOR3xp33_ASAP7_75t_SL g1826 ( 
.A(n_1817),
.B(n_1813),
.C(n_1823),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_SL g1827 ( 
.A(n_1824),
.B(n_1738),
.C(n_1729),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_L g1828 ( 
.A(n_1815),
.B(n_1734),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1824),
.A2(n_1748),
.B(n_1729),
.C(n_1745),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_L g1830 ( 
.A(n_1821),
.B(n_1745),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1828),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1827),
.B(n_1820),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1829),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1830),
.Y(n_1834)
);

NOR3x2_ASAP7_75t_L g1835 ( 
.A(n_1826),
.B(n_1819),
.C(n_1816),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1825),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1827),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1834),
.B(n_1814),
.Y(n_1838)
);

NAND4xp75_ASAP7_75t_L g1839 ( 
.A(n_1832),
.B(n_1818),
.C(n_1748),
.D(n_1728),
.Y(n_1839)
);

NAND4xp25_ASAP7_75t_L g1840 ( 
.A(n_1834),
.B(n_1836),
.C(n_1831),
.D(n_1833),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1835),
.B(n_1747),
.C(n_1749),
.Y(n_1841)
);

NAND4xp75_ASAP7_75t_L g1842 ( 
.A(n_1837),
.B(n_1712),
.C(n_1606),
.D(n_1572),
.Y(n_1842)
);

NAND4xp75_ASAP7_75t_L g1843 ( 
.A(n_1837),
.B(n_1557),
.C(n_1571),
.D(n_1627),
.Y(n_1843)
);

XNOR2xp5_ASAP7_75t_L g1844 ( 
.A(n_1839),
.B(n_1578),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1838),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1842),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1845),
.Y(n_1847)
);

NAND5xp2_ASAP7_75t_L g1848 ( 
.A(n_1847),
.B(n_1840),
.C(n_1846),
.D(n_1841),
.E(n_1844),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1848),
.B(n_1843),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1848),
.A2(n_1593),
.B(n_1578),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1849),
.A2(n_1611),
.B1(n_1634),
.B2(n_1576),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1850),
.A2(n_1589),
.B(n_1627),
.Y(n_1852)
);

AOI21xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1851),
.A2(n_1329),
.B(n_1309),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1852),
.A2(n_1629),
.B(n_1601),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1853),
.A2(n_1591),
.B(n_1629),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1855),
.A2(n_1854),
.B1(n_1629),
.B2(n_1364),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1629),
.B1(n_1585),
.B2(n_1630),
.C(n_1611),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1473),
.B(n_1364),
.C(n_1419),
.Y(n_1858)
);


endmodule