module real_jpeg_25263_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_0),
.A2(n_51),
.B1(n_52),
.B2(n_66),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_0),
.A2(n_36),
.B1(n_40),
.B2(n_66),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_0),
.A2(n_22),
.B1(n_24),
.B2(n_66),
.Y(n_207)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_5),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_25),
.B1(n_36),
.B2(n_40),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_31),
.B1(n_36),
.B2(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_31),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_36),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_8),
.A2(n_22),
.B1(n_24),
.B2(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_43),
.B1(n_65),
.B2(n_72),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_8),
.A2(n_62),
.B(n_73),
.C(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_60),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_8),
.A2(n_49),
.B(n_51),
.C(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_8),
.B(n_24),
.C(n_39),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_8),
.B(n_150),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_8),
.B(n_213),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_8),
.B(n_41),
.Y(n_223)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_133),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_132),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_111),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_16),
.B(n_111),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_77),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.C(n_58),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_18),
.A2(n_19),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_20),
.B(n_32),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_28),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_21),
.A2(n_83),
.B(n_87),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_22),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_24),
.B(n_219),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_26),
.B(n_30),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_26),
.A2(n_84),
.B(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_26),
.B(n_86),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_26),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_27),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_29),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_29),
.B(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_44),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_33),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_42),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_34),
.B(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_34),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_40),
.B1(n_49),
.B2(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_36),
.B(n_195),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_40),
.A2(n_43),
.B(n_54),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_41),
.B(n_182),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_42),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_43),
.A2(n_51),
.B(n_61),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_44),
.A2(n_90),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_44),
.B(n_181),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_46),
.A2(n_58),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_46),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_55),
.B(n_56),
.Y(n_46)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_47),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_47),
.B(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_55),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_48)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_55),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_56),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_57),
.B(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_58),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_69),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_59),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_60),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_74),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_70),
.Y(n_97)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_96),
.Y(n_142)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_105),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_92),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_81),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_87),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_89),
.A2(n_109),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_89),
.B(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_91),
.B(n_192),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_123),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_103),
.B(n_149),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_106),
.A2(n_110),
.B1(n_176),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.C(n_131),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_112),
.A2(n_113),
.B1(n_131),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_118),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_131),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_169),
.B(n_244),
.C(n_249),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_157),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_135),
.B(n_157),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_153),
.B2(n_156),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_151),
.B2(n_152),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_138),
.B(n_152),
.C(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_146),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_141),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_163),
.C(n_164),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_159),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_164),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_243),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_186),
.B(n_242),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_183),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_172),
.B(n_183),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_178),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_175),
.B(n_178),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_176),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_237),
.B(n_241),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_228),
.B(n_236),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_209),
.B(n_227),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_196),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_193),
.B1(n_194),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_203),
.B2(n_208),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_202),
.C(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_216),
.B(n_226),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_222),
.B(n_225),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_239),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);


endmodule