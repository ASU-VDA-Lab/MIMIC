module real_jpeg_33947_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_682, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_682;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_666;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_620;
wire n_332;
wire n_456;
wire n_366;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_675;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_313;
wire n_268;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_0),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_0),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_1),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_3),
.A2(n_342),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_3),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_3),
.A2(n_370),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_3),
.A2(n_370),
.B1(n_495),
.B2(n_498),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_3),
.A2(n_370),
.B1(n_594),
.B2(n_597),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_4),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_4),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_138),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_4),
.A2(n_138),
.B1(n_224),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_4),
.A2(n_138),
.B1(n_410),
.B2(n_413),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_5),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_5),
.A2(n_82),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_5),
.A2(n_82),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_5),
.A2(n_82),
.B1(n_576),
.B2(n_578),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_6),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_6),
.A2(n_130),
.B1(n_348),
.B2(n_352),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_6),
.A2(n_423),
.B(n_426),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_6),
.B(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_6),
.A2(n_130),
.B1(n_604),
.B2(n_607),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_7),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_7),
.A2(n_226),
.B1(n_374),
.B2(n_377),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_7),
.A2(n_226),
.B1(n_443),
.B2(n_448),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_7),
.A2(n_226),
.B1(n_257),
.B2(n_552),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_43),
.B1(n_46),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_8),
.A2(n_49),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_8),
.A2(n_49),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_8),
.A2(n_49),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_11),
.Y(n_364)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_12),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_13),
.A2(n_107),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_13),
.A2(n_107),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_13),
.A2(n_107),
.B1(n_547),
.B2(n_548),
.Y(n_546)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_14),
.A2(n_153),
.A3(n_333),
.B1(n_337),
.B2(n_340),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_14),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_14),
.A2(n_214),
.B1(n_341),
.B2(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_14),
.B(n_176),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_14),
.A2(n_32),
.B1(n_510),
.B2(n_516),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_14),
.A2(n_117),
.B(n_539),
.C(n_542),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_14),
.B(n_543),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_15),
.Y(n_672)
);

CKINVDCx11_ASAP7_75t_R g680 ( 
.A(n_15),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_16),
.A2(n_387),
.B1(n_389),
.B2(n_391),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_16),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_16),
.A2(n_205),
.B1(n_391),
.B2(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_16),
.A2(n_391),
.B1(n_496),
.B2(n_511),
.Y(n_510)
);

AO22x1_ASAP7_75t_L g536 ( 
.A1(n_16),
.A2(n_112),
.B1(n_391),
.B2(n_537),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_18),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_18),
.A2(n_89),
.B1(n_193),
.B2(n_196),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_18),
.A2(n_89),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_18),
.A2(n_89),
.B1(n_131),
.B2(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_19),
.Y(n_141)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_19),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_19),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_663),
.B(n_674),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_21),
.A2(n_675),
.B(n_677),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_321),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_311),
.B(n_320),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_294),
.B(n_310),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_266),
.B(n_293),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_232),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_26),
.B(n_232),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_135),
.C(n_189),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_28),
.B(n_135),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_93),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_29),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_50),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_30),
.A2(n_264),
.B1(n_265),
.B2(n_682),
.Y(n_263)
);

XOR2x2_ASAP7_75t_SL g642 ( 
.A(n_30),
.B(n_50),
.Y(n_642)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_38),
.B(n_41),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_31),
.A2(n_347),
.B1(n_355),
.B2(n_359),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_31),
.A2(n_359),
.B1(n_406),
.B2(n_409),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_31),
.A2(n_493),
.B1(n_502),
.B2(n_503),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_31),
.B(n_409),
.Y(n_580)
);

AO22x1_ASAP7_75t_L g614 ( 
.A1(n_31),
.A2(n_355),
.B1(n_615),
.B2(n_616),
.Y(n_614)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_32),
.A2(n_42),
.B1(n_192),
.B2(n_198),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_32),
.A2(n_442),
.B1(n_450),
.B2(n_454),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_32),
.A2(n_198),
.B1(n_494),
.B2(n_510),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_35),
.Y(n_453)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_35),
.Y(n_505)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_36),
.Y(n_197)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_36),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_37),
.Y(n_351)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_37),
.Y(n_512)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_45),
.Y(n_412)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_75),
.B1(n_83),
.B2(n_84),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_51),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_51),
.A2(n_75),
.B1(n_83),
.B2(n_203),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_51),
.A2(n_83),
.B(n_181),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_51),
.A2(n_83),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_51),
.A2(n_83),
.B1(n_369),
.B2(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_51),
.A2(n_83),
.B1(n_422),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_51),
.Y(n_619)
);

AO21x2_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_60),
.B(n_67),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_59),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_60),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_62),
.Y(n_186)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_62),
.Y(n_345)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_62),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_63),
.Y(n_208)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_78),
.Y(n_204)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_79),
.Y(n_549)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_80),
.Y(n_378)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_81),
.Y(n_438)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_83),
.B(n_341),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_84),
.Y(n_178)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_94),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_106),
.B(n_116),
.Y(n_94)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_95),
.Y(n_237)
);

AOI22x1_ASAP7_75t_L g591 ( 
.A1(n_95),
.A2(n_246),
.B1(n_536),
.B2(n_592),
.Y(n_591)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_96),
.A2(n_221),
.B1(n_222),
.B2(n_231),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_96),
.A2(n_238),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_96),
.A2(n_275),
.B1(n_277),
.B2(n_304),
.Y(n_303)
);

OAI22x1_ASAP7_75t_R g312 ( 
.A1(n_96),
.A2(n_221),
.B1(n_304),
.B2(n_313),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g403 ( 
.A(n_96),
.B(n_341),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_96),
.A2(n_221),
.B1(n_222),
.B2(n_593),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_96),
.A2(n_275),
.B(n_313),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_100),
.Y(n_397)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_102),
.Y(n_572)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_103),
.Y(n_217)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_106),
.Y(n_247)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_110),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_115),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_115),
.Y(n_244)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_115),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_115),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_115),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_128),
.Y(n_116)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_117),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_121),
.Y(n_596)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_123),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_133),
.Y(n_541)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_134),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_134),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_177),
.B(n_188),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_177),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_145),
.B1(n_169),
.B2(n_176),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_137),
.B(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_140),
.Y(n_288)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_145),
.A2(n_211),
.B(n_218),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_145),
.A2(n_176),
.B(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_146),
.A2(n_251),
.B1(n_252),
.B2(n_260),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_146),
.A2(n_252),
.B1(n_260),
.B2(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_146),
.A2(n_260),
.B1(n_381),
.B2(n_386),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_146),
.A2(n_260),
.B1(n_386),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_146),
.A2(n_260),
.B1(n_395),
.B2(n_551),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_146),
.A2(n_260),
.B1(n_551),
.B2(n_603),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_146),
.A2(n_212),
.B1(n_260),
.B2(n_603),
.Y(n_630)
);

AO21x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_153),
.B(n_161),
.Y(n_146)
);

NAND2xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_156),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_156),
.Y(n_606)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_162),
.B1(n_165),
.B2(n_167),
.Y(n_161)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_162),
.Y(n_425)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_164),
.Y(n_472)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_165),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_166),
.Y(n_372)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_169),
.Y(n_251)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_187),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_179),
.A2(n_187),
.B1(n_368),
.B2(n_373),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_179),
.A2(n_187),
.B1(n_435),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g617 ( 
.A1(n_187),
.A2(n_618),
.B1(n_619),
.B2(n_620),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_189),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_209),
.C(n_219),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_190),
.B(n_644),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_202),
.Y(n_190)
);

XOR2x2_ASAP7_75t_SL g636 ( 
.A(n_191),
.B(n_202),
.Y(n_636)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_192),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_194),
.Y(n_414)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_195),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_195),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_203),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_207),
.Y(n_427)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_208),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_210),
.B(n_220),
.Y(n_644)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx4f_ASAP7_75t_L g390 ( 
.A(n_217),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_263),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_263),
.C(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_248),
.Y(n_235)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_245),
.B2(n_247),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_237),
.A2(n_535),
.B(n_538),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_261),
.B2(n_262),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_249),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_249),
.A2(n_262),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_274),
.C(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_262),
.C(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_257),
.B(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_269),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_271),
.C(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_273),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_282),
.Y(n_601)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_292),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_292),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_308),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_308),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_301),
.C(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_319),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_312),
.B(n_666),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_312),
.Y(n_669)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.C(n_327),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_584),
.B(n_658),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_429),
.B(n_527),
.C(n_582),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_392),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_330),
.B(n_392),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_367),
.C(n_379),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_331),
.B(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_346),
.B1(n_365),
.B2(n_366),
.Y(n_331)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_332),
.B(n_366),
.Y(n_418)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_SL g464 ( 
.A1(n_341),
.A2(n_465),
.B(n_469),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_341),
.B(n_470),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_341),
.B(n_451),
.Y(n_519)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_351),
.Y(n_577)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_353),
.Y(n_578)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_355),
.Y(n_579)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_364),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_364),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_367),
.A2(n_379),
.B1(n_380),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_385),
.Y(n_388)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_415),
.B1(n_416),
.B2(n_428),
.Y(n_392)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_393),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_394),
.B(n_403),
.C(n_404),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_397),
.Y(n_554)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_400),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_417),
.B(n_420),
.C(n_428),
.Y(n_531)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_458),
.B(n_526),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_455),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_432),
.B(n_455),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_439),
.C(n_441),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_433),
.A2(n_439),
.B1(n_440),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_433),
.Y(n_489)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_488),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_443),
.A2(n_475),
.B1(n_485),
.B2(n_486),
.Y(n_474)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_490),
.B(n_525),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_487),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_461),
.B(n_487),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_473),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_462),
.A2(n_463),
.B1(n_473),
.B2(n_474),
.Y(n_506)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_480),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_507),
.B(n_524),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_506),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_492),
.B(n_506),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx2_ASAP7_75t_SL g522 ( 
.A(n_497),
.Y(n_522)
);

BUFx2_ASAP7_75t_SL g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_508),
.A2(n_514),
.B(n_523),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_513),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_509),
.B(n_513),
.Y(n_523)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_518),
.Y(n_514)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_532),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_531),
.B(n_583),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_532),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_555),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_533),
.B(n_556),
.C(n_581),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_544),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_534),
.B(n_545),
.C(n_550),
.Y(n_611)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_537),
.Y(n_543)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx3_ASAP7_75t_SL g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_542),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_550),
.Y(n_544)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_581),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_574),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_557),
.B(n_574),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_562),
.B1(n_568),
.B2(n_573),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_566),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx3_ASAP7_75t_SL g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_575),
.A2(n_579),
.B(n_580),
.Y(n_574)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_575),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

NAND4xp25_ASAP7_75t_SL g584 ( 
.A(n_585),
.B(n_622),
.C(n_645),
.D(n_651),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_587),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_586),
.B(n_587),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_610),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_588),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_590),
.Y(n_588)
);

MAJx2_ASAP7_75t_L g633 ( 
.A(n_589),
.B(n_634),
.C(n_635),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_602),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx4_ASAP7_75t_SL g595 ( 
.A(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_602),
.Y(n_634)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_611),
.A2(n_612),
.B1(n_613),
.B2(n_621),
.Y(n_610)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_611),
.Y(n_621)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

HB1xp67_ASAP7_75t_SL g654 ( 
.A(n_613),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_614),
.B(n_617),
.Y(n_613)
);

NAND2x1_ASAP7_75t_SL g626 ( 
.A(n_614),
.B(n_617),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_621),
.Y(n_655)
);

A2O1A1O1Ixp25_ASAP7_75t_L g658 ( 
.A1(n_622),
.A2(n_645),
.B(n_659),
.C(n_661),
.D(n_662),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_637),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_623),
.B(n_637),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_632),
.C(n_636),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_625),
.B(n_636),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_626),
.B(n_627),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_626),
.B(n_639),
.C(n_640),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_628),
.A2(n_629),
.B1(n_630),
.B2(n_631),
.Y(n_627)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_628),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_629),
.Y(n_640)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_631),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_633),
.Y(n_632)
);

XNOR2x1_ASAP7_75t_L g656 ( 
.A(n_633),
.B(n_657),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_638),
.B(n_641),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_638),
.B(n_642),
.C(n_647),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_642),
.B(n_643),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_643),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_646),
.B(n_648),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_646),
.B(n_648),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_650),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_652),
.B(n_656),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_652),
.B(n_656),
.C(n_660),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_653),
.B(n_654),
.C(n_655),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_664),
.B(n_670),
.Y(n_663)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_664),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_665),
.B(n_668),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g666 ( 
.A(n_667),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_667),
.B(n_669),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_670),
.B(n_676),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_670),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_671),
.B(n_673),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_672),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_678),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_679),
.B(n_680),
.Y(n_678)
);


endmodule