module fake_netlist_6_1035_n_580 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_580);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_580;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_16),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_40),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_48),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_18),
.Y(n_137)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_37),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_58),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_61),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_71),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_49),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_26),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_114),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_19),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_31),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_60),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_21),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_25),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_99),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_20),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_74),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_72),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_24),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_87),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_42),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_52),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_30),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_35),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_23),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_34),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_46),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_45),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_0),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

INVxp33_ASAP7_75t_SL g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_137),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_0),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_139),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_134),
.B(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_149),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_2),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_147),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_151),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_154),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_156),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_157),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_158),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_3),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_159),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_138),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_195),
.B(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_196),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_146),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_190),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_133),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_218),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_172),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_198),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_180),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_246),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_186),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_250),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_161),
.Y(n_290)
);

NAND3x1_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_188),
.C(n_184),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_185),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_162),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_183),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_178),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_181),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_167),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_275),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_168),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_257),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_169),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_173),
.Y(n_307)
);

BUFx4f_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_148),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_182),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

AND2x6_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_148),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_265),
.Y(n_314)
);

AND3x4_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_4),
.C(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_273),
.B(n_174),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_273),
.B(n_267),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_179),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_176),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_239),
.B(n_13),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_269),
.A2(n_148),
.B1(n_5),
.B2(n_6),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_240),
.B(n_148),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_250),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_4),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_270),
.B(n_14),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_240),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_264),
.B(n_7),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_240),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_266),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_243),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_249),
.B(n_8),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_252),
.B(n_8),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_289),
.A2(n_288),
.B1(n_244),
.B2(n_337),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_237),
.B1(n_241),
.B2(n_248),
.Y(n_342)
);

OA22x2_ASAP7_75t_L g343 ( 
.A1(n_300),
.A2(n_252),
.B1(n_284),
.B2(n_261),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_251),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_259),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_286),
.B(n_314),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_296),
.B(n_262),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_248),
.B1(n_10),
.B2(n_11),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

NOR2x1p5_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_243),
.Y(n_353)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_285),
.A2(n_247),
.B1(n_242),
.B2(n_254),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_247),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_328),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_299),
.A2(n_260),
.B1(n_254),
.B2(n_253),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_306),
.Y(n_361)
);

AO22x2_ASAP7_75t_L g362 ( 
.A1(n_317),
.A2(n_9),
.B1(n_10),
.B2(n_260),
.Y(n_362)
);

OAI221xp5_ASAP7_75t_L g363 ( 
.A1(n_322),
.A2(n_253),
.B1(n_245),
.B2(n_284),
.C(n_9),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_319),
.B(n_331),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

AO22x2_ASAP7_75t_L g370 ( 
.A1(n_298),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_307),
.B(n_38),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g374 ( 
.A1(n_332),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_51),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g378 ( 
.A1(n_299),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_295),
.B(n_126),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_310),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_308),
.B(n_64),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_293),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_308),
.B(n_65),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_316),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_346),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_341),
.B(n_320),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_344),
.B(n_297),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_344),
.B(n_323),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_294),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_330),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_345),
.B(n_323),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_371),
.B(n_324),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_367),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_340),
.B(n_324),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_359),
.B(n_287),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_353),
.B(n_291),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_382),
.B(n_287),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_383),
.B(n_287),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_309),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_368),
.B(n_325),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_380),
.B(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_357),
.B(n_313),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_385),
.B(n_66),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_SL g408 ( 
.A(n_387),
.B(n_67),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_68),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_351),
.B(n_69),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_352),
.B(n_70),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_73),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_355),
.B(n_76),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_343),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_360),
.B(n_365),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_78),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_381),
.B(n_81),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_342),
.B(n_82),
.Y(n_418)
);

AO31x2_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_377),
.A3(n_373),
.B(n_369),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_397),
.A2(n_366),
.B(n_356),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_405),
.A2(n_386),
.B(n_384),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_363),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_379),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_354),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_394),
.Y(n_426)
);

AO22x1_ASAP7_75t_L g427 ( 
.A1(n_418),
.A2(n_354),
.B1(n_350),
.B2(n_372),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_374),
.B1(n_372),
.B2(n_370),
.Y(n_428)
);

CKINVDCx8_ASAP7_75t_R g429 ( 
.A(n_416),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_414),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_R g432 ( 
.A(n_394),
.B(n_342),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_350),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_83),
.Y(n_435)
);

AOI21x1_ASAP7_75t_L g436 ( 
.A1(n_412),
.A2(n_374),
.B(n_378),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_84),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_406),
.A2(n_378),
.B(n_370),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_396),
.A2(n_362),
.B1(n_90),
.B2(n_93),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_88),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_362),
.B(n_95),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_402),
.Y(n_442)
);

NAND3x1_ASAP7_75t_L g443 ( 
.A(n_388),
.B(n_94),
.C(n_97),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_100),
.C(n_105),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g445 ( 
.A1(n_421),
.A2(n_398),
.B(n_417),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_420),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_430),
.A2(n_411),
.B(n_410),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_423),
.A2(n_408),
.B(n_407),
.C(n_399),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

AO21x2_ASAP7_75t_L g451 ( 
.A1(n_441),
.A2(n_106),
.B(n_109),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_110),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

BUFx12f_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_428),
.A2(n_111),
.B1(n_113),
.B2(n_117),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_437),
.A2(n_123),
.B(n_124),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

AOI221xp5_ASAP7_75t_L g461 ( 
.A1(n_427),
.A2(n_439),
.B1(n_438),
.B2(n_444),
.C(n_440),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_432),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_435),
.A2(n_422),
.B1(n_424),
.B2(n_443),
.Y(n_463)
);

INVx8_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_436),
.Y(n_465)
);

AO21x2_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_405),
.B(n_361),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_467),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_467),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_449),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

AO21x2_ASAP7_75t_L g480 ( 
.A1(n_445),
.A2(n_466),
.B(n_458),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_464),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_466),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_451),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_452),
.Y(n_486)
);

NOR2x1_ASAP7_75t_SL g487 ( 
.A(n_454),
.B(n_457),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_463),
.B(n_448),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

AOI21x1_ASAP7_75t_L g493 ( 
.A1(n_461),
.A2(n_463),
.B(n_456),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_462),
.A2(n_429),
.B1(n_375),
.B2(n_461),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_449),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_496),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_472),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_R g500 ( 
.A(n_489),
.B(n_486),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_489),
.B(n_468),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_481),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_482),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_R g504 ( 
.A(n_496),
.B(n_493),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_R g505 ( 
.A(n_468),
.B(n_495),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_475),
.B(n_491),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_494),
.B(n_488),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_469),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_493),
.B(n_492),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_474),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_478),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_R g513 ( 
.A(n_490),
.B(n_479),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_471),
.B(n_490),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_471),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_482),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_476),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_484),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_480),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_517),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_515),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_505),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_508),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_502),
.B(n_470),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_514),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_483),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_502),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_484),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_483),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_511),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_512),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_521),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_523),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_516),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_500),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_533),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_497),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_522),
.B(n_501),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_532),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_537),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_534),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_538),
.B(n_527),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_536),
.B(n_530),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_534),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_529),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_541),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_543),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_535),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_524),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_537),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_553),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_549),
.B(n_542),
.Y(n_555)
);

AO21x2_ASAP7_75t_L g556 ( 
.A1(n_550),
.A2(n_543),
.B(n_504),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_551),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_552),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_557),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_542),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_537),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_560),
.B(n_555),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_558),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_562),
.Y(n_564)
);

AOI211x1_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_563),
.B(n_556),
.C(n_561),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_SL g566 ( 
.A(n_565),
.B(n_540),
.C(n_564),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_567),
.B(n_540),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_568),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_569),
.Y(n_570)
);

XNOR2x1_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_497),
.Y(n_571)
);

AOI31xp33_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_507),
.A3(n_513),
.B(n_531),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_539),
.Y(n_573)
);

XNOR2x1_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_539),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_573),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_511),
.B1(n_510),
.B2(n_525),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_575),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_576),
.Y(n_578)
);

OAI221xp5_ASAP7_75t_R g579 ( 
.A1(n_577),
.A2(n_520),
.B1(n_519),
.B2(n_480),
.C(n_526),
.Y(n_579)
);

AOI211xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_578),
.B(n_520),
.C(n_485),
.Y(n_580)
);


endmodule