module fake_jpeg_6811_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_62),
.B1(n_23),
.B2(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_33),
.B1(n_24),
.B2(n_17),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_64),
.Y(n_94)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_27),
.B1(n_29),
.B2(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_16),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_16),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_38),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_38),
.B1(n_35),
.B2(n_17),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_28),
.C(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_33),
.B1(n_23),
.B2(n_18),
.Y(n_85)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_43),
.B1(n_41),
.B2(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_87),
.B1(n_93),
.B2(n_50),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_43),
.B1(n_41),
.B2(n_29),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_92),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_47),
.B(n_61),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_64),
.B1(n_54),
.B2(n_66),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_48),
.B(n_23),
.C(n_65),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_38),
.B1(n_19),
.B2(n_23),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_74),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_82),
.B1(n_57),
.B2(n_50),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_38),
.B1(n_19),
.B2(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_96),
.Y(n_126)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_59),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_73),
.C(n_49),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_104),
.B1(n_114),
.B2(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_103),
.B1(n_48),
.B2(n_89),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_66),
.C(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_56),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_68),
.B(n_51),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_127),
.C(n_34),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_51),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_57),
.B1(n_46),
.B2(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_47),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_144)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_125),
.B1(n_114),
.B2(n_127),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_91),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_34),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_23),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_104),
.B1(n_110),
.B2(n_107),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_75),
.B1(n_79),
.B2(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_150),
.B1(n_152),
.B2(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_137),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_91),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_20),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_134),
.B(n_147),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_73),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_116),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_155),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_84),
.B1(n_95),
.B2(n_81),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_84),
.B1(n_81),
.B2(n_46),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_96),
.B1(n_60),
.B2(n_58),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_110),
.B1(n_135),
.B2(n_118),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_34),
.C(n_40),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_141),
.B(n_131),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_164),
.B(n_172),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_120),
.B(n_112),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_146),
.B(n_143),
.C(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_170),
.B1(n_173),
.B2(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_167),
.B1(n_181),
.B2(n_19),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_106),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_101),
.B1(n_113),
.B2(n_121),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_113),
.B1(n_92),
.B2(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_175),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_34),
.B(n_40),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_40),
.B(n_25),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_152),
.B1(n_129),
.B2(n_144),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_34),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_145),
.C(n_137),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_140),
.B1(n_154),
.B2(n_141),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_184),
.B(n_185),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_195),
.C(n_200),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_133),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_199),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_140),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_205),
.B(n_174),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_191),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_180),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_40),
.C(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_92),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_18),
.C(n_25),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_159),
.B(n_166),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_158),
.B1(n_18),
.B2(n_25),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_25),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_25),
.C(n_20),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_172),
.C(n_171),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_167),
.B1(n_177),
.B2(n_165),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_219),
.B1(n_230),
.B2(n_235),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_165),
.B1(n_181),
.B2(n_166),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_186),
.C(n_210),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_188),
.A2(n_158),
.B1(n_164),
.B2(n_168),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_191),
.B1(n_209),
.B2(n_197),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_20),
.B1(n_18),
.B2(n_22),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_20),
.B1(n_18),
.B2(n_22),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_212),
.B1(n_234),
.B2(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_236),
.B(n_0),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_22),
.B(n_1),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_195),
.C(n_189),
.Y(n_237)
);

AOI221xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_236),
.B1(n_216),
.B2(n_228),
.C(n_221),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_245),
.C(n_251),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_201),
.B(n_191),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_247),
.B1(n_249),
.B2(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_246),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_224),
.C(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_213),
.B(n_189),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_193),
.C(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_258),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_216),
.A2(n_197),
.B1(n_15),
.B2(n_13),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_0),
.C(n_1),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_257),
.C(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_213),
.B(n_2),
.CI(n_3),
.CON(n_258),
.SN(n_258)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_276),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_250),
.B(n_245),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_259),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_270),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_221),
.B1(n_220),
.B2(n_233),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_251),
.B1(n_250),
.B2(n_239),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_3),
.C(n_4),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_4),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_284),
.B(n_289),
.Y(n_299)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_267),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_248),
.B1(n_238),
.B2(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_258),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_273),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_5),
.B(n_6),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_294),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_272),
.B1(n_268),
.B2(n_275),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_282),
.B1(n_293),
.B2(n_285),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_260),
.B(n_269),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_300),
.B(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_260),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_303),
.C(n_306),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_261),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_273),
.B(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_276),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_288),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_309),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_290),
.C(n_6),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_303),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_10),
.B1(n_13),
.B2(n_11),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_10),
.B1(n_15),
.B2(n_8),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_10),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_302),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_304),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_323),
.B(n_325),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_306),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_312),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_311),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_312),
.B(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_314),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.C(n_15),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_5),
.B(n_7),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_330),
.B(n_329),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_335),
.C(n_8),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_7),
.B(n_8),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.C(n_324),
.Y(n_339)
);


endmodule