module fake_jpeg_10534_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_19),
.B1(n_22),
.B2(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_53),
.B1(n_18),
.B2(n_21),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_21),
.B1(n_34),
.B2(n_23),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.C(n_37),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_43),
.C(n_44),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_19),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_62),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_1),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_17),
.B1(n_22),
.B2(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_63),
.B1(n_31),
.B2(n_25),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_34),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_34),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_75),
.B(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_67),
.Y(n_103)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_83),
.B1(n_23),
.B2(n_34),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_71),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_23),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_27),
.B1(n_31),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_79),
.B1(n_3),
.B2(n_5),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_84),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_27),
.B1(n_25),
.B2(n_18),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_52),
.B1(n_62),
.B2(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_85),
.B1(n_92),
.B2(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_86),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_42),
.C(n_34),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_61),
.B1(n_47),
.B2(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_23),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_42),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_105),
.B1(n_70),
.B2(n_95),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_44),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_100),
.B(n_42),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_41),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_3),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_80),
.B1(n_79),
.B2(n_67),
.Y(n_126)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_42),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_119),
.B(n_112),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_130),
.B(n_133),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_121),
.B1(n_117),
.B2(n_97),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_85),
.B1(n_96),
.B2(n_91),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_141),
.B1(n_145),
.B2(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_136),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_135),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_77),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_5),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_148),
.B(n_129),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_90),
.B1(n_66),
.B2(n_84),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_121),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_15),
.C(n_6),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_14),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_14),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_7),
.B(n_8),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_118),
.B(n_116),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_152),
.B(n_168),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_118),
.B(n_97),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_161),
.B1(n_170),
.B2(n_172),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_127),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_99),
.B1(n_120),
.B2(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_108),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_99),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_143),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_100),
.B(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_173),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_109),
.B1(n_108),
.B2(n_9),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_129),
.B(n_7),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_125),
.B(n_130),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_8),
.B(n_11),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_140),
.C(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_173),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_134),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_182),
.C(n_186),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_141),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_140),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_137),
.C(n_149),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_189),
.C(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_145),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_172),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_109),
.B(n_9),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_156),
.B(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_166),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_203),
.C(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_163),
.B1(n_161),
.B2(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_168),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_184),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_208),
.B(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_207),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_202),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_162),
.C(n_150),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_180),
.B(n_184),
.Y(n_217)
);

AOI321xp33_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_156),
.A3(n_109),
.B1(n_11),
.B2(n_12),
.C(n_10),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_208),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_109),
.B1(n_10),
.B2(n_11),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_218),
.C(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_181),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_220),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_179),
.C(n_185),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_230),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_194),
.B(n_205),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_227),
.B(n_229),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_190),
.B1(n_193),
.B2(n_183),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_196),
.B1(n_193),
.B2(n_202),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_175),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_192),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_226),
.B(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_175),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_220),
.C(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_237),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_204),
.B(n_179),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_241),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_195),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_206),
.Y(n_241)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_232),
.B(n_229),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_218),
.B1(n_189),
.B2(n_12),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_239),
.A2(n_234),
.B(n_228),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_243),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_247),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_12),
.Y(n_251)
);


endmodule