module fake_jpeg_25998_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_42),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.C(n_1),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_34),
.C(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_8),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_27),
.B1(n_21),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_34),
.B1(n_21),
.B2(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_62),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_27),
.B1(n_33),
.B2(n_17),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_64),
.B1(n_40),
.B2(n_27),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_51),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_42),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_21),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_57),
.B(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_58),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_29),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_27),
.B1(n_30),
.B2(n_22),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_40),
.B1(n_41),
.B2(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_79),
.B1(n_86),
.B2(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_63),
.B1(n_60),
.B2(n_46),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_79),
.B(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_84),
.Y(n_98)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_19),
.B1(n_30),
.B2(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_19),
.B1(n_18),
.B2(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_18),
.B1(n_32),
.B2(n_31),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_56),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_38),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_56),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_47),
.C(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_70),
.C(n_90),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_49),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_20),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_56),
.B1(n_63),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_112),
.B1(n_118),
.B2(n_72),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_113),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_63),
.B1(n_60),
.B2(n_29),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_0),
.B(n_1),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_0),
.B(n_1),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_68),
.B1(n_74),
.B2(n_84),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_25),
.Y(n_119)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_123),
.B1(n_127),
.B2(n_145),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_65),
.B1(n_71),
.B2(n_67),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_142),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_134),
.B(n_138),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_66),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_143),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_107),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_66),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_137),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_23),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_110),
.B1(n_113),
.B2(n_75),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_23),
.C(n_25),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_117),
.C(n_118),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_87),
.B1(n_20),
.B2(n_75),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_46),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_104),
.B1(n_115),
.B2(n_109),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_149),
.B1(n_76),
.B2(n_77),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_109),
.B1(n_107),
.B2(n_112),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_99),
.B(n_112),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_173),
.B(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_163),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_160),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_97),
.C(n_99),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_166),
.C(n_170),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_129),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_118),
.B1(n_106),
.B2(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_165),
.B1(n_131),
.B2(n_143),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_100),
.B1(n_103),
.B2(n_119),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_103),
.C(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_11),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_96),
.C(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_114),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_23),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_23),
.B(n_76),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_186),
.C(n_158),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_192),
.B(n_164),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_200),
.B1(n_149),
.B2(n_173),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_193),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_144),
.C(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_R g191 ( 
.A(n_150),
.B(n_134),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_153),
.B(n_3),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_132),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_157),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_154),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_10),
.B1(n_13),
.B2(n_6),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_77),
.B1(n_76),
.B2(n_5),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_205),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_210),
.B1(n_212),
.B2(n_216),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_167),
.C(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_163),
.C(n_162),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_170),
.C(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_172),
.C(n_165),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_218),
.C(n_219),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_153),
.B1(n_77),
.B2(n_2),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_10),
.A3(n_14),
.B1(n_6),
.B2(n_7),
.C1(n_9),
.C2(n_15),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_181),
.A3(n_200),
.B1(n_184),
.B2(n_183),
.C1(n_15),
.C2(n_12),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_9),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_10),
.C(n_12),
.Y(n_219)
);

OA21x2_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_6),
.B(n_7),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_236),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_227),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_184),
.B1(n_190),
.B2(n_188),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_193),
.B1(n_219),
.B2(n_218),
.Y(n_247)
);

NAND4xp25_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_212),
.C(n_216),
.D(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_177),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_197),
.C(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_208),
.C(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_238),
.C(n_248),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_204),
.C(n_201),
.Y(n_238)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_229),
.Y(n_250)
);

HB1xp67_ASAP7_75t_SL g252 ( 
.A(n_242),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_211),
.B1(n_187),
.B2(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_195),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_226),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_231),
.B(n_233),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_11),
.C(n_12),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_258),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_229),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_15),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_2),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_262),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_241),
.B1(n_239),
.B2(n_246),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_249),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_252),
.A2(n_240),
.B(n_248),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_238),
.B(n_3),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_3),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_268),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_254),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_270),
.B(n_260),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_271),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_273),
.A2(n_259),
.B1(n_253),
.B2(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_272),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_275),
.Y(n_277)
);


endmodule