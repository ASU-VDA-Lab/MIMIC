module real_aes_16918_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_2000, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_2000;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1441;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_1250;
wire n_1987;
wire n_859;
wire n_1465;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_1632;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_1945;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_1951;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_1971;
wire n_964;
wire n_731;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1671;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1691;
wire n_1176;
wire n_1931;
wire n_640;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1584;
wire n_466;
wire n_1277;
wire n_1049;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_1647;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1972 ( .A1(n_0), .A2(n_108), .B1(n_576), .B2(n_694), .C(n_1018), .Y(n_1972) );
AOI22xp33_ASAP7_75t_SL g1984 ( .A1(n_0), .A2(n_237), .B1(n_1375), .B2(n_1985), .Y(n_1984) );
AOI22xp33_ASAP7_75t_L g1699 ( .A1(n_1), .A2(n_92), .B1(n_1691), .B2(n_1694), .Y(n_1699) );
AOI22xp33_ASAP7_75t_L g1649 ( .A1(n_2), .A2(n_292), .B1(n_1028), .B2(n_1381), .Y(n_1649) );
AOI22xp33_ASAP7_75t_L g1664 ( .A1(n_2), .A2(n_251), .B1(n_525), .B2(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1180 ( .A(n_3), .Y(n_1180) );
INVx1_ASAP7_75t_L g389 ( .A(n_4), .Y(n_389) );
AND2x2_ASAP7_75t_L g417 ( .A(n_4), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g533 ( .A(n_4), .B(n_258), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_4), .B(n_399), .Y(n_559) );
INVx1_ASAP7_75t_L g1010 ( .A(n_5), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_5), .A2(n_85), .B1(n_439), .B2(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1122 ( .A(n_6), .Y(n_1122) );
INVx1_ASAP7_75t_L g1964 ( .A(n_7), .Y(n_1964) );
OAI22xp33_ASAP7_75t_L g1989 ( .A1(n_7), .A2(n_96), .B1(n_1207), .B2(n_1990), .Y(n_1989) );
INVx1_ASAP7_75t_L g998 ( .A(n_8), .Y(n_998) );
INVx1_ASAP7_75t_L g727 ( .A(n_9), .Y(n_727) );
OA222x2_ASAP7_75t_L g749 ( .A1(n_9), .A2(n_144), .B1(n_175), .B2(n_750), .C1(n_752), .C2(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g1422 ( .A(n_10), .Y(n_1422) );
OAI211xp5_ASAP7_75t_SL g1546 ( .A1(n_11), .A2(n_1038), .B(n_1547), .C(n_1550), .Y(n_1546) );
INVx1_ASAP7_75t_L g1570 ( .A(n_11), .Y(n_1570) );
AOI22xp33_ASAP7_75t_SL g1650 ( .A1(n_12), .A2(n_210), .B1(n_708), .B2(n_742), .Y(n_1650) );
AOI221xp5_ASAP7_75t_L g1663 ( .A1(n_12), .A2(n_117), .B1(n_546), .B2(n_666), .C(n_759), .Y(n_1663) );
AOI221xp5_ASAP7_75t_L g1380 ( .A1(n_13), .A2(n_30), .B1(n_967), .B2(n_1381), .C(n_1382), .Y(n_1380) );
INVx1_ASAP7_75t_L g1400 ( .A(n_13), .Y(n_1400) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_14), .A2(n_370), .B1(n_439), .B2(n_444), .C(n_450), .Y(n_1049) );
OAI21xp33_ASAP7_75t_SL g1077 ( .A1(n_14), .A2(n_595), .B(n_753), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_15), .A2(n_73), .B1(n_712), .B2(n_934), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_15), .A2(n_335), .B1(n_1017), .B2(n_1308), .C(n_1309), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1958 ( .A1(n_16), .A2(n_95), .B1(n_576), .B2(n_1174), .C(n_1249), .Y(n_1958) );
AOI22xp33_ASAP7_75t_SL g1988 ( .A1(n_16), .A2(n_200), .B1(n_479), .B2(n_638), .Y(n_1988) );
INVx2_ASAP7_75t_L g434 ( .A(n_17), .Y(n_434) );
INVx1_ASAP7_75t_L g1179 ( .A(n_18), .Y(n_1179) );
OAI322xp33_ASAP7_75t_L g1181 ( .A1(n_18), .A2(n_1182), .A3(n_1188), .B1(n_1189), .B2(n_1193), .C1(n_1198), .C2(n_1201), .Y(n_1181) );
INVxp67_ASAP7_75t_SL g1409 ( .A(n_19), .Y(n_1409) );
OAI211xp5_ASAP7_75t_L g1441 ( .A1(n_19), .A2(n_450), .B(n_1038), .C(n_1442), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_20), .A2(n_177), .B1(n_709), .B2(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_20), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g1171 ( .A1(n_21), .A2(n_235), .B1(n_761), .B2(n_1172), .C(n_1174), .Y(n_1171) );
INVx1_ASAP7_75t_L g1191 ( .A(n_21), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_22), .A2(n_303), .B1(n_487), .B2(n_490), .Y(n_1060) );
INVx1_ASAP7_75t_L g1076 ( .A(n_22), .Y(n_1076) );
INVx1_ASAP7_75t_L g1598 ( .A(n_23), .Y(n_1598) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_24), .A2(n_369), .B1(n_619), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_24), .A2(n_158), .B1(n_579), .B2(n_580), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_25), .Y(n_1279) );
INVx1_ASAP7_75t_L g1411 ( .A(n_26), .Y(n_1411) );
XOR2x1_ASAP7_75t_L g408 ( .A(n_27), .B(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_28), .A2(n_339), .B1(n_487), .B2(n_490), .Y(n_1123) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_28), .Y(n_1125) );
INVx1_ASAP7_75t_L g968 ( .A(n_29), .Y(n_968) );
AOI221x1_ASAP7_75t_SL g973 ( .A1(n_29), .A2(n_198), .B1(n_525), .B2(n_885), .C(n_974), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g1392 ( .A1(n_30), .A2(n_152), .B1(n_661), .B2(n_692), .C(n_1393), .Y(n_1392) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_31), .Y(n_384) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_31), .B(n_382), .Y(n_1685) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_32), .A2(n_229), .B1(n_628), .B2(n_722), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_32), .A2(n_314), .B1(n_779), .B2(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_33), .A2(n_313), .B1(n_983), .B2(n_1176), .Y(n_1175) );
INVxp67_ASAP7_75t_L g1186 ( .A(n_33), .Y(n_1186) );
INVx1_ASAP7_75t_L g1924 ( .A(n_34), .Y(n_1924) );
INVx1_ASAP7_75t_L g962 ( .A(n_35), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_35), .A2(n_181), .B1(n_547), .B2(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g1225 ( .A(n_36), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_36), .A2(n_66), .B1(n_987), .B2(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1153 ( .A(n_37), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_38), .A2(n_273), .B1(n_456), .B2(n_463), .Y(n_455) );
INVxp33_ASAP7_75t_L g593 ( .A(n_38), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_39), .A2(n_333), .B1(n_487), .B2(n_490), .Y(n_1379) );
INVxp67_ASAP7_75t_SL g1403 ( .A(n_39), .Y(n_1403) );
OAI211xp5_ASAP7_75t_SL g1594 ( .A1(n_40), .A2(n_1595), .B(n_1597), .C(n_1600), .Y(n_1594) );
OAI22xp5_ASAP7_75t_L g1631 ( .A1(n_40), .A2(n_291), .B1(n_649), .B2(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g1115 ( .A(n_41), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_42), .A2(n_311), .B1(n_983), .B2(n_1165), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_42), .A2(n_235), .B1(n_479), .B2(n_711), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1697 ( .A1(n_43), .A2(n_70), .B1(n_1684), .B2(n_1698), .Y(n_1697) );
AOI22xp33_ASAP7_75t_L g1648 ( .A1(n_44), .A2(n_251), .B1(n_1028), .B2(n_1381), .Y(n_1648) );
AOI221xp5_ASAP7_75t_L g1660 ( .A1(n_44), .A2(n_292), .B1(n_577), .B2(n_888), .C(n_1088), .Y(n_1660) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_45), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_45), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_46), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_47), .A2(n_288), .B1(n_706), .B2(n_709), .Y(n_705) );
INVxp67_ASAP7_75t_SL g763 ( .A(n_47), .Y(n_763) );
AOI22xp33_ASAP7_75t_SL g1565 ( .A1(n_48), .A2(n_245), .B1(n_502), .B2(n_722), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_48), .A2(n_286), .B1(n_779), .B2(n_847), .Y(n_1579) );
CKINVDCx5p33_ASAP7_75t_R g1641 ( .A(n_49), .Y(n_1641) );
OAI221xp5_ASAP7_75t_L g1603 ( .A1(n_50), .A2(n_118), .B1(n_680), .B2(n_1604), .C(n_1605), .Y(n_1603) );
OAI22xp33_ASAP7_75t_L g1624 ( .A1(n_50), .A2(n_118), .B1(n_1625), .B2(n_1627), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_51), .A2(n_193), .B1(n_525), .B2(n_778), .Y(n_889) );
INVx1_ASAP7_75t_L g924 ( .A(n_51), .Y(n_924) );
INVx1_ASAP7_75t_L g1369 ( .A(n_52), .Y(n_1369) );
INVx1_ASAP7_75t_L g1102 ( .A(n_53), .Y(n_1102) );
AOI22xp33_ASAP7_75t_SL g1609 ( .A1(n_54), .A2(n_265), .B1(n_1610), .B2(n_1611), .Y(n_1609) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_54), .A2(n_371), .B1(n_479), .B2(n_639), .Y(n_1619) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_55), .A2(n_124), .B1(n_614), .B2(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_55), .Y(n_690) );
INVx1_ASAP7_75t_L g1424 ( .A(n_56), .Y(n_1424) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_57), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g1241 ( .A1(n_58), .A2(n_351), .B1(n_721), .B2(n_724), .C(n_1242), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_58), .A2(n_168), .B1(n_1017), .B2(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1929 ( .A(n_59), .Y(n_1929) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_60), .A2(n_479), .B(n_724), .Y(n_1107) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_60), .Y(n_1134) );
INVx1_ASAP7_75t_L g1654 ( .A(n_61), .Y(n_1654) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_62), .A2(n_199), .B1(n_456), .B2(n_463), .Y(n_1222) );
CKINVDCx5p33_ASAP7_75t_R g1255 ( .A(n_62), .Y(n_1255) );
INVx1_ASAP7_75t_L g1504 ( .A(n_63), .Y(n_1504) );
OAI211xp5_ASAP7_75t_L g1516 ( .A1(n_63), .A2(n_1517), .B(n_1519), .C(n_1521), .Y(n_1516) );
AOI22xp5_ASAP7_75t_L g1710 ( .A1(n_64), .A2(n_111), .B1(n_1684), .B2(n_1698), .Y(n_1710) );
AOI22xp5_ASAP7_75t_L g1717 ( .A1(n_65), .A2(n_263), .B1(n_1684), .B2(n_1698), .Y(n_1717) );
INVx1_ASAP7_75t_L g1245 ( .A(n_66), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_67), .A2(n_221), .B1(n_839), .B2(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g918 ( .A(n_67), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_68), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1103 ( .A1(n_69), .A2(n_261), .B1(n_439), .B2(n_444), .C(n_450), .Y(n_1103) );
OAI221xp5_ASAP7_75t_L g1147 ( .A1(n_69), .A2(n_339), .B1(n_595), .B2(n_985), .C(n_987), .Y(n_1147) );
OAI21xp5_ASAP7_75t_L g1427 ( .A1(n_71), .A2(n_1266), .B(n_1428), .Y(n_1427) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_71), .A2(n_78), .B1(n_456), .B2(n_463), .Y(n_1429) );
INVx1_ASAP7_75t_L g1406 ( .A(n_72), .Y(n_1406) );
AOI22xp33_ASAP7_75t_SL g1305 ( .A1(n_73), .A2(n_143), .B1(n_579), .B2(n_580), .Y(n_1305) );
AOI21xp33_ASAP7_75t_L g1061 ( .A1(n_74), .A2(n_1062), .B(n_1065), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_74), .A2(n_107), .B1(n_576), .B2(n_1087), .C(n_1089), .Y(n_1086) );
INVx1_ASAP7_75t_L g789 ( .A(n_75), .Y(n_789) );
INVx1_ASAP7_75t_L g1226 ( .A(n_76), .Y(n_1226) );
OAI21xp33_ASAP7_75t_L g1270 ( .A1(n_76), .A2(n_595), .B(n_753), .Y(n_1270) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_77), .Y(n_1205) );
INVxp33_ASAP7_75t_L g1426 ( .A(n_78), .Y(n_1426) );
INVx1_ASAP7_75t_L g1167 ( .A(n_79), .Y(n_1167) );
OAI211xp5_ASAP7_75t_L g1206 ( .A1(n_79), .A2(n_1207), .B(n_1210), .C(n_1213), .Y(n_1206) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_80), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g1727 ( .A1(n_81), .A2(n_247), .B1(n_1684), .B2(n_1698), .Y(n_1727) );
XOR2x2_ASAP7_75t_L g1887 ( .A(n_81), .B(n_1888), .Y(n_1887) );
AOI22xp33_ASAP7_75t_L g1944 ( .A1(n_81), .A2(n_1945), .B1(n_1948), .B2(n_1993), .Y(n_1944) );
INVx1_ASAP7_75t_L g612 ( .A(n_82), .Y(n_612) );
AOI21xp33_ASAP7_75t_L g1608 ( .A1(n_83), .A2(n_693), .B(n_694), .Y(n_1608) );
INVx1_ASAP7_75t_L g1615 ( .A(n_83), .Y(n_1615) );
XOR2x2_ASAP7_75t_L g1044 ( .A(n_84), .B(n_1045), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1703 ( .A1(n_84), .A2(n_256), .B1(n_1691), .B2(n_1694), .Y(n_1703) );
INVx1_ASAP7_75t_L g1003 ( .A(n_85), .Y(n_1003) );
AOI22xp5_ASAP7_75t_L g1704 ( .A1(n_86), .A2(n_104), .B1(n_1684), .B2(n_1705), .Y(n_1704) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_87), .B(n_600), .Y(n_599) );
AO22x1_ASAP7_75t_L g1690 ( .A1(n_87), .A2(n_266), .B1(n_1691), .B2(n_1694), .Y(n_1690) );
INVx1_ASAP7_75t_L g1892 ( .A(n_88), .Y(n_1892) );
OAI221xp5_ASAP7_75t_L g867 ( .A1(n_89), .A2(n_123), .B1(n_764), .B2(n_868), .C(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g898 ( .A(n_89), .Y(n_898) );
CKINVDCx5p33_ASAP7_75t_R g1231 ( .A(n_90), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_91), .A2(n_201), .B1(n_487), .B2(n_490), .Y(n_486) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_91), .Y(n_543) );
XOR2xp5_ASAP7_75t_L g1637 ( .A(n_92), .B(n_1638), .Y(n_1637) );
OAI22xp5_ASAP7_75t_L g1976 ( .A1(n_93), .A2(n_206), .B1(n_647), .B2(n_649), .Y(n_1976) );
INVx1_ASAP7_75t_L g871 ( .A(n_94), .Y(n_871) );
OAI221xp5_ASAP7_75t_SL g906 ( .A1(n_94), .A2(n_121), .B1(n_442), .B2(n_610), .C(n_814), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g1983 ( .A1(n_95), .A2(n_290), .B1(n_638), .B2(n_1374), .Y(n_1983) );
INVx1_ASAP7_75t_L g1962 ( .A(n_96), .Y(n_1962) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_97), .A2(n_344), .B1(n_934), .B2(n_1235), .C(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1359 ( .A(n_97), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_98), .A2(n_215), .B1(n_456), .B2(n_463), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1085 ( .A(n_98), .Y(n_1085) );
AND2x2_ASAP7_75t_L g484 ( .A(n_99), .B(n_485), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_99), .A2(n_226), .B1(n_579), .B2(n_580), .C(n_582), .Y(n_578) );
INVx1_ASAP7_75t_L g1668 ( .A(n_100), .Y(n_1668) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_101), .A2(n_116), .B1(n_721), .B2(n_722), .C(n_724), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_101), .A2(n_288), .B1(n_778), .B2(n_779), .Y(n_777) );
AOI222xp33_ASAP7_75t_L g1066 ( .A1(n_102), .A2(n_148), .B1(n_354), .B2(n_465), .C1(n_619), .C2(n_961), .Y(n_1066) );
INVx1_ASAP7_75t_L g1091 ( .A(n_102), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_103), .B(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_103), .A2(n_174), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_105), .A2(n_196), .B1(n_624), .B2(n_625), .Y(n_623) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_105), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g1373 ( .A1(n_106), .A2(n_319), .B1(n_1374), .B2(n_1375), .C(n_1376), .Y(n_1373) );
INVx1_ASAP7_75t_L g1394 ( .A(n_106), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_107), .A2(n_228), .B1(n_1053), .B2(n_1055), .C(n_1057), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1987 ( .A1(n_108), .A2(n_294), .B1(n_628), .B2(n_631), .Y(n_1987) );
INVx1_ASAP7_75t_L g382 ( .A(n_109), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g1458 ( .A(n_110), .Y(n_1458) );
INVx1_ASAP7_75t_L g1541 ( .A(n_112), .Y(n_1541) );
AO221x2_ASAP7_75t_L g1769 ( .A1(n_112), .A2(n_355), .B1(n_1691), .B2(n_1694), .C(n_1770), .Y(n_1769) );
AOI221xp5_ASAP7_75t_L g890 ( .A1(n_113), .A2(n_150), .B1(n_761), .B2(n_885), .C(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g912 ( .A(n_113), .Y(n_912) );
INVx1_ASAP7_75t_L g1048 ( .A(n_114), .Y(n_1048) );
OAI21xp33_ASAP7_75t_L g1073 ( .A1(n_114), .A2(n_520), .B(n_1074), .Y(n_1073) );
OAI211xp5_ASAP7_75t_L g1890 ( .A1(n_115), .A2(n_1140), .B(n_1495), .C(n_1891), .Y(n_1890) );
INVx1_ASAP7_75t_L g1913 ( .A(n_115), .Y(n_1913) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_116), .A2(n_155), .B1(n_759), .B2(n_761), .C(n_762), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g1645 ( .A1(n_117), .A2(n_257), .B1(n_1646), .B2(n_1647), .Y(n_1645) );
XOR2x2_ASAP7_75t_L g1316 ( .A(n_119), .B(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1567 ( .A(n_120), .Y(n_1567) );
INVx1_ASAP7_75t_L g880 ( .A(n_121), .Y(n_880) );
INVx1_ASAP7_75t_L g937 ( .A(n_122), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_122), .A2(n_253), .B1(n_985), .B2(n_987), .Y(n_984) );
INVx1_ASAP7_75t_L g896 ( .A(n_123), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_124), .A2(n_196), .B1(n_659), .B2(n_664), .C(n_666), .Y(n_658) );
INVx1_ASAP7_75t_L g1330 ( .A(n_125), .Y(n_1330) );
INVx1_ASAP7_75t_L g1335 ( .A(n_126), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1602 ( .A1(n_127), .A2(n_241), .B1(n_580), .B2(n_779), .Y(n_1602) );
INVx1_ASAP7_75t_L g1618 ( .A(n_127), .Y(n_1618) );
INVx1_ASAP7_75t_L g1932 ( .A(n_128), .Y(n_1932) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_129), .A2(n_786), .B1(n_787), .B2(n_855), .Y(n_785) );
INVx1_ASAP7_75t_L g855 ( .A(n_129), .Y(n_855) );
INVx1_ASAP7_75t_L g1334 ( .A(n_130), .Y(n_1334) );
INVx1_ASAP7_75t_L g875 ( .A(n_131), .Y(n_875) );
OAI21xp33_ASAP7_75t_L g904 ( .A1(n_131), .A2(n_642), .B(n_905), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_132), .Y(n_1280) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_133), .A2(n_332), .B1(n_439), .B2(n_444), .C(n_450), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_133), .B(n_551), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_134), .A2(n_204), .B1(n_487), .B2(n_490), .Y(n_1331) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_134), .A2(n_299), .B1(n_530), .B2(n_539), .Y(n_1345) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_135), .A2(n_269), .B1(n_779), .B2(n_893), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_135), .A2(n_353), .B1(n_479), .B2(n_721), .C(n_724), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1895 ( .A1(n_136), .A2(n_349), .B1(n_1896), .B2(n_1897), .Y(n_1895) );
OAI22xp5_ASAP7_75t_L g1904 ( .A1(n_136), .A2(n_349), .B1(n_1905), .B2(n_1906), .Y(n_1904) );
INVx1_ASAP7_75t_L g1166 ( .A(n_137), .Y(n_1166) );
AOI22xp33_ASAP7_75t_SL g1286 ( .A1(n_138), .A2(n_318), .B1(n_1287), .B2(n_1289), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_138), .A2(n_305), .B1(n_579), .B2(n_580), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1322 ( .A1(n_139), .A2(n_225), .B1(n_456), .B2(n_463), .Y(n_1322) );
INVxp67_ASAP7_75t_SL g1343 ( .A(n_139), .Y(n_1343) );
AO22x1_ASAP7_75t_L g1714 ( .A1(n_140), .A2(n_361), .B1(n_1691), .B2(n_1694), .Y(n_1714) );
OAI22xp33_ASAP7_75t_L g1899 ( .A1(n_141), .A2(n_173), .B1(n_1900), .B2(n_1901), .Y(n_1899) );
OAI22xp33_ASAP7_75t_L g1914 ( .A1(n_141), .A2(n_173), .B1(n_1512), .B2(n_1915), .Y(n_1914) );
INVx1_ASAP7_75t_L g1552 ( .A(n_142), .Y(n_1552) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_143), .A2(n_335), .B1(n_485), .B2(n_619), .Y(n_1291) );
INVx1_ASAP7_75t_L g743 ( .A(n_144), .Y(n_743) );
AOI221xp5_ASAP7_75t_SL g884 ( .A1(n_145), .A2(n_331), .B1(n_761), .B2(n_885), .C(n_888), .Y(n_884) );
INVx1_ASAP7_75t_L g921 ( .A(n_145), .Y(n_921) );
OAI222xp33_ASAP7_75t_L g640 ( .A1(n_146), .A2(n_252), .B1(n_262), .B2(n_641), .C1(n_647), .C2(n_649), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_146), .A2(n_654), .B(n_657), .C(n_669), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_147), .Y(n_882) );
INVx1_ASAP7_75t_L g1082 ( .A(n_148), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1160 ( .A1(n_149), .A2(n_214), .B1(n_546), .B2(n_1161), .C(n_1163), .Y(n_1160) );
INVxp67_ASAP7_75t_L g1183 ( .A(n_149), .Y(n_1183) );
INVx1_ASAP7_75t_L g925 ( .A(n_150), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g1601 ( .A1(n_151), .A2(n_371), .B1(n_563), .B2(n_891), .C(n_1308), .Y(n_1601) );
AOI22xp33_ASAP7_75t_L g1622 ( .A1(n_151), .A2(n_265), .B1(n_479), .B2(n_625), .Y(n_1622) );
INVx1_ASAP7_75t_L g1378 ( .A(n_152), .Y(n_1378) );
INVx1_ASAP7_75t_L g1232 ( .A(n_153), .Y(n_1232) );
AOI22xp33_ASAP7_75t_SL g1251 ( .A1(n_153), .A2(n_163), .B1(n_1252), .B2(n_1253), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_154), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_155), .A2(n_191), .B1(n_711), .B2(n_712), .C(n_715), .Y(n_710) );
AO22x1_ASAP7_75t_L g1683 ( .A1(n_156), .A2(n_362), .B1(n_1684), .B2(n_1688), .Y(n_1683) );
CKINVDCx16_ASAP7_75t_R g1771 ( .A(n_157), .Y(n_1771) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_158), .A2(n_368), .B1(n_631), .B2(n_633), .Y(n_630) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_159), .Y(n_794) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_159), .A2(n_450), .B1(n_456), .B2(n_811), .C(n_820), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_160), .A2(n_186), .B1(n_456), .B2(n_463), .Y(n_1371) );
INVxp67_ASAP7_75t_SL g1386 ( .A(n_160), .Y(n_1386) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_161), .A2(n_631), .B(n_715), .Y(n_808) );
INVx1_ASAP7_75t_L g835 ( .A(n_161), .Y(n_835) );
INVx1_ASAP7_75t_L g819 ( .A(n_162), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g837 ( .A1(n_162), .A2(n_229), .B1(n_838), .B2(n_839), .Y(n_837) );
INVx1_ASAP7_75t_L g1240 ( .A(n_163), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_164), .A2(n_373), .B1(n_465), .B2(n_723), .Y(n_1118) );
INVxp67_ASAP7_75t_SL g1144 ( .A(n_164), .Y(n_1144) );
INVx1_ASAP7_75t_L g1640 ( .A(n_165), .Y(n_1640) );
OAI221xp5_ASAP7_75t_L g1321 ( .A1(n_166), .A2(n_299), .B1(n_439), .B2(n_444), .C(n_450), .Y(n_1321) );
INVxp67_ASAP7_75t_SL g1341 ( .A(n_166), .Y(n_1341) );
INVx1_ASAP7_75t_L g1106 ( .A(n_167), .Y(n_1106) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_168), .A2(n_320), .B1(n_715), .B2(n_1234), .C(n_1235), .Y(n_1233) );
OAI22xp33_ASAP7_75t_L g1478 ( .A1(n_169), .A2(n_189), .B1(n_391), .B2(n_1479), .Y(n_1478) );
OAI22xp33_ASAP7_75t_L g1509 ( .A1(n_169), .A2(n_189), .B1(n_1510), .B2(n_1513), .Y(n_1509) );
INVx1_ASAP7_75t_L g1927 ( .A(n_170), .Y(n_1927) );
INVx1_ASAP7_75t_L g604 ( .A(n_171), .Y(n_604) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_171), .A2(n_183), .B1(n_676), .B2(n_680), .C(n_684), .Y(n_675) );
INVx1_ASAP7_75t_L g1894 ( .A(n_172), .Y(n_1894) );
OAI211xp5_ASAP7_75t_L g1907 ( .A1(n_172), .A2(n_1908), .B(n_1910), .C(n_1911), .Y(n_1907) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_174), .A2(n_209), .B1(n_494), .B2(n_499), .C(n_500), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_175), .A2(n_176), .B1(n_734), .B2(n_735), .C(n_739), .Y(n_733) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_176), .Y(n_755) );
INVxp33_ASAP7_75t_SL g765 ( .A(n_177), .Y(n_765) );
INVx1_ASAP7_75t_L g1549 ( .A(n_178), .Y(n_1549) );
INVx1_ASAP7_75t_L g437 ( .A(n_179), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_180), .Y(n_1500) );
INVx1_ASAP7_75t_L g952 ( .A(n_181), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g1415 ( .A1(n_182), .A2(n_264), .B1(n_885), .B2(n_1416), .C(n_1418), .Y(n_1415) );
INVx1_ASAP7_75t_L g1436 ( .A(n_182), .Y(n_1436) );
INVx1_ASAP7_75t_L g607 ( .A(n_183), .Y(n_607) );
INVx2_ASAP7_75t_L g1687 ( .A(n_184), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_184), .B(n_316), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_184), .B(n_1693), .Y(n_1695) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_185), .A2(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g566 ( .A(n_185), .Y(n_566) );
INVxp67_ASAP7_75t_SL g1401 ( .A(n_186), .Y(n_1401) );
CKINVDCx5p33_ASAP7_75t_R g1457 ( .A(n_187), .Y(n_1457) );
XNOR2xp5_ASAP7_75t_L g1591 ( .A(n_188), .B(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1656 ( .A(n_190), .Y(n_1656) );
INVx1_ASAP7_75t_L g773 ( .A(n_191), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g1000 ( .A1(n_192), .A2(n_750), .B(n_1001), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_192), .A2(n_301), .B1(n_823), .B2(n_1035), .C(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g911 ( .A(n_193), .Y(n_911) );
INVx1_ASAP7_75t_L g1113 ( .A(n_194), .Y(n_1113) );
OAI21xp5_ASAP7_75t_SL g1220 ( .A1(n_195), .A2(n_747), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1244 ( .A(n_195), .Y(n_1244) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_197), .Y(n_946) );
INVx1_ASAP7_75t_L g956 ( .A(n_198), .Y(n_956) );
INVx1_ASAP7_75t_L g1264 ( .A(n_199), .Y(n_1264) );
INVxp67_ASAP7_75t_SL g1971 ( .A(n_200), .Y(n_1971) );
INVx1_ASAP7_75t_L g410 ( .A(n_201), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_202), .A2(n_363), .B1(n_1017), .B2(n_1018), .Y(n_1413) );
AOI21xp33_ASAP7_75t_L g1438 ( .A1(n_202), .A2(n_715), .B(n_967), .Y(n_1438) );
CKINVDCx5p33_ASAP7_75t_R g1284 ( .A(n_203), .Y(n_1284) );
OAI211xp5_ASAP7_75t_L g1338 ( .A1(n_204), .A2(n_747), .B(n_1339), .C(n_1342), .Y(n_1338) );
INVx1_ASAP7_75t_L g741 ( .A(n_205), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_205), .A2(n_239), .B1(n_530), .B2(n_539), .Y(n_782) );
OAI211xp5_ASAP7_75t_L g1956 ( .A1(n_206), .A2(n_654), .B(n_1957), .C(n_1961), .Y(n_1956) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_207), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_208), .A2(n_340), .B1(n_575), .B2(n_887), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_208), .A2(n_234), .B1(n_715), .B2(n_721), .C(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g568 ( .A(n_209), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_210), .A2(n_257), .B1(n_779), .B2(n_893), .Y(n_1661) );
AOI22xp33_ASAP7_75t_SL g1293 ( .A1(n_211), .A2(n_305), .B1(n_614), .B2(n_1289), .Y(n_1293) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_211), .A2(n_318), .B1(n_576), .B2(n_666), .C(n_1302), .Y(n_1301) );
INVx2_ASAP7_75t_L g436 ( .A(n_212), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_212), .B(n_434), .Y(n_459) );
INVx1_ASAP7_75t_L g505 ( .A(n_212), .Y(n_505) );
INVx1_ASAP7_75t_L g1630 ( .A(n_213), .Y(n_1630) );
INVxp67_ASAP7_75t_L g1195 ( .A(n_214), .Y(n_1195) );
INVxp67_ASAP7_75t_SL g1069 ( .A(n_215), .Y(n_1069) );
OAI211xp5_ASAP7_75t_L g1223 ( .A1(n_216), .A2(n_450), .B(n_1038), .C(n_1224), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g1269 ( .A(n_216), .Y(n_1269) );
INVxp67_ASAP7_75t_SL g1563 ( .A(n_217), .Y(n_1563) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_217), .A2(n_222), .B1(n_1575), .B2(n_1577), .Y(n_1574) );
XOR2xp5_ASAP7_75t_L g927 ( .A(n_218), .B(n_928), .Y(n_927) );
OAI221xp5_ASAP7_75t_SL g1965 ( .A1(n_219), .A2(n_317), .B1(n_1966), .B2(n_1967), .C(n_1968), .Y(n_1965) );
INVx1_ASAP7_75t_L g1980 ( .A(n_219), .Y(n_1980) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_220), .A2(n_327), .B1(n_497), .B2(n_713), .Y(n_938) );
INVx1_ASAP7_75t_L g991 ( .A(n_220), .Y(n_991) );
INVx1_ASAP7_75t_L g922 ( .A(n_221), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g1558 ( .A1(n_222), .A2(n_310), .B1(n_724), .B2(n_1559), .C(n_1560), .Y(n_1558) );
CKINVDCx5p33_ASAP7_75t_R g1297 ( .A(n_223), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_224), .A2(n_352), .B1(n_893), .B2(n_1014), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_224), .A2(n_269), .B1(n_479), .B2(n_502), .Y(n_1026) );
INVxp67_ASAP7_75t_SL g1340 ( .A(n_225), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_226), .A2(n_282), .B1(n_472), .B2(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g428 ( .A(n_227), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_228), .B(n_692), .Y(n_1079) );
INVx1_ASAP7_75t_L g1058 ( .A(n_230), .Y(n_1058) );
OAI21xp5_ASAP7_75t_SL g1314 ( .A1(n_231), .A2(n_647), .B(n_1315), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1728 ( .A1(n_232), .A2(n_236), .B1(n_1691), .B2(n_1694), .Y(n_1728) );
INVx1_ASAP7_75t_L g1002 ( .A(n_233), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_234), .A2(n_353), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1959 ( .A1(n_237), .A2(n_294), .B1(n_1014), .B2(n_1960), .Y(n_1959) );
INVx1_ASAP7_75t_L g1921 ( .A(n_238), .Y(n_1921) );
INVx1_ASAP7_75t_L g726 ( .A(n_239), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g1452 ( .A(n_240), .Y(n_1452) );
INVx1_ASAP7_75t_L g1621 ( .A(n_241), .Y(n_1621) );
CKINVDCx5p33_ASAP7_75t_R g1975 ( .A(n_242), .Y(n_1975) );
INVx1_ASAP7_75t_L g1121 ( .A(n_243), .Y(n_1121) );
INVx1_ASAP7_75t_L g1568 ( .A(n_244), .Y(n_1568) );
OAI221xp5_ASAP7_75t_L g1572 ( .A1(n_244), .A2(n_330), .B1(n_987), .B2(n_1272), .C(n_1573), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_245), .A2(n_310), .B1(n_656), .B2(n_847), .Y(n_1584) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_246), .Y(n_793) );
OAI211xp5_ASAP7_75t_L g1492 ( .A1(n_248), .A2(n_1493), .B(n_1495), .C(n_1498), .Y(n_1492) );
INVx1_ASAP7_75t_L g1529 ( .A(n_248), .Y(n_1529) );
INVx1_ASAP7_75t_L g1328 ( .A(n_249), .Y(n_1328) );
INVx1_ASAP7_75t_L g469 ( .A(n_250), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_253), .A2(n_279), .B1(n_442), .B2(n_610), .C(n_913), .Y(n_942) );
INVx1_ASAP7_75t_L g1320 ( .A(n_254), .Y(n_1320) );
INVx1_ASAP7_75t_L g1599 ( .A(n_255), .Y(n_1599) );
BUFx3_ASAP7_75t_L g399 ( .A(n_258), .Y(n_399) );
INVx1_ASAP7_75t_L g418 ( .A(n_258), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g1773 ( .A(n_259), .Y(n_1773) );
AOI22xp5_ASAP7_75t_L g1716 ( .A1(n_260), .A2(n_283), .B1(n_1691), .B2(n_1694), .Y(n_1716) );
INVxp67_ASAP7_75t_SL g1149 ( .A(n_261), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1434 ( .A1(n_264), .A2(n_268), .B1(n_614), .B2(n_625), .C(n_724), .Y(n_1434) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_267), .A2(n_307), .B1(n_1483), .B2(n_1486), .Y(n_1482) );
OAI22xp33_ASAP7_75t_L g1530 ( .A1(n_267), .A2(n_307), .B1(n_1531), .B2(n_1533), .Y(n_1530) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_268), .A2(n_356), .B1(n_525), .B2(n_983), .Y(n_1414) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_270), .B(n_852), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_271), .Y(n_964) );
INVx1_ASAP7_75t_L g1555 ( .A(n_272), .Y(n_1555) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_273), .Y(n_511) );
INVxp67_ASAP7_75t_SL g994 ( .A(n_274), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_275), .Y(n_870) );
INVx1_ASAP7_75t_L g801 ( .A(n_276), .Y(n_801) );
INVx1_ASAP7_75t_L g1383 ( .A(n_277), .Y(n_1383) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_277), .A2(n_328), .B1(n_661), .B2(n_692), .C(n_1398), .Y(n_1397) );
AOI21xp33_ASAP7_75t_L g1564 ( .A1(n_278), .A2(n_619), .B(n_715), .Y(n_1564) );
INVx1_ASAP7_75t_L g1583 ( .A(n_278), .Y(n_1583) );
OA222x2_ASAP7_75t_L g988 ( .A1(n_279), .A2(n_298), .B1(n_357), .B2(n_520), .C1(n_750), .C2(n_753), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_280), .Y(n_1451) );
INVx1_ASAP7_75t_L g1923 ( .A(n_281), .Y(n_1923) );
AOI32xp33_ASAP7_75t_L g545 ( .A1(n_282), .A2(n_546), .A3(n_549), .B1(n_554), .B2(n_2000), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g1670 ( .A1(n_284), .A2(n_647), .B(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_L g1059 ( .A(n_285), .Y(n_1059) );
INVx1_ASAP7_75t_L g1557 ( .A(n_286), .Y(n_1557) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_287), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_289), .Y(n_1461) );
INVxp67_ASAP7_75t_SL g1969 ( .A(n_290), .Y(n_1969) );
AOI211xp5_ASAP7_75t_L g1324 ( .A1(n_293), .A2(n_721), .B(n_1325), .C(n_1327), .Y(n_1324) );
INVx1_ASAP7_75t_L g1355 ( .A(n_293), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1709 ( .A1(n_295), .A2(n_367), .B1(n_1691), .B2(n_1694), .Y(n_1709) );
AO22x1_ASAP7_75t_L g1713 ( .A1(n_296), .A2(n_302), .B1(n_1684), .B2(n_1698), .Y(n_1713) );
INVx1_ASAP7_75t_L g431 ( .A(n_297), .Y(n_431) );
INVx1_ASAP7_75t_L g449 ( .A(n_297), .Y(n_449) );
INVx1_ASAP7_75t_L g940 ( .A(n_298), .Y(n_940) );
INVx1_ASAP7_75t_L g1011 ( .A(n_300), .Y(n_1011) );
INVxp67_ASAP7_75t_SL g1041 ( .A(n_301), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_303), .Y(n_1072) );
AOI21xp33_ASAP7_75t_L g1117 ( .A1(n_304), .A2(n_714), .B(n_715), .Y(n_1117) );
INVxp67_ASAP7_75t_L g1137 ( .A(n_304), .Y(n_1137) );
INVx1_ASAP7_75t_L g1384 ( .A(n_306), .Y(n_1384) );
INVx1_ASAP7_75t_L g740 ( .A(n_308), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_308), .B(n_747), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g1299 ( .A(n_309), .Y(n_1299) );
INVxp33_ASAP7_75t_L g1190 ( .A(n_311), .Y(n_1190) );
CKINVDCx5p33_ASAP7_75t_R g1606 ( .A(n_312), .Y(n_1606) );
INVx1_ASAP7_75t_L g1196 ( .A(n_313), .Y(n_1196) );
INVx1_ASAP7_75t_L g825 ( .A(n_314), .Y(n_825) );
INVx1_ASAP7_75t_L g617 ( .A(n_315), .Y(n_617) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_316), .B(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1693 ( .A(n_316), .Y(n_1693) );
INVx1_ASAP7_75t_L g1981 ( .A(n_317), .Y(n_1981) );
INVx1_ASAP7_75t_L g1399 ( .A(n_319), .Y(n_1399) );
AOI221xp5_ASAP7_75t_SL g1256 ( .A1(n_320), .A2(n_322), .B1(n_1249), .B2(n_1257), .C(n_1258), .Y(n_1256) );
INVx1_ASAP7_75t_L g1920 ( .A(n_321), .Y(n_1920) );
INVx1_ASAP7_75t_L g1239 ( .A(n_322), .Y(n_1239) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_323), .A2(n_1218), .B1(n_1219), .B2(n_1273), .Y(n_1217) );
INVx1_ASAP7_75t_L g1273 ( .A(n_323), .Y(n_1273) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_324), .A2(n_343), .B1(n_439), .B2(n_444), .C(n_450), .Y(n_1370) );
OAI21xp33_ASAP7_75t_L g1389 ( .A1(n_324), .A2(n_595), .B(n_753), .Y(n_1389) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_325), .A2(n_1544), .B1(n_1586), .B2(n_1587), .Y(n_1543) );
INVx1_ASAP7_75t_L g1587 ( .A(n_325), .Y(n_1587) );
XOR2x2_ASAP7_75t_L g1098 ( .A(n_326), .B(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g990 ( .A(n_327), .Y(n_990) );
INVx1_ASAP7_75t_L g1377 ( .A(n_328), .Y(n_1377) );
INVx1_ASAP7_75t_L g1419 ( .A(n_329), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_329), .A2(n_356), .B1(n_502), .B2(n_1242), .Y(n_1439) );
INVx1_ASAP7_75t_L g1551 ( .A(n_330), .Y(n_1551) );
INVx1_ASAP7_75t_L g915 ( .A(n_331), .Y(n_915) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_332), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_333), .A2(n_343), .B1(n_987), .B2(n_1272), .Y(n_1390) );
INVx1_ASAP7_75t_L g1326 ( .A(n_334), .Y(n_1326) );
INVx1_ASAP7_75t_L g1667 ( .A(n_336), .Y(n_1667) );
INVx1_ASAP7_75t_L g1410 ( .A(n_337), .Y(n_1410) );
INVx1_ASAP7_75t_L g802 ( .A(n_338), .Y(n_802) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_338), .A2(n_753), .B1(n_841), .B2(n_849), .C(n_850), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_340), .A2(n_352), .B1(n_502), .B2(n_1031), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1949 ( .A1(n_341), .A2(n_1950), .B1(n_1951), .B2(n_1992), .Y(n_1949) );
INVxp67_ASAP7_75t_SL g1950 ( .A(n_341), .Y(n_1950) );
INVx1_ASAP7_75t_L g1170 ( .A(n_342), .Y(n_1170) );
INVx1_ASAP7_75t_L g1349 ( .A(n_344), .Y(n_1349) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_345), .Y(n_395) );
INVx1_ASAP7_75t_L g1110 ( .A(n_346), .Y(n_1110) );
XNOR2x1_ASAP7_75t_L g1365 ( .A(n_347), .B(n_1366), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g1283 ( .A(n_348), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1455 ( .A(n_350), .Y(n_1455) );
INVx1_ASAP7_75t_L g1259 ( .A(n_351), .Y(n_1259) );
AOI21xp33_ASAP7_75t_L g1083 ( .A1(n_354), .A2(n_546), .B(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g935 ( .A(n_357), .Y(n_935) );
INVx1_ASAP7_75t_L g1443 ( .A(n_358), .Y(n_1443) );
INVx1_ASAP7_75t_L g1931 ( .A(n_359), .Y(n_1931) );
CKINVDCx5p33_ASAP7_75t_R g1454 ( .A(n_360), .Y(n_1454) );
INVx1_ASAP7_75t_L g783 ( .A(n_361), .Y(n_783) );
INVx1_ASAP7_75t_L g1433 ( .A(n_363), .Y(n_1433) );
XOR2xp5_ASAP7_75t_L g1276 ( .A(n_364), .B(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1548 ( .A(n_365), .Y(n_1548) );
INVx1_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
INVx2_ASAP7_75t_L g509 ( .A(n_366), .Y(n_509) );
INVx1_ASAP7_75t_L g524 ( .A(n_366), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_368), .A2(n_369), .B1(n_546), .B2(n_692), .C(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g1075 ( .A(n_370), .Y(n_1075) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_372), .Y(n_804) );
INVxp67_ASAP7_75t_SL g1132 ( .A(n_373), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g1157 ( .A(n_374), .Y(n_1157) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_400), .B(n_1674), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1943 ( .A(n_379), .B(n_388), .Y(n_1943) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1947 ( .A(n_381), .B(n_384), .Y(n_1947) );
INVx1_ASAP7_75t_L g1996 ( .A(n_381), .Y(n_1996) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1998 ( .A(n_384), .B(n_1996), .Y(n_1998) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g1506 ( .A(n_388), .B(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g586 ( .A(n_389), .B(n_399), .Y(n_586) );
AND2x4_ASAP7_75t_L g695 ( .A(n_389), .B(n_398), .Y(n_695) );
AND2x4_ASAP7_75t_SL g1942 ( .A(n_390), .B(n_1943), .Y(n_1942) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
BUFx4f_ASAP7_75t_L g567 ( .A(n_392), .Y(n_567) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_392), .Y(n_1396) );
INVx1_ASAP7_75t_L g1421 ( .A(n_392), .Y(n_1421) );
OR2x6_ASAP7_75t_L g1485 ( .A(n_392), .B(n_1481), .Y(n_1485) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx4f_ASAP7_75t_L g687 ( .A(n_393), .Y(n_687) );
INVx3_ASAP7_75t_L g976 ( .A(n_393), .Y(n_976) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
AND2x2_ASAP7_75t_L g515 ( .A(n_395), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g528 ( .A(n_395), .Y(n_528) );
INVx1_ASAP7_75t_L g542 ( .A(n_395), .Y(n_542) );
AND2x2_ASAP7_75t_L g548 ( .A(n_395), .B(n_396), .Y(n_548) );
NAND2x1_ASAP7_75t_L g553 ( .A(n_395), .B(n_396), .Y(n_553) );
INVx1_ASAP7_75t_L g421 ( .A(n_396), .Y(n_421) );
INVx2_ASAP7_75t_L g516 ( .A(n_396), .Y(n_516) );
AND2x2_ASAP7_75t_L g527 ( .A(n_396), .B(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g536 ( .A(n_396), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_396), .B(n_528), .Y(n_573) );
OR2x2_ASAP7_75t_L g772 ( .A(n_396), .B(n_420), .Y(n_772) );
OR2x6_ASAP7_75t_L g1900 ( .A(n_397), .B(n_976), .Y(n_1900) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g1497 ( .A(n_398), .Y(n_1497) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g1491 ( .A(n_399), .Y(n_1491) );
AND2x4_ASAP7_75t_L g1503 ( .A(n_399), .B(n_541), .Y(n_1503) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_1361), .B2(n_1673), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_1094), .Y(n_402) );
XNOR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_857), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_699), .B2(n_856), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OA22x2_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_598), .B2(n_599), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AO211x2_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_422), .C(n_517), .Y(n_409) );
INVx3_ASAP7_75t_L g747 ( .A(n_411), .Y(n_747) );
AOI222xp33_ASAP7_75t_L g788 ( .A1(n_411), .A2(n_512), .B1(n_789), .B2(n_790), .C1(n_793), .C2(n_794), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_411), .A2(n_512), .B1(n_990), .B2(n_991), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_411), .B(n_998), .Y(n_997) );
AOI211xp5_ASAP7_75t_L g1071 ( .A1(n_411), .A2(n_1072), .B(n_1073), .C(n_1077), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_411), .B(n_1403), .Y(n_1402) );
AOI211x1_ASAP7_75t_L g1405 ( .A1(n_411), .A2(n_1406), .B(n_1407), .C(n_1427), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_411), .A2(n_1265), .B1(n_1548), .B2(n_1567), .Y(n_1585) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
AND2x4_ASAP7_75t_L g512 ( .A(n_412), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g539 ( .A(n_413), .B(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_L g650 ( .A(n_413), .Y(n_650) );
OR2x2_ASAP7_75t_L g987 ( .A(n_413), .B(n_540), .Y(n_987) );
INVx1_ASAP7_75t_L g1507 ( .A(n_413), .Y(n_1507) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g585 ( .A(n_414), .Y(n_585) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g671 ( .A(n_416), .Y(n_671) );
BUFx6f_ASAP7_75t_L g1298 ( .A(n_416), .Y(n_1298) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_L g513 ( .A(n_417), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_417), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g655 ( .A(n_417), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g674 ( .A(n_417), .B(n_514), .Y(n_674) );
AND2x4_ASAP7_75t_SL g679 ( .A(n_417), .B(n_547), .Y(n_679) );
BUFx2_ASAP7_75t_L g872 ( .A(n_417), .Y(n_872) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_417), .B(n_525), .Y(n_1596) );
HB1xp67_ASAP7_75t_L g1481 ( .A(n_418), .Y(n_1481) );
INVx3_ASAP7_75t_L g581 ( .A(n_419), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_419), .B(n_533), .Y(n_592) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_419), .Y(n_778) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_466), .B(n_506), .C(n_510), .Y(n_422) );
AOI211xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_437), .B(n_438), .C(n_455), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_424), .A2(n_730), .B1(n_733), .B2(n_743), .Y(n_729) );
INVx2_ASAP7_75t_L g1038 ( .A(n_424), .Y(n_1038) );
AOI211xp5_ASAP7_75t_SL g1047 ( .A1(n_424), .A2(n_1048), .B(n_1049), .C(n_1050), .Y(n_1047) );
AOI211xp5_ASAP7_75t_L g1101 ( .A1(n_424), .A2(n_1102), .B(n_1103), .C(n_1104), .Y(n_1101) );
AOI211xp5_ASAP7_75t_L g1319 ( .A1(n_424), .A2(n_1320), .B(n_1321), .C(n_1322), .Y(n_1319) );
AOI211xp5_ASAP7_75t_L g1368 ( .A1(n_424), .A2(n_1369), .B(n_1370), .C(n_1371), .Y(n_1368) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x6_ASAP7_75t_L g649 ( .A(n_425), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g791 ( .A(n_425), .B(n_650), .Y(n_791) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_426), .B(n_432), .Y(n_425) );
INVx8_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
AND2x2_ASAP7_75t_L g488 ( .A(n_426), .B(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g708 ( .A(n_426), .Y(n_708) );
BUFx3_ASAP7_75t_L g723 ( .A(n_426), .Y(n_723) );
HB1xp67_ASAP7_75t_L g1646 ( .A(n_426), .Y(n_1646) );
AND2x4_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
AND2x4_ASAP7_75t_L g461 ( .A(n_427), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_428), .Y(n_443) );
AND2x4_ASAP7_75t_L g492 ( .A(n_428), .B(n_448), .Y(n_492) );
OR2x2_ASAP7_75t_L g498 ( .A(n_428), .B(n_430), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_428), .B(n_449), .Y(n_645) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
AND2x6_ASAP7_75t_L g440 ( .A(n_432), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g445 ( .A(n_432), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g454 ( .A(n_432), .Y(n_454) );
AND2x4_ASAP7_75t_L g606 ( .A(n_432), .B(n_590), .Y(n_606) );
AND2x4_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_433), .B(n_505), .Y(n_504) );
NAND3x1_ASAP7_75t_L g635 ( .A(n_433), .B(n_505), .C(n_636), .Y(n_635) );
OR2x4_ASAP7_75t_L g1512 ( .A(n_433), .B(n_498), .Y(n_1512) );
INVx1_ASAP7_75t_L g1515 ( .A(n_433), .Y(n_1515) );
AND2x4_ASAP7_75t_L g1520 ( .A(n_433), .B(n_492), .Y(n_1520) );
OR2x6_ASAP7_75t_L g1535 ( .A(n_433), .B(n_738), .Y(n_1535) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
NAND2xp33_ASAP7_75t_SL g716 ( .A(n_434), .B(n_436), .Y(n_716) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g482 ( .A(n_436), .B(n_483), .Y(n_482) );
AND3x4_ASAP7_75t_L g622 ( .A(n_436), .B(n_483), .C(n_508), .Y(n_622) );
HB1xp67_ASAP7_75t_L g1538 ( .A(n_436), .Y(n_1538) );
AOI222xp33_ASAP7_75t_L g518 ( .A1(n_437), .A2(n_519), .B1(n_529), .B2(n_537), .C1(n_538), .C2(n_543), .Y(n_518) );
INVx4_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_440), .A2(n_445), .B1(n_726), .B2(n_727), .C(n_728), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_440), .A2(n_445), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_440), .A2(n_445), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_440), .A2(n_445), .B1(n_1410), .B2(n_1424), .Y(n_1442) );
AOI221xp5_ASAP7_75t_L g1550 ( .A1(n_440), .A2(n_445), .B1(n_728), .B2(n_1551), .C(n_1552), .Y(n_1550) );
AND2x2_ASAP7_75t_L g605 ( .A(n_441), .B(n_606), .Y(n_605) );
NAND2x1_ASAP7_75t_L g1212 ( .A(n_441), .B(n_606), .Y(n_1212) );
AND2x4_ASAP7_75t_SL g1626 ( .A(n_441), .B(n_606), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_441), .B(n_606), .Y(n_1655) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_443), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g465 ( .A(n_443), .B(n_447), .Y(n_465) );
BUFx2_ASAP7_75t_L g1525 ( .A(n_443), .Y(n_1525) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_445), .Y(n_1024) );
INVx1_ASAP7_75t_L g610 ( .A(n_446), .Y(n_610) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g453 ( .A(n_449), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_450), .Y(n_728) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
INVx1_ASAP7_75t_L g1064 ( .A(n_451), .Y(n_1064) );
INVx1_ASAP7_75t_L g1518 ( .A(n_451), .Y(n_1518) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
BUFx3_ASAP7_75t_L g814 ( .A(n_452), .Y(n_814) );
BUFx2_ASAP7_75t_L g1528 ( .A(n_453), .Y(n_1528) );
INVx1_ASAP7_75t_L g943 ( .A(n_454), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_456), .Y(n_1120) );
OR2x6_ASAP7_75t_SL g456 ( .A(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g464 ( .A(n_458), .B(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_458), .Y(n_732) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g489 ( .A(n_459), .Y(n_489) );
OR2x2_ASAP7_75t_L g616 ( .A(n_459), .B(n_585), .Y(n_616) );
INVx3_ASAP7_75t_L g900 ( .A(n_460), .Y(n_900) );
INVx1_ASAP7_75t_L g1185 ( .A(n_460), .Y(n_1185) );
BUFx2_ASAP7_75t_L g1937 ( .A(n_460), .Y(n_1937) );
BUFx2_ASAP7_75t_L g1986 ( .A(n_460), .Y(n_1986) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_461), .Y(n_472) );
BUFx8_ASAP7_75t_L g619 ( .A(n_461), .Y(n_619) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_461), .Y(n_714) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_464), .B(n_745), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_464), .A2(n_1120), .B1(n_1121), .B2(n_1122), .C(n_1123), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1547 ( .A1(n_464), .A2(n_1120), .B1(n_1548), .B2(n_1549), .Y(n_1547) );
BUFx3_ASAP7_75t_L g485 ( .A(n_465), .Y(n_485) );
BUFx12f_ASAP7_75t_L g502 ( .A(n_465), .Y(n_502) );
INVx5_ASAP7_75t_L g629 ( .A(n_465), .Y(n_629) );
BUFx2_ASAP7_75t_L g709 ( .A(n_465), .Y(n_709) );
BUFx3_ASAP7_75t_L g934 ( .A(n_465), .Y(n_934) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_486), .C(n_493), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_473), .C(n_484), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_469), .B(n_550), .Y(n_561) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g1194 ( .A(n_471), .Y(n_1194) );
INVx1_ASAP7_75t_L g1238 ( .A(n_471), .Y(n_1238) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g967 ( .A(n_472), .Y(n_967) );
INVx2_ASAP7_75t_L g1035 ( .A(n_472), .Y(n_1035) );
INVx1_ASAP7_75t_L g1054 ( .A(n_472), .Y(n_1054) );
INVx2_ASAP7_75t_L g1236 ( .A(n_472), .Y(n_1236) );
AND2x4_ASAP7_75t_L g1514 ( .A(n_472), .B(n_1515), .Y(n_1514) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_476), .A2(n_955), .B1(n_1461), .B2(n_1462), .Y(n_1460) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g648 ( .A(n_477), .B(n_616), .Y(n_648) );
INVx3_ASAP7_75t_L g807 ( .A(n_477), .Y(n_807) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_477), .Y(n_913) );
INVx4_ASAP7_75t_L g954 ( .A(n_477), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_479), .A2(n_711), .B1(n_793), .B2(n_799), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g905 ( .A1(n_479), .A2(n_606), .B(n_870), .C(n_906), .Y(n_905) );
INVx8_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g614 ( .A(n_480), .Y(n_614) );
INVx2_ASAP7_75t_L g624 ( .A(n_480), .Y(n_624) );
INVx3_ASAP7_75t_L g941 ( .A(n_480), .Y(n_941) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_482), .A2(n_964), .B1(n_965), .B2(n_966), .C(n_968), .Y(n_963) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_482), .A2(n_629), .B1(n_707), .B2(n_1058), .C(n_1059), .Y(n_1057) );
OAI21xp33_ASAP7_75t_L g1325 ( .A1(n_482), .A2(n_1032), .B(n_1326), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g1376 ( .A1(n_482), .A2(n_821), .B1(n_1116), .B2(n_1377), .C(n_1378), .Y(n_1376) );
INVx3_ASAP7_75t_L g1524 ( .A(n_483), .Y(n_1524) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_488), .A2(n_491), .B1(n_1244), .B2(n_1245), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_488), .A2(n_491), .B1(n_1406), .B2(n_1411), .Y(n_1440) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_488), .A2(n_491), .B1(n_1567), .B2(n_1568), .Y(n_1566) );
AND2x2_ASAP7_75t_L g491 ( .A(n_489), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g626 ( .A(n_492), .Y(n_626) );
BUFx2_ASAP7_75t_L g639 ( .A(n_492), .Y(n_639) );
BUFx2_ASAP7_75t_L g711 ( .A(n_492), .Y(n_711) );
BUFx3_ASAP7_75t_L g721 ( .A(n_492), .Y(n_721) );
BUFx2_ASAP7_75t_L g742 ( .A(n_492), .Y(n_742) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_492), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1559 ( .A(n_492), .Y(n_1559) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI221xp5_ASAP7_75t_L g1333 ( .A1(n_497), .A2(n_503), .B1(n_814), .B2(n_1334), .C(n_1335), .Y(n_1333) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx4f_ASAP7_75t_L g818 ( .A(n_498), .Y(n_818) );
BUFx3_ASAP7_75t_L g955 ( .A(n_498), .Y(n_955) );
INVx2_ASAP7_75t_L g961 ( .A(n_498), .Y(n_961) );
OR2x4_ASAP7_75t_L g1532 ( .A(n_498), .B(n_1515), .Y(n_1532) );
INVx1_ASAP7_75t_L g1437 ( .A(n_499), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
BUFx2_ASAP7_75t_L g1375 ( .A(n_502), .Y(n_1375) );
INVx3_ASAP7_75t_L g724 ( .A(n_503), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g811 ( .A1(n_503), .A2(n_812), .B1(n_815), .B2(n_816), .C(n_819), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_503), .A2(n_952), .B1(n_953), .B2(n_955), .C(n_956), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_503), .B(n_1066), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1382 ( .A1(n_503), .A2(n_955), .B1(n_1116), .B2(n_1383), .C(n_1384), .Y(n_1382) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g926 ( .A(n_504), .B(n_558), .Y(n_926) );
OR2x6_ASAP7_75t_L g1652 ( .A(n_504), .B(n_558), .Y(n_1652) );
OAI21xp33_ASAP7_75t_L g1593 ( .A1(n_506), .A2(n_1594), .B(n_1603), .Y(n_1593) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g698 ( .A(n_507), .Y(n_698) );
BUFx2_ASAP7_75t_L g1973 ( .A(n_507), .Y(n_1973) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_508), .A2(n_1020), .B1(n_1039), .B2(n_1041), .Y(n_1019) );
INVx2_ASAP7_75t_SL g1067 ( .A(n_508), .Y(n_1067) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_509), .B(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g558 ( .A(n_509), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_512), .Y(n_756) );
INVx1_ASAP7_75t_L g1040 ( .A(n_512), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_512), .B(n_1069), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_512), .B(n_1121), .Y(n_1150) );
INVx1_ASAP7_75t_L g1266 ( .A(n_512), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_512), .B(n_1343), .Y(n_1342) );
INVx2_ASAP7_75t_L g564 ( .A(n_514), .Y(n_564) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_514), .Y(n_693) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx3_ASAP7_75t_L g577 ( .A(n_515), .Y(n_577) );
INVx2_ASAP7_75t_L g760 ( .A(n_515), .Y(n_760) );
AND2x4_ASAP7_75t_L g1480 ( .A(n_515), .B(n_1481), .Y(n_1480) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_544), .C(n_587), .Y(n_517) );
INVxp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_L g752 ( .A(n_521), .Y(n_752) );
INVx1_ASAP7_75t_L g792 ( .A(n_521), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_521), .A2(n_1002), .B1(n_1003), .B2(n_1004), .Y(n_1001) );
AOI222xp33_ASAP7_75t_L g1148 ( .A1(n_521), .A2(n_588), .B1(n_1004), .B2(n_1102), .C1(n_1122), .C2(n_1149), .Y(n_1148) );
AOI211xp5_ASAP7_75t_L g1268 ( .A1(n_521), .A2(n_1269), .B(n_1270), .C(n_1271), .Y(n_1268) );
AOI222xp33_ASAP7_75t_L g1339 ( .A1(n_521), .A2(n_588), .B1(n_1004), .B2(n_1320), .C1(n_1340), .C2(n_1341), .Y(n_1339) );
AOI211xp5_ASAP7_75t_L g1388 ( .A1(n_521), .A2(n_1369), .B(n_1389), .C(n_1390), .Y(n_1388) );
AOI222xp33_ASAP7_75t_L g1408 ( .A1(n_521), .A2(n_529), .B1(n_538), .B2(n_1409), .C1(n_1410), .C2(n_1411), .Y(n_1408) );
AOI222xp33_ASAP7_75t_L g1569 ( .A1(n_521), .A2(n_588), .B1(n_1004), .B2(n_1549), .C1(n_1552), .C2(n_1570), .Y(n_1569) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g551 ( .A(n_523), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g753 ( .A(n_523), .B(n_552), .Y(n_753) );
INVx1_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
INVx1_ASAP7_75t_L g636 ( .A(n_524), .Y(n_636) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g1611 ( .A(n_526), .Y(n_1611) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g579 ( .A(n_527), .Y(n_579) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_527), .Y(n_656) );
BUFx3_ASAP7_75t_L g779 ( .A(n_527), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_529), .A2(n_538), .B1(n_799), .B2(n_801), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g1009 ( .A1(n_529), .A2(n_538), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_529), .A2(n_538), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_SL g986 ( .A(n_530), .Y(n_986) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_530), .Y(n_1272) );
NAND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_533), .B(n_541), .Y(n_540) );
AND2x6_ASAP7_75t_L g668 ( .A(n_533), .B(n_547), .Y(n_668) );
INVx1_ASAP7_75t_L g683 ( .A(n_533), .Y(n_683) );
AND2x2_ASAP7_75t_L g878 ( .A(n_533), .B(n_879), .Y(n_878) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g682 ( .A(n_536), .Y(n_682) );
BUFx2_ASAP7_75t_L g879 ( .A(n_536), .Y(n_879) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_536), .B(n_1491), .Y(n_1499) );
AND2x4_ASAP7_75t_L g1893 ( .A(n_536), .B(n_1491), .Y(n_1893) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g647 ( .A(n_539), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g1632 ( .A(n_539), .B(n_648), .Y(n_1632) );
INVx1_ASAP7_75t_L g881 ( .A(n_540), .Y(n_881) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_560), .B1(n_574), .B2(n_578), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_546), .A2(n_579), .B1(n_870), .B2(n_871), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_546), .A2(n_847), .B(n_875), .C(n_876), .Y(n_874) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g575 ( .A(n_547), .Y(n_575) );
BUFx3_ASAP7_75t_L g761 ( .A(n_547), .Y(n_761) );
BUFx6f_ASAP7_75t_L g1088 ( .A(n_547), .Y(n_1088) );
BUFx3_ASAP7_75t_L g1308 ( .A(n_547), .Y(n_1308) );
INVx1_ASAP7_75t_L g1417 ( .A(n_547), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_547), .B(n_1497), .Y(n_1496) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g663 ( .A(n_548), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_549), .A2(n_561), .B1(n_562), .B2(n_565), .Y(n_560) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g1004 ( .A(n_551), .Y(n_1004) );
BUFx3_ASAP7_75t_L g977 ( .A(n_552), .Y(n_977) );
INVx2_ASAP7_75t_SL g1472 ( .A(n_552), .Y(n_1472) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_553), .Y(n_596) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_SL g831 ( .A(n_556), .Y(n_831) );
INVx4_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g781 ( .A(n_557), .Y(n_781) );
HB1xp67_ASAP7_75t_L g972 ( .A(n_557), .Y(n_972) );
AOI31xp33_ASAP7_75t_L g1006 ( .A1(n_557), .A2(n_594), .A3(n_1007), .B(n_1008), .Y(n_1006) );
INVx2_ASAP7_75t_L g1084 ( .A(n_557), .Y(n_1084) );
INVx2_ASAP7_75t_L g1130 ( .A(n_557), .Y(n_1130) );
INVx1_ASAP7_75t_L g1464 ( .A(n_557), .Y(n_1464) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g745 ( .A(n_558), .Y(n_745) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g665 ( .A(n_563), .Y(n_665) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g1162 ( .A(n_564), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_567), .A2(n_569), .B1(n_1059), .B2(n_1082), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_567), .A2(n_1135), .B1(n_1399), .B2(n_1400), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1930 ( .A1(n_567), .A2(n_569), .B1(n_1931), .B2(n_1932), .Y(n_1930) );
INVx5_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx6_ASAP7_75t_L g689 ( .A(n_570), .Y(n_689) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g1092 ( .A(n_571), .Y(n_1092) );
INVx2_ASAP7_75t_SL g1261 ( .A(n_571), .Y(n_1261) );
INVx4_ASAP7_75t_L g1423 ( .A(n_571), .Y(n_1423) );
INVx1_ASAP7_75t_L g1476 ( .A(n_571), .Y(n_1476) );
INVx1_ASAP7_75t_L g1970 ( .A(n_571), .Y(n_1970) );
INVx8_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_572), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1490 ( .A(n_572), .B(n_1491), .Y(n_1490) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g1576 ( .A(n_577), .Y(n_1576) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_579), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_579), .Y(n_1176) );
INVx1_ASAP7_75t_SL g1254 ( .A(n_579), .Y(n_1254) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g838 ( .A(n_581), .Y(n_838) );
INVx2_ASAP7_75t_L g983 ( .A(n_581), .Y(n_983) );
INVx1_ASAP7_75t_L g1252 ( .A(n_581), .Y(n_1252) );
INVx1_ASAP7_75t_L g1610 ( .A(n_581), .Y(n_1610) );
INVx1_ASAP7_75t_L g1578 ( .A(n_582), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
AND2x4_ASAP7_75t_L g766 ( .A(n_583), .B(n_586), .Y(n_766) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g909 ( .A(n_585), .B(n_716), .Y(n_909) );
AND2x2_ASAP7_75t_SL g1146 ( .A(n_585), .B(n_586), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1540 ( .A(n_585), .Y(n_1540) );
INVx4_ASAP7_75t_L g666 ( .A(n_586), .Y(n_666) );
INVx4_ASAP7_75t_L g891 ( .A(n_586), .Y(n_891) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_593), .B(n_594), .Y(n_587) );
AOI322xp5_ASAP7_75t_L g1078 ( .A1(n_588), .A2(n_766), .A3(n_1079), .B1(n_1080), .B2(n_1083), .C1(n_1085), .C2(n_1086), .Y(n_1078) );
AOI322xp5_ASAP7_75t_L g1247 ( .A1(n_588), .A2(n_766), .A3(n_1248), .B1(n_1251), .B2(n_1255), .C1(n_1256), .C2(n_1262), .Y(n_1247) );
AOI222xp33_ASAP7_75t_L g1391 ( .A1(n_588), .A2(n_766), .B1(n_972), .B2(n_1392), .C1(n_1397), .C2(n_1401), .Y(n_1391) );
AOI21xp33_ASAP7_75t_L g1425 ( .A1(n_588), .A2(n_594), .B(n_1426), .Y(n_1425) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g646 ( .A(n_590), .B(n_592), .Y(n_646) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR3x1_ASAP7_75t_L g1344 ( .A(n_594), .B(n_1345), .C(n_1346), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_595), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_595), .A2(n_768), .B(n_780), .Y(n_767) );
OAI21xp5_ASAP7_75t_SL g828 ( .A1(n_595), .A2(n_829), .B(n_832), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g978 ( .A1(n_595), .A2(n_849), .B(n_979), .Y(n_978) );
OAI21xp5_ASAP7_75t_L g1580 ( .A1(n_595), .A2(n_1581), .B(n_1582), .Y(n_1580) );
OR2x6_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx4_ASAP7_75t_L g775 ( .A(n_596), .Y(n_775) );
BUFx4f_ASAP7_75t_L g836 ( .A(n_596), .Y(n_836) );
BUFx4f_ASAP7_75t_L g845 ( .A(n_596), .Y(n_845) );
BUFx6f_ASAP7_75t_L g1140 ( .A(n_596), .Y(n_1140) );
BUFx4f_ASAP7_75t_L g1348 ( .A(n_596), .Y(n_1348) );
BUFx4f_ASAP7_75t_L g1607 ( .A(n_596), .Y(n_1607) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_652), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_640), .C(n_651), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_611), .C(n_620), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_607), .B2(n_608), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g1979 ( .A1(n_605), .A2(n_608), .B1(n_1980), .B2(n_1981), .Y(n_1979) );
AND2x4_ASAP7_75t_L g608 ( .A(n_606), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g651 ( .A(n_606), .B(n_639), .Y(n_651) );
AND2x4_ASAP7_75t_SL g1628 ( .A(n_606), .B(n_609), .Y(n_1628) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_608), .A2(n_1166), .B1(n_1170), .B2(n_1211), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_608), .A2(n_1211), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1653 ( .A1(n_608), .A2(n_1654), .B1(n_1655), .B2(n_1656), .Y(n_1653) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_617), .B2(n_618), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_612), .A2(n_617), .B1(n_670), .B2(n_672), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_613), .B(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_613), .A2(n_618), .B1(n_1297), .B2(n_1299), .Y(n_1315) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x4_ASAP7_75t_L g1634 ( .A(n_614), .B(n_615), .Y(n_1634) );
AND2x4_ASAP7_75t_L g618 ( .A(n_615), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g642 ( .A(n_616), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g901 ( .A(n_616), .Y(n_901) );
INVx2_ASAP7_75t_L g1201 ( .A(n_618), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1633 ( .A1(n_618), .A2(n_1598), .B1(n_1599), .B2(n_1634), .Y(n_1633) );
INVx2_ASAP7_75t_L g1990 ( .A(n_618), .Y(n_1990) );
INVx3_ASAP7_75t_L g632 ( .A(n_619), .Y(n_632) );
INVx2_ASAP7_75t_SL g821 ( .A(n_619), .Y(n_821) );
INVx3_ASAP7_75t_L g1032 ( .A(n_619), .Y(n_1032) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_619), .Y(n_1109) );
AOI33xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .A3(n_627), .B1(n_630), .B2(n_634), .B3(n_637), .Y(n_620) );
AOI33xp33_ASAP7_75t_L g1285 ( .A1(n_621), .A2(n_1286), .A3(n_1290), .B1(n_1291), .B2(n_1292), .B3(n_1293), .Y(n_1285) );
AOI33xp33_ASAP7_75t_L g1982 ( .A1(n_621), .A2(n_634), .A3(n_1983), .B1(n_1984), .B2(n_1987), .B3(n_1988), .Y(n_1982) );
BUFx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI33xp33_ASAP7_75t_L g1644 ( .A1(n_622), .A2(n_1645), .A3(n_1648), .B1(n_1649), .B2(n_1650), .B3(n_1651), .Y(n_1644) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_624), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g936 ( .A(n_626), .Y(n_936) );
INVx2_ASAP7_75t_L g1647 ( .A(n_626), .Y(n_1647) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g633 ( .A(n_629), .Y(n_633) );
INVx2_ASAP7_75t_R g1381 ( .A(n_629), .Y(n_1381) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g1459 ( .A(n_634), .Y(n_1459) );
CKINVDCx5p33_ASAP7_75t_R g1623 ( .A(n_634), .Y(n_1623) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g1200 ( .A(n_635), .Y(n_1200) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_639), .A2(n_941), .B1(n_998), .B2(n_1011), .Y(n_1036) );
INVx8_ASAP7_75t_L g1204 ( .A(n_641), .Y(n_1204) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_646), .Y(n_641) );
INVx1_ASAP7_75t_L g1112 ( .A(n_643), .Y(n_1112) );
BUFx3_ASAP7_75t_L g1187 ( .A(n_643), .Y(n_1187) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_644), .Y(n_824) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g738 ( .A(n_645), .Y(n_738) );
INVx1_ASAP7_75t_L g751 ( .A(n_646), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_646), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g1156 ( .A(n_647), .Y(n_1156) );
INVx2_ASAP7_75t_L g902 ( .A(n_648), .Y(n_902) );
INVx3_ASAP7_75t_L g1203 ( .A(n_649), .Y(n_1203) );
INVx3_ASAP7_75t_L g1213 ( .A(n_651), .Y(n_1213) );
NOR3xp33_ASAP7_75t_L g1612 ( .A(n_651), .B(n_1613), .C(n_1624), .Y(n_1612) );
INVx3_ASAP7_75t_L g1643 ( .A(n_651), .Y(n_1643) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_675), .B(n_696), .Y(n_652) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g1177 ( .A1(n_655), .A2(n_1178), .B1(n_1179), .B2(n_1180), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_655), .A2(n_668), .B1(n_1279), .B2(n_1301), .C(n_1305), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1662 ( .A1(n_655), .A2(n_668), .B1(n_1640), .B2(n_1663), .C(n_1664), .Y(n_1662) );
BUFx2_ASAP7_75t_L g839 ( .A(n_656), .Y(n_839) );
INVx1_ASAP7_75t_L g1015 ( .A(n_656), .Y(n_1015) );
AOI21xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_667), .B(n_668), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g1018 ( .A(n_662), .Y(n_1018) );
INVx1_ASAP7_75t_L g1577 ( .A(n_662), .Y(n_1577) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g1304 ( .A(n_663), .Y(n_1304) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_SL g1174 ( .A(n_666), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_668), .A2(n_1169), .B1(n_1170), .B2(n_1171), .C(n_1175), .Y(n_1168) );
AOI21xp5_ASAP7_75t_L g1600 ( .A1(n_668), .A2(n_1601), .B(n_1602), .Y(n_1600) );
AOI21xp5_ASAP7_75t_L g1957 ( .A1(n_668), .A2(n_1958), .B(n_1959), .Y(n_1957) );
AOI222xp33_ASAP7_75t_L g1159 ( .A1(n_670), .A2(n_878), .B1(n_1160), .B2(n_1164), .C1(n_1166), .C2(n_1167), .Y(n_1159) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g1961 ( .A1(n_672), .A2(n_1962), .B1(n_1963), .B2(n_1964), .Y(n_1961) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx6f_ASAP7_75t_L g1178 ( .A(n_674), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_674), .A2(n_1298), .B1(n_1598), .B2(n_1599), .Y(n_1597) );
AOI22xp33_ASAP7_75t_L g1666 ( .A1(n_674), .A2(n_1298), .B1(n_1667), .B2(n_1668), .Y(n_1666) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g1604 ( .A(n_677), .Y(n_1604) );
INVx2_ASAP7_75t_L g1966 ( .A(n_677), .Y(n_1966) );
INVx4_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx3_ASAP7_75t_L g1169 ( .A(n_679), .Y(n_1169) );
BUFx2_ASAP7_75t_L g1967 ( .A(n_680), .Y(n_1967) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g876 ( .A(n_683), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B1(n_689), .B2(n_690), .C(n_691), .Y(n_684) );
OAI22xp5_ASAP7_75t_SL g1258 ( .A1(n_685), .A2(n_1231), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1968 ( .A1(n_685), .A2(n_1969), .B1(n_1970), .B2(n_1971), .C(n_1972), .Y(n_1968) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g1351 ( .A(n_686), .Y(n_1351) );
INVx2_ASAP7_75t_L g1466 ( .A(n_686), .Y(n_1466) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g764 ( .A(n_687), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_689), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g979 ( .A1(n_689), .A2(n_949), .B1(n_964), .B2(n_980), .C(n_982), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_689), .A2(n_1451), .B1(n_1461), .B2(n_1466), .Y(n_1465) );
BUFx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g888 ( .A(n_695), .Y(n_888) );
INVx2_ASAP7_75t_L g1163 ( .A(n_695), .Y(n_1163) );
INVx1_ASAP7_75t_L g1309 ( .A(n_695), .Y(n_1309) );
AOI221xp5_ASAP7_75t_L g1155 ( .A1(n_696), .A2(n_1156), .B1(n_1157), .B2(n_1158), .C(n_1181), .Y(n_1155) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g826 ( .A(n_698), .Y(n_826) );
A2O1A1Ixp33_ASAP7_75t_SL g1100 ( .A1(n_698), .A2(n_1101), .B(n_1119), .C(n_1124), .Y(n_1100) );
INVx2_ASAP7_75t_SL g856 ( .A(n_699), .Y(n_856) );
XNOR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_785), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_783), .B(n_784), .Y(n_700) );
AND3x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_748), .C(n_757), .Y(n_701) );
AOI31xp33_ASAP7_75t_L g784 ( .A1(n_702), .A2(n_748), .A3(n_757), .B(n_783), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_744), .B(n_746), .Y(n_702) );
NAND3xp33_ASAP7_75t_SL g703 ( .A(n_704), .B(n_725), .C(n_729), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_710), .B1(n_717), .B2(n_720), .Y(n_704) );
BUFx2_ASAP7_75t_SL g1374 ( .A(n_706), .Y(n_1374) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
BUFx3_ASAP7_75t_L g1242 ( .A(n_708), .Y(n_1242) );
INVx1_ASAP7_75t_L g1288 ( .A(n_708), .Y(n_1288) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g719 ( .A(n_714), .Y(n_719) );
INVx3_ASAP7_75t_L g734 ( .A(n_714), .Y(n_734) );
INVx5_ASAP7_75t_L g916 ( .A(n_714), .Y(n_916) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_714), .Y(n_948) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1561 ( .A(n_723), .Y(n_1561) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_728), .B(n_1022), .Y(n_1021) );
INVxp67_ASAP7_75t_L g797 ( .A(n_730), .Y(n_797) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g932 ( .A(n_732), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_735), .A2(n_958), .B1(n_959), .B2(n_962), .Y(n_957) );
OAI21xp33_ASAP7_75t_L g1617 ( .A1(n_735), .A2(n_1618), .B(n_1619), .Y(n_1617) );
INVx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g917 ( .A(n_737), .Y(n_917) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
BUFx3_ASAP7_75t_L g950 ( .A(n_738), .Y(n_950) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_742), .Y(n_1234) );
OAI31xp33_ASAP7_75t_SL g1221 ( .A1(n_744), .A2(n_1222), .A3(n_1223), .B(n_1227), .Y(n_1221) );
INVx1_ASAP7_75t_L g1313 ( .A(n_744), .Y(n_1313) );
INVx2_ASAP7_75t_L g1337 ( .A(n_744), .Y(n_1337) );
OAI21xp5_ASAP7_75t_L g1545 ( .A1(n_744), .A2(n_1546), .B(n_1553), .Y(n_1545) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_SL g865 ( .A1(n_745), .A2(n_866), .B(n_883), .Y(n_865) );
INVx1_ASAP7_75t_L g970 ( .A(n_745), .Y(n_970) );
INVx1_ASAP7_75t_L g1126 ( .A(n_747), .Y(n_1126) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_754), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
AOI211xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_766), .B(n_767), .C(n_782), .Y(n_757) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g887 ( .A(n_760), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_766), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g1012 ( .A(n_766), .B(n_1013), .C(n_1016), .Y(n_1012) );
AOI322xp5_ASAP7_75t_L g1412 ( .A1(n_766), .A2(n_1004), .A3(n_1262), .B1(n_1413), .B2(n_1414), .C1(n_1415), .C2(n_1424), .Y(n_1412) );
INVx2_ASAP7_75t_L g1473 ( .A(n_766), .Y(n_1473) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_773), .B1(n_774), .B2(n_776), .C(n_777), .Y(n_768) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g834 ( .A(n_772), .Y(n_834) );
BUFx2_ASAP7_75t_L g844 ( .A(n_772), .Y(n_844) );
INVx1_ASAP7_75t_L g981 ( .A(n_772), .Y(n_981) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_772), .Y(n_1139) );
OAI221xp5_ASAP7_75t_L g1582 ( .A1(n_774), .A2(n_842), .B1(n_1555), .B2(n_1583), .C(n_1584), .Y(n_1582) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g1356 ( .A(n_775), .Y(n_1356) );
INVx2_ASAP7_75t_L g1928 ( .A(n_775), .Y(n_1928) );
INVx3_ASAP7_75t_L g848 ( .A(n_778), .Y(n_848) );
BUFx6f_ASAP7_75t_L g893 ( .A(n_778), .Y(n_893) );
INVx1_ASAP7_75t_L g1262 ( .A(n_780), .Y(n_1262) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_795), .C(n_827), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
OAI21xp33_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_810), .B(n_826), .Y(n_795) );
OAI211xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B(n_800), .C(n_803), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_805), .B(n_808), .C(n_809), .Y(n_803) );
OAI221xp5_ASAP7_75t_L g841 ( .A1(n_804), .A2(n_815), .B1(n_842), .B2(n_845), .C(n_846), .Y(n_841) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI211xp5_ASAP7_75t_L g1562 ( .A1(n_806), .A2(n_1563), .B(n_1564), .C(n_1565), .Y(n_1562) );
OAI22xp33_ASAP7_75t_L g1935 ( .A1(n_806), .A2(n_960), .B1(n_1920), .B2(n_1927), .Y(n_1935) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx3_ASAP7_75t_L g1116 ( .A(n_807), .Y(n_1116) );
INVx2_ASAP7_75t_L g1192 ( .A(n_807), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g1450 ( .A1(n_812), .A2(n_955), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_814), .A2(n_818), .B1(n_924), .B2(n_925), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g1940 ( .A1(n_814), .A2(n_960), .B1(n_1921), .B2(n_1929), .Y(n_1940) );
OAI22xp33_ASAP7_75t_L g1189 ( .A1(n_816), .A2(n_1190), .B1(n_1191), .B2(n_1192), .Y(n_1189) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_818), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_825), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g1938 ( .A1(n_821), .A2(n_1924), .B1(n_1932), .B2(n_1939), .Y(n_1938) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_822), .A2(n_833), .B1(n_835), .B2(n_836), .C(n_837), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g1431 ( .A1(n_823), .A2(n_1422), .B1(n_1432), .B2(n_1433), .C(n_1434), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g1453 ( .A1(n_823), .A2(n_1194), .B1(n_1454), .B2(n_1455), .Y(n_1453) );
OAI221xp5_ASAP7_75t_L g1620 ( .A1(n_823), .A2(n_966), .B1(n_1606), .B2(n_1621), .C(n_1622), .Y(n_1620) );
CKINVDCx8_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g1329 ( .A(n_824), .Y(n_1329) );
INVx3_ASAP7_75t_L g1556 ( .A(n_824), .Y(n_1556) );
INVx3_ASAP7_75t_L g1939 ( .A(n_824), .Y(n_1939) );
INVx1_ASAP7_75t_L g1669 ( .A(n_826), .Y(n_1669) );
NOR3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_840), .C(n_851), .Y(n_827) );
INVxp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g1467 ( .A1(n_833), .A2(n_836), .B1(n_1454), .B2(n_1457), .Y(n_1467) );
INVx1_ASAP7_75t_L g1470 ( .A(n_833), .Y(n_1470) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx2_ASAP7_75t_L g1354 ( .A(n_834), .Y(n_1354) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g868 ( .A(n_843), .Y(n_868) );
INVx4_ASAP7_75t_L g1926 ( .A(n_843), .Y(n_1926) );
INVx4_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g1665 ( .A(n_848), .Y(n_1665) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
XNOR2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_992), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
XNOR2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_927), .Y(n_860) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_894), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_872), .B(n_873), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_868), .A2(n_1326), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_877), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_878), .A2(n_880), .B1(n_881), .B2(n_882), .Y(n_877) );
INVx1_ASAP7_75t_L g1312 ( .A(n_878), .Y(n_1312) );
AOI222xp33_ASAP7_75t_L g1659 ( .A1(n_878), .A2(n_1169), .B1(n_1654), .B2(n_1656), .C1(n_1660), .C2(n_1661), .Y(n_1659) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_882), .A2(n_898), .B1(n_899), .B2(n_902), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_889), .B1(n_890), .B2(n_892), .Y(n_883) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g1017 ( .A(n_886), .Y(n_1017) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g1173 ( .A(n_887), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1257 ( .A(n_887), .Y(n_1257) );
HB1xp67_ASAP7_75t_L g1960 ( .A(n_893), .Y(n_1960) );
NAND3xp33_ASAP7_75t_SL g894 ( .A(n_895), .B(n_897), .C(n_903), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1671 ( .A1(n_899), .A2(n_1634), .B1(n_1667), .B2(n_1668), .Y(n_1671) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
INVx2_ASAP7_75t_L g920 ( .A(n_900), .Y(n_920) );
INVx2_ASAP7_75t_L g1432 ( .A(n_900), .Y(n_1432) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_901), .Y(n_1209) );
NOR2xp33_ASAP7_75t_SL g903 ( .A(n_904), .B(n_907), .Y(n_903) );
OAI33xp33_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_910), .A3(n_914), .B1(n_919), .B2(n_923), .B3(n_926), .Y(n_907) );
BUFx4f_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx8_ASAP7_75t_L g1188 ( .A(n_909), .Y(n_1188) );
BUFx2_ASAP7_75t_L g1934 ( .A(n_909), .Y(n_1934) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_914) );
INVx8_ASAP7_75t_L g1028 ( .A(n_916), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1554 ( .A1(n_916), .A2(n_1555), .B1(n_1556), .B2(n_1557), .C(n_1558), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_917), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_920), .A2(n_950), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
NAND4xp75_ASAP7_75t_L g928 ( .A(n_929), .B(n_971), .C(n_988), .D(n_989), .Y(n_928) );
OAI21x1_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_944), .B(n_969), .Y(n_929) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_933), .B(n_939), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_932), .A2(n_1002), .B1(n_1034), .B2(n_1037), .Y(n_1033) );
AOI221xp5_ASAP7_75t_SL g933 ( .A1(n_934), .A2(n_935), .B1(n_936), .B2(n_937), .C(n_938), .Y(n_933) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_941), .B(n_942), .C(n_943), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_951), .B1(n_957), .B2(n_963), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_949), .B2(n_950), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_946), .A2(n_958), .B1(n_975), .B2(n_977), .Y(n_974) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_950), .A2(n_1194), .B1(n_1195), .B2(n_1196), .C(n_1197), .Y(n_1193) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g965 ( .A(n_954), .Y(n_965) );
INVx2_ASAP7_75t_L g1056 ( .A(n_954), .Y(n_1056) );
INVx2_ASAP7_75t_L g1909 ( .A(n_954), .Y(n_1909) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_955), .A2(n_1328), .B1(n_1329), .B2(n_1330), .Y(n_1327) );
BUFx4f_ASAP7_75t_SL g959 ( .A(n_960), .Y(n_959) );
INVx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx2_ASAP7_75t_SL g1208 ( .A(n_961), .Y(n_1208) );
OAI21xp33_ASAP7_75t_L g1105 ( .A1(n_965), .A2(n_1106), .B(n_1107), .Y(n_1105) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
OAI31xp33_ASAP7_75t_L g1428 ( .A1(n_969), .A2(n_1429), .A3(n_1430), .B(n_1441), .Y(n_1428) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AOI211x1_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B(n_978), .C(n_984), .Y(n_971) );
BUFx3_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
BUFx3_ASAP7_75t_L g1090 ( .A(n_976), .Y(n_1090) );
BUFx6f_ASAP7_75t_L g1133 ( .A(n_976), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1143 ( .A(n_976), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_977), .A2(n_980), .B1(n_1110), .B2(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_1043), .B1(n_1044), .B2(n_1093), .Y(n_992) );
INVx1_ASAP7_75t_L g1093 ( .A(n_993), .Y(n_1093) );
OAI21x1_ASAP7_75t_SL g993 ( .A1(n_994), .A2(n_995), .B(n_1042), .Y(n_993) );
NAND4xp25_ASAP7_75t_L g1042 ( .A(n_994), .B(n_997), .C(n_999), .D(n_1019), .Y(n_1042) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_999), .C(n_1019), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1005), .Y(n_999) );
NAND3xp33_ASAP7_75t_SL g1005 ( .A(n_1006), .B(n_1009), .C(n_1012), .Y(n_1005) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
NAND3xp33_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1025), .C(n_1033), .Y(n_1020) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .B1(n_1029), .B2(n_1030), .Y(n_1025) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OAI21xp5_ASAP7_75t_L g1614 ( .A1(n_1032), .A2(n_1615), .B(n_1616), .Y(n_1614) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
NOR2x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1070), .Y(n_1045) );
A2O1A1Ixp33_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1051), .B(n_1067), .C(n_1068), .Y(n_1046) );
NOR3xp33_ASAP7_75t_SL g1051 ( .A(n_1052), .B(n_1060), .C(n_1061), .Y(n_1051) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_1058), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1089) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1078), .Y(n_1070) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
OAI33xp33_ASAP7_75t_L g1346 ( .A1(n_1084), .A2(n_1347), .A3(n_1350), .B1(n_1352), .B2(n_1357), .B3(n_1358), .Y(n_1346) );
OAI33xp33_ASAP7_75t_L g1918 ( .A1(n_1084), .A2(n_1357), .A3(n_1919), .B1(n_1922), .B2(n_1925), .B3(n_1930), .Y(n_1918) );
BUFx2_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1088), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_1090), .A2(n_1261), .B1(n_1330), .B2(n_1359), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_1092), .A2(n_1328), .B1(n_1335), .B2(n_1351), .Y(n_1350) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .B1(n_1215), .B2(n_1216), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_1097), .A2(n_1151), .B1(n_1152), .B2(n_1214), .Y(n_1096) );
BUFx2_ASAP7_75t_SL g1097 ( .A(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1098), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1127), .Y(n_1099) );
OAI21xp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1108), .B(n_1114), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_1106), .A2(n_1115), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1110), .B1(n_1111), .B2(n_1113), .Y(n_1108) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_1113), .A2(n_1135), .B1(n_1142), .B2(n_1144), .Y(n_1141) );
OAI211xp5_ASAP7_75t_L g1114 ( .A1(n_1115), .A2(n_1116), .B(n_1117), .C(n_1118), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1126), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1148), .C(n_1150), .Y(n_1127) );
NOR2xp33_ASAP7_75t_SL g1128 ( .A(n_1129), .B(n_1147), .Y(n_1128) );
OAI33xp33_ASAP7_75t_L g1129 ( .A1(n_1130), .A2(n_1131), .A3(n_1136), .B1(n_1138), .B2(n_1141), .B3(n_1145), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_1132), .A2(n_1133), .B1(n_1134), .B2(n_1135), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1919 ( .A1(n_1133), .A2(n_1423), .B1(n_1920), .B2(n_1921), .Y(n_1919) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_1135), .A2(n_1384), .B1(n_1394), .B2(n_1395), .Y(n_1393) );
OAI22xp5_ASAP7_75t_SL g1922 ( .A1(n_1139), .A2(n_1356), .B1(n_1923), .B2(n_1924), .Y(n_1922) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1146), .Y(n_1357) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
XNOR2x1_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1154), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1202), .Y(n_1154) );
NAND3xp33_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1168), .C(n_1177), .Y(n_1158) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
AOI222xp33_ASAP7_75t_L g1306 ( .A1(n_1169), .A2(n_1283), .B1(n_1284), .B2(n_1307), .C1(n_1310), .C2(n_1311), .Y(n_1306) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_1178), .A2(n_1297), .B1(n_1298), .B2(n_1299), .Y(n_1296) );
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_1180), .A2(n_1203), .B1(n_1204), .B2(n_1205), .C(n_1206), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1184), .B1(n_1186), .B2(n_1187), .Y(n_1182) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_1187), .A2(n_1229), .B1(n_1231), .B2(n_1232), .C(n_1233), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1237 ( .A1(n_1187), .A2(n_1238), .B1(n_1239), .B2(n_1240), .C(n_1241), .Y(n_1237) );
OAI33xp33_ASAP7_75t_L g1449 ( .A1(n_1188), .A2(n_1450), .A3(n_1453), .B1(n_1456), .B2(n_1459), .B3(n_1460), .Y(n_1449) );
CKINVDCx20_ASAP7_75t_R g1616 ( .A(n_1188), .Y(n_1616) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
BUFx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
BUFx2_ASAP7_75t_L g1292 ( .A(n_1200), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1278 ( .A1(n_1203), .A2(n_1204), .B1(n_1279), .B2(n_1280), .C(n_1281), .Y(n_1278) );
AOI221xp5_ASAP7_75t_L g1639 ( .A1(n_1203), .A2(n_1204), .B1(n_1640), .B2(n_1641), .C(n_1642), .Y(n_1639) );
AOI21xp5_ASAP7_75t_L g1629 ( .A1(n_1204), .A2(n_1630), .B(n_1631), .Y(n_1629) );
AOI21xp5_ASAP7_75t_L g1974 ( .A1(n_1204), .A2(n_1975), .B(n_1976), .Y(n_1974) );
OR2x6_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1230 ( .A(n_1208), .Y(n_1230) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND3xp33_ASAP7_75t_SL g1281 ( .A(n_1213), .B(n_1282), .C(n_1285), .Y(n_1281) );
INVx2_ASAP7_75t_SL g1991 ( .A(n_1213), .Y(n_1991) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
OA22x2_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1274), .B1(n_1275), .B2(n_1360), .Y(n_1216) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1217), .Y(n_1360) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NOR2x1_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1246), .Y(n_1219) );
NAND3xp33_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1237), .C(n_1243), .Y(n_1227) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1263), .Y(n_1246) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_SL g1253 ( .A(n_1254), .Y(n_1253) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1262), .Y(n_1581) );
AOI21xp5_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B(n_1267), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1265), .B(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1316), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1294), .Y(n_1277) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
AOI21xp5_ASAP7_75t_SL g1294 ( .A1(n_1295), .A2(n_1313), .B(n_1314), .Y(n_1294) );
NAND3xp33_ASAP7_75t_SL g1295 ( .A(n_1296), .B(n_1300), .C(n_1306), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g1963 ( .A(n_1298), .Y(n_1963) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
A2O1A1Ixp33_ASAP7_75t_SL g1367 ( .A1(n_1313), .A2(n_1368), .B(n_1372), .C(n_1385), .Y(n_1367) );
AOI211x1_ASAP7_75t_L g1317 ( .A1(n_1318), .A2(n_1336), .B(n_1338), .C(n_1344), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1323), .Y(n_1318) );
NOR3xp33_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1331), .C(n_1332), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1936 ( .A1(n_1329), .A2(n_1923), .B1(n_1931), .B2(n_1937), .Y(n_1936) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_1334), .A2(n_1353), .B1(n_1355), .B2(n_1356), .Y(n_1352) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1348), .Y(n_1494) );
INVx4_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1361), .Y(n_1673) );
AOI22xp5_ASAP7_75t_L g1361 ( .A1(n_1362), .A2(n_1363), .B1(n_1588), .B2(n_1589), .Y(n_1361) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
XOR2x2_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1444), .Y(n_1363) );
XOR2xp5_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1404), .Y(n_1364) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1387), .Y(n_1366) );
NOR3xp33_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1379), .C(n_1380), .Y(n_1372) );
NAND3xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .C(n_1402), .Y(n_1387) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
XOR2x2_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1443), .Y(n_1404) );
NAND3xp33_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1412), .C(n_1425), .Y(n_1407) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
OAI22xp5_ASAP7_75t_L g1418 ( .A1(n_1419), .A2(n_1420), .B1(n_1422), .B2(n_1423), .Y(n_1418) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
NAND3xp33_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1435), .C(n_1440), .Y(n_1430) );
OAI211xp5_ASAP7_75t_L g1435 ( .A1(n_1436), .A2(n_1437), .B(n_1438), .C(n_1439), .Y(n_1435) );
AOI22xp5_ASAP7_75t_L g1444 ( .A1(n_1445), .A2(n_1446), .B1(n_1542), .B2(n_1543), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
XOR2x2_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1541), .Y(n_1446) );
AND3x1_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1477), .C(n_1508), .Y(n_1447) );
NOR2xp33_ASAP7_75t_SL g1448 ( .A(n_1449), .B(n_1463), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1468 ( .A1(n_1452), .A2(n_1462), .B1(n_1469), .B2(n_1471), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g1474 ( .A1(n_1455), .A2(n_1458), .B1(n_1466), .B2(n_1475), .Y(n_1474) );
OAI33xp33_ASAP7_75t_L g1463 ( .A1(n_1464), .A2(n_1465), .A3(n_1467), .B1(n_1468), .B2(n_1473), .B3(n_1474), .Y(n_1463) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx5_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
BUFx3_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
OAI31xp33_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1482), .A3(n_1492), .B(n_1505), .Y(n_1477) );
INVx4_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
CKINVDCx16_ASAP7_75t_R g1901 ( .A(n_1480), .Y(n_1901) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
BUFx6f_ASAP7_75t_L g1896 ( .A(n_1485), .Y(n_1896) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx2_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx2_ASAP7_75t_L g1898 ( .A(n_1490), .Y(n_1898) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx3_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1500), .B1(n_1501), .B2(n_1504), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_1500), .A2(n_1522), .B1(n_1526), .B2(n_1529), .Y(n_1521) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
AOI22xp33_ASAP7_75t_L g1891 ( .A1(n_1503), .A2(n_1892), .B1(n_1893), .B2(n_1894), .Y(n_1891) );
BUFx3_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
BUFx2_ASAP7_75t_SL g1902 ( .A(n_1506), .Y(n_1902) );
OAI31xp33_ASAP7_75t_L g1508 ( .A1(n_1509), .A2(n_1516), .A3(n_1530), .B(n_1536), .Y(n_1508) );
INVx2_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVx2_ASAP7_75t_SL g1511 ( .A(n_1512), .Y(n_1511) );
INVx2_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1915 ( .A(n_1514), .Y(n_1915) );
INVxp67_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
CKINVDCx8_ASAP7_75t_R g1519 ( .A(n_1520), .Y(n_1519) );
CKINVDCx8_ASAP7_75t_R g1910 ( .A(n_1520), .Y(n_1910) );
BUFx3_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1525), .Y(n_1523) );
AND2x4_ASAP7_75t_L g1527 ( .A(n_1524), .B(n_1528), .Y(n_1527) );
AND2x4_ASAP7_75t_L g1912 ( .A(n_1524), .B(n_1525), .Y(n_1912) );
BUFx6f_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g1911 ( .A1(n_1527), .A2(n_1892), .B1(n_1912), .B2(n_1913), .Y(n_1911) );
BUFx2_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
BUFx2_ASAP7_75t_L g1905 ( .A(n_1532), .Y(n_1905) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx2_ASAP7_75t_L g1906 ( .A(n_1534), .Y(n_1906) );
INVx2_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
AND2x2_ASAP7_75t_SL g1536 ( .A(n_1537), .B(n_1539), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1916 ( .A(n_1537), .B(n_1539), .Y(n_1916) );
INVx1_ASAP7_75t_SL g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1544), .Y(n_1586) );
NAND4xp25_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1569), .C(n_1571), .D(n_1585), .Y(n_1544) );
NAND3xp33_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1562), .C(n_1566), .Y(n_1553) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1580), .Y(n_1571) );
NAND3xp33_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1578), .C(n_1579), .Y(n_1573) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
CKINVDCx5p33_ASAP7_75t_R g1588 ( .A(n_1589), .Y(n_1588) );
AO22x1_ASAP7_75t_L g1589 ( .A1(n_1590), .A2(n_1635), .B1(n_1636), .B2(n_1672), .Y(n_1589) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1590), .Y(n_1672) );
HB1xp67_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
AND4x1_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1612), .C(n_1629), .D(n_1633), .Y(n_1592) );
INVx2_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
OAI211xp5_ASAP7_75t_L g1605 ( .A1(n_1606), .A2(n_1607), .B(n_1608), .C(n_1609), .Y(n_1605) );
OAI22xp5_ASAP7_75t_L g1613 ( .A1(n_1614), .A2(n_1617), .B1(n_1620), .B2(n_1623), .Y(n_1613) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
HB1xp67_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1657), .Y(n_1638) );
NAND3xp33_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1644), .C(n_1653), .Y(n_1642) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
OAI33xp33_ASAP7_75t_L g1933 ( .A1(n_1652), .A2(n_1934), .A3(n_1935), .B1(n_1936), .B2(n_1938), .B3(n_1940), .Y(n_1933) );
AOI21xp5_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1669), .B(n_1670), .Y(n_1657) );
NAND3xp33_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1662), .C(n_1666), .Y(n_1658) );
OAI221xp5_ASAP7_75t_L g1674 ( .A1(n_1675), .A2(n_1885), .B1(n_1887), .B2(n_1941), .C(n_1944), .Y(n_1674) );
NOR3xp33_ASAP7_75t_L g1675 ( .A(n_1676), .B(n_1847), .C(n_1860), .Y(n_1675) );
NAND4xp25_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1775), .C(n_1797), .D(n_1830), .Y(n_1676) );
OAI31xp33_ASAP7_75t_L g1677 ( .A1(n_1678), .A2(n_1729), .A3(n_1759), .B(n_1768), .Y(n_1677) );
OAI21xp33_ASAP7_75t_L g1678 ( .A1(n_1679), .A2(n_1700), .B(n_1718), .Y(n_1678) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1680), .B(n_1795), .Y(n_1794) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_1680), .B(n_1804), .Y(n_1803) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1696), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1681), .B(n_1742), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1681), .B(n_1724), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1681), .B(n_1766), .Y(n_1765) );
OR2x2_ASAP7_75t_L g1790 ( .A(n_1681), .B(n_1696), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1801 ( .A(n_1681), .B(n_1768), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1812 ( .A(n_1681), .B(n_1733), .Y(n_1812) );
NAND3xp33_ASAP7_75t_L g1842 ( .A(n_1681), .B(n_1737), .C(n_1843), .Y(n_1842) );
CKINVDCx6p67_ASAP7_75t_R g1681 ( .A(n_1682), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1730 ( .A(n_1682), .B(n_1731), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1782 ( .A(n_1682), .B(n_1696), .Y(n_1782) );
OR2x2_ASAP7_75t_L g1791 ( .A(n_1682), .B(n_1696), .Y(n_1791) );
CKINVDCx5p33_ASAP7_75t_R g1816 ( .A(n_1682), .Y(n_1816) );
NAND2xp5_ASAP7_75t_L g1828 ( .A(n_1682), .B(n_1769), .Y(n_1828) );
OR2x6_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1690), .Y(n_1682) );
OR2x2_ASAP7_75t_L g1809 ( .A(n_1683), .B(n_1690), .Y(n_1809) );
INVx2_ASAP7_75t_L g1772 ( .A(n_1684), .Y(n_1772) );
AND2x6_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1686), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1685), .B(n_1689), .Y(n_1688) );
AND2x4_ASAP7_75t_L g1691 ( .A(n_1685), .B(n_1692), .Y(n_1691) );
AND2x6_ASAP7_75t_L g1694 ( .A(n_1685), .B(n_1695), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1685), .B(n_1689), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1685), .B(n_1689), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1687), .B(n_1693), .Y(n_1692) );
OAI21xp5_ASAP7_75t_L g1995 ( .A1(n_1689), .A2(n_1996), .B(n_1997), .Y(n_1995) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1696), .B(n_1726), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1696), .B(n_1733), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1696), .B(n_1726), .Y(n_1758) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1696), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1837 ( .A(n_1696), .B(n_1838), .Y(n_1837) );
INVx3_ASAP7_75t_L g1853 ( .A(n_1696), .Y(n_1853) );
OAI21xp5_ASAP7_75t_L g1863 ( .A1(n_1696), .A2(n_1778), .B(n_1864), .Y(n_1863) );
AND2x4_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1699), .Y(n_1696) );
INVxp67_ASAP7_75t_L g1774 ( .A(n_1698), .Y(n_1774) );
HB1xp67_ASAP7_75t_L g1886 ( .A(n_1698), .Y(n_1886) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1700), .Y(n_1858) );
OR2x2_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1706), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1701), .B(n_1707), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1781 ( .A(n_1701), .B(n_1756), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1800 ( .A(n_1701), .B(n_1719), .Y(n_1800) );
NAND2xp5_ASAP7_75t_L g1827 ( .A(n_1701), .B(n_1720), .Y(n_1827) );
OR2x2_ASAP7_75t_L g1832 ( .A(n_1701), .B(n_1833), .Y(n_1832) );
AND3x1_ASAP7_75t_L g1868 ( .A(n_1701), .B(n_1715), .C(n_1720), .Y(n_1868) );
INVx2_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
BUFx2_ASAP7_75t_L g1740 ( .A(n_1702), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1702), .B(n_1756), .Y(n_1763) );
OR2x2_ASAP7_75t_L g1821 ( .A(n_1702), .B(n_1822), .Y(n_1821) );
OR2x2_ASAP7_75t_L g1865 ( .A(n_1702), .B(n_1745), .Y(n_1865) );
AND2x2_ASAP7_75t_L g1874 ( .A(n_1702), .B(n_1711), .Y(n_1874) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1704), .Y(n_1702) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1706), .Y(n_1882) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1711), .Y(n_1706) );
NOR2xp33_ASAP7_75t_L g1735 ( .A(n_1707), .B(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1707), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1751 ( .A(n_1707), .B(n_1742), .Y(n_1751) );
NOR2xp33_ASAP7_75t_L g1819 ( .A(n_1707), .B(n_1820), .Y(n_1819) );
NAND2xp5_ASAP7_75t_L g1841 ( .A(n_1707), .B(n_1750), .Y(n_1841) );
INVx2_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1708), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1745 ( .A(n_1708), .B(n_1711), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1708), .B(n_1740), .Y(n_1757) );
NOR2xp33_ASAP7_75t_L g1804 ( .A(n_1708), .B(n_1805), .Y(n_1804) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1708), .B(n_1733), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1838 ( .A(n_1708), .B(n_1726), .Y(n_1838) );
OR2x2_ASAP7_75t_L g1844 ( .A(n_1708), .B(n_1726), .Y(n_1844) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1709), .B(n_1710), .Y(n_1708) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1711), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1715), .Y(n_1711) );
INVx2_ASAP7_75t_L g1720 ( .A(n_1712), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1712), .B(n_1721), .Y(n_1756) );
OR2x2_ASAP7_75t_L g1712 ( .A(n_1713), .B(n_1714), .Y(n_1712) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1715), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1715), .B(n_1720), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1715), .B(n_1740), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1820 ( .A(n_1715), .B(n_1740), .Y(n_1820) );
AOI32xp33_ASAP7_75t_L g1836 ( .A1(n_1715), .A2(n_1816), .A3(n_1837), .B1(n_1839), .B2(n_1840), .Y(n_1836) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1717), .Y(n_1715) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1722), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1753 ( .A(n_1719), .B(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1719), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1833 ( .A(n_1719), .B(n_1723), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1720), .B(n_1721), .Y(n_1719) );
OR2x2_ASAP7_75t_L g1805 ( .A(n_1720), .B(n_1740), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_1720), .B(n_1740), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1721), .B(n_1740), .Y(n_1739) );
OAI211xp5_ASAP7_75t_L g1806 ( .A1(n_1722), .A2(n_1807), .B(n_1808), .C(n_1809), .Y(n_1806) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1724), .Y(n_1722) );
INVx2_ASAP7_75t_L g1762 ( .A(n_1723), .Y(n_1762) );
INVx2_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
AOI211xp5_ASAP7_75t_L g1824 ( .A1(n_1725), .A2(n_1762), .B(n_1816), .C(n_1825), .Y(n_1824) );
OAI22xp5_ASAP7_75t_L g1848 ( .A1(n_1725), .A2(n_1849), .B1(n_1853), .B2(n_1854), .Y(n_1848) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1726), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1726), .B(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1728), .Y(n_1726) );
OAI211xp5_ASAP7_75t_SL g1729 ( .A1(n_1730), .A2(n_1734), .B(n_1738), .C(n_1752), .Y(n_1729) );
OAI21xp5_ASAP7_75t_L g1759 ( .A1(n_1731), .A2(n_1760), .B(n_1764), .Y(n_1759) );
A2O1A1Ixp33_ASAP7_75t_L g1869 ( .A1(n_1731), .A2(n_1845), .B(n_1870), .C(n_1871), .Y(n_1869) );
CKINVDCx6p67_ASAP7_75t_R g1731 ( .A(n_1732), .Y(n_1731) );
AOI31xp33_ASAP7_75t_L g1813 ( .A1(n_1732), .A2(n_1757), .A3(n_1814), .B(n_1816), .Y(n_1813) );
INVx2_ASAP7_75t_L g1742 ( .A(n_1733), .Y(n_1742) );
OAI211xp5_ASAP7_75t_SL g1835 ( .A1(n_1734), .A2(n_1790), .B(n_1836), .C(n_1842), .Y(n_1835) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
AOI211xp5_ASAP7_75t_L g1826 ( .A1(n_1736), .A2(n_1827), .B(n_1828), .C(n_1829), .Y(n_1826) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1737), .B(n_1754), .Y(n_1793) );
OR2x2_ASAP7_75t_L g1815 ( .A(n_1737), .B(n_1756), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1879 ( .A(n_1737), .B(n_1740), .Y(n_1879) );
AOI321xp33_ASAP7_75t_L g1738 ( .A1(n_1739), .A2(n_1741), .A3(n_1743), .B1(n_1744), .B2(n_1746), .C(n_1748), .Y(n_1738) );
AOI221xp5_ASAP7_75t_L g1810 ( .A1(n_1741), .A2(n_1792), .B1(n_1811), .B2(n_1812), .C(n_1813), .Y(n_1810) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1741), .Y(n_1834) );
INVx2_ASAP7_75t_L g1779 ( .A(n_1742), .Y(n_1779) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
AOI21xp33_ASAP7_75t_SL g1831 ( .A1(n_1745), .A2(n_1832), .B(n_1834), .Y(n_1831) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
NOR2xp33_ASAP7_75t_L g1748 ( .A(n_1749), .B(n_1751), .Y(n_1748) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
OAI21xp33_ASAP7_75t_L g1752 ( .A1(n_1753), .A2(n_1755), .B(n_1758), .Y(n_1752) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1753), .B(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1753), .Y(n_1811) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1755), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_1756), .B(n_1757), .Y(n_1755) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1756), .B(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1757), .Y(n_1788) );
INVx2_ASAP7_75t_L g1859 ( .A(n_1758), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1761), .B(n_1763), .Y(n_1760) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1762), .B(n_1781), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1852 ( .A(n_1762), .B(n_1800), .Y(n_1852) );
AND2x2_ASAP7_75t_L g1867 ( .A(n_1762), .B(n_1868), .Y(n_1867) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1763), .Y(n_1825) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1765), .Y(n_1823) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1766), .Y(n_1857) );
AOI211xp5_ASAP7_75t_L g1873 ( .A1(n_1766), .A2(n_1776), .B(n_1874), .C(n_1875), .Y(n_1873) );
OAI32xp33_ASAP7_75t_L g1880 ( .A1(n_1767), .A2(n_1845), .A3(n_1881), .B1(n_1882), .B2(n_1883), .Y(n_1880) );
OAI321xp33_ASAP7_75t_L g1798 ( .A1(n_1768), .A2(n_1778), .A3(n_1799), .B1(n_1801), .B2(n_1802), .C(n_1806), .Y(n_1798) );
INVx2_ASAP7_75t_SL g1768 ( .A(n_1769), .Y(n_1768) );
INVx2_ASAP7_75t_SL g1846 ( .A(n_1769), .Y(n_1846) );
OAI22xp5_ASAP7_75t_SL g1770 ( .A1(n_1771), .A2(n_1772), .B1(n_1773), .B2(n_1774), .Y(n_1770) );
O2A1O1Ixp33_ASAP7_75t_L g1775 ( .A1(n_1776), .A2(n_1780), .B(n_1782), .C(n_1783), .Y(n_1775) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1778), .B(n_1786), .Y(n_1785) );
A2O1A1Ixp33_ASAP7_75t_L g1861 ( .A1(n_1778), .A2(n_1804), .B(n_1853), .C(n_1862), .Y(n_1861) );
INVx2_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
NOR2xp33_ASAP7_75t_L g1795 ( .A(n_1779), .B(n_1796), .Y(n_1795) );
NAND2xp5_ASAP7_75t_L g1850 ( .A(n_1779), .B(n_1851), .Y(n_1850) );
NAND2xp5_ASAP7_75t_L g1855 ( .A(n_1779), .B(n_1780), .Y(n_1855) );
AOI21xp33_ASAP7_75t_SL g1866 ( .A1(n_1779), .A2(n_1867), .B(n_1869), .Y(n_1866) );
OAI221xp5_ASAP7_75t_L g1783 ( .A1(n_1784), .A2(n_1790), .B1(n_1791), .B2(n_1792), .C(n_1794), .Y(n_1783) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1788), .B(n_1789), .Y(n_1787) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1791), .Y(n_1839) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1793), .Y(n_1792) );
NOR5xp2_ASAP7_75t_SL g1797 ( .A(n_1798), .B(n_1810), .C(n_1817), .D(n_1824), .E(n_1826), .Y(n_1797) );
NAND2xp5_ASAP7_75t_L g1877 ( .A(n_1799), .B(n_1878), .Y(n_1877) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1801), .Y(n_1884) );
INVxp67_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1805), .Y(n_1808) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
AOI21xp33_ASAP7_75t_SL g1817 ( .A1(n_1818), .A2(n_1821), .B(n_1823), .Y(n_1817) );
INVxp33_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1821), .Y(n_1881) );
O2A1O1Ixp33_ASAP7_75t_L g1847 ( .A1(n_1825), .A2(n_1828), .B(n_1848), .C(n_1856), .Y(n_1847) );
OAI211xp5_ASAP7_75t_L g1862 ( .A1(n_1825), .A2(n_1844), .B(n_1852), .C(n_1863), .Y(n_1862) );
OAI21xp5_ASAP7_75t_L g1830 ( .A1(n_1831), .A2(n_1835), .B(n_1845), .Y(n_1830) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1833), .Y(n_1872) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1844), .Y(n_1843) );
INVx3_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
NAND2xp5_ASAP7_75t_L g1883 ( .A(n_1846), .B(n_1853), .Y(n_1883) );
INVxp67_ASAP7_75t_L g1849 ( .A(n_1850), .Y(n_1849) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
AOI221xp5_ASAP7_75t_L g1860 ( .A1(n_1855), .A2(n_1861), .B1(n_1866), .B2(n_1873), .C(n_1884), .Y(n_1860) );
OAI21xp5_ASAP7_75t_SL g1856 ( .A1(n_1857), .A2(n_1858), .B(n_1859), .Y(n_1856) );
OAI21xp5_ASAP7_75t_SL g1875 ( .A1(n_1859), .A2(n_1876), .B(n_1880), .Y(n_1875) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
INVx2_ASAP7_75t_L g1870 ( .A(n_1868), .Y(n_1870) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1879), .Y(n_1878) );
INVx4_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
NAND3xp33_ASAP7_75t_L g1888 ( .A(n_1889), .B(n_1903), .C(n_1917), .Y(n_1888) );
OAI31xp33_ASAP7_75t_L g1889 ( .A1(n_1890), .A2(n_1895), .A3(n_1899), .B(n_1902), .Y(n_1889) );
INVx2_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
OAI31xp33_ASAP7_75t_L g1903 ( .A1(n_1904), .A2(n_1907), .A3(n_1914), .B(n_1916), .Y(n_1903) );
HB1xp67_ASAP7_75t_L g1908 ( .A(n_1909), .Y(n_1908) );
NOR2xp33_ASAP7_75t_SL g1917 ( .A(n_1918), .B(n_1933), .Y(n_1917) );
OAI22xp5_ASAP7_75t_L g1925 ( .A1(n_1926), .A2(n_1927), .B1(n_1928), .B2(n_1929), .Y(n_1925) );
INVx3_ASAP7_75t_L g1941 ( .A(n_1942), .Y(n_1941) );
HB1xp67_ASAP7_75t_L g1945 ( .A(n_1946), .Y(n_1945) );
BUFx3_ASAP7_75t_L g1946 ( .A(n_1947), .Y(n_1946) );
INVx1_ASAP7_75t_SL g1948 ( .A(n_1949), .Y(n_1948) );
INVx1_ASAP7_75t_L g1951 ( .A(n_1952), .Y(n_1951) );
INVx1_ASAP7_75t_L g1952 ( .A(n_1953), .Y(n_1952) );
INVx1_ASAP7_75t_L g1992 ( .A(n_1953), .Y(n_1992) );
INVx1_ASAP7_75t_L g1953 ( .A(n_1954), .Y(n_1953) );
NAND3xp33_ASAP7_75t_SL g1954 ( .A(n_1955), .B(n_1974), .C(n_1977), .Y(n_1954) );
OAI21xp33_ASAP7_75t_L g1955 ( .A1(n_1956), .A2(n_1965), .B(n_1973), .Y(n_1955) );
NOR3xp33_ASAP7_75t_L g1977 ( .A(n_1978), .B(n_1989), .C(n_1991), .Y(n_1977) );
NAND2xp5_ASAP7_75t_L g1978 ( .A(n_1979), .B(n_1982), .Y(n_1978) );
INVx1_ASAP7_75t_L g1985 ( .A(n_1986), .Y(n_1985) );
INVx1_ASAP7_75t_L g1993 ( .A(n_1994), .Y(n_1993) );
INVx1_ASAP7_75t_L g1994 ( .A(n_1995), .Y(n_1994) );
INVx1_ASAP7_75t_L g1997 ( .A(n_1998), .Y(n_1997) );
endmodule