module fake_jpeg_1223_n_112 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_40),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_43),
.B1(n_31),
.B2(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_64),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_52),
.B1(n_51),
.B2(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_0),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_35),
.C(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_69),
.B(n_4),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_35),
.B1(n_31),
.B2(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_55),
.B1(n_62),
.B2(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_56),
.B1(n_5),
.B2(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_15),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_74),
.B1(n_72),
.B2(n_9),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_16),
.Y(n_80)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.C(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_85),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_56),
.B(n_5),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_7),
.B(n_8),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_4),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_86),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_18),
.C(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_93),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_96),
.B1(n_76),
.B2(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_92),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_74),
.B(n_13),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_14),
.B(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_80),
.B1(n_9),
.B2(n_10),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_8),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_23),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_100),
.C(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_97),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_103),
.B1(n_102),
.B2(n_96),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_93),
.A3(n_95),
.B1(n_102),
.B2(n_92),
.C1(n_87),
.C2(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_10),
.Y(n_112)
);


endmodule