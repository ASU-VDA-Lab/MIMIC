module fake_jpeg_792_n_184 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_51),
.B1(n_60),
.B2(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_51),
.B1(n_69),
.B2(n_46),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_70),
.Y(n_99)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_68),
.C(n_59),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_56),
.C(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_92),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_93),
.B1(n_45),
.B2(n_50),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_65),
.B1(n_61),
.B2(n_71),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_75),
.B1(n_84),
.B2(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_58),
.C(n_53),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_70),
.B1(n_71),
.B2(n_55),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_4),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_84),
.B1(n_45),
.B2(n_48),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_115),
.B1(n_20),
.B2(n_40),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_113),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_84),
.B(n_45),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_102),
.B(n_105),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_45),
.B1(n_48),
.B2(n_2),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_25),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_0),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_9),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_112),
.B1(n_116),
.B2(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_27),
.B(n_37),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_22),
.C(n_42),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_10),
.C(n_11),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_6),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_7),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_139),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_145),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_15),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_13),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_156),
.B1(n_12),
.B2(n_13),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_26),
.C(n_34),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_155),
.C(n_19),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_125),
.B1(n_126),
.B2(n_14),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_145),
.C(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_160),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_155),
.C(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

AOI31xp67_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_162),
.A3(n_159),
.B(n_157),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_164),
.B1(n_146),
.B2(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_154),
.C(n_158),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_166),
.B(n_175),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_171),
.C(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_148),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_156),
.B(n_28),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_17),
.B(n_30),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_33),
.Y(n_184)
);


endmodule