module fake_jpeg_29952_n_516 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_516);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_516;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_9),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_55),
.Y(n_151)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g106 ( 
.A(n_57),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_18),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_32),
.B(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_34),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_8),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_94),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_27),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_77),
.A2(n_33),
.B1(n_44),
.B2(n_20),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_32),
.B(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_49),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_38),
.B(n_10),
.CON(n_80),
.SN(n_80)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_82),
.Y(n_120)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_33),
.B(n_7),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_22),
.B1(n_37),
.B2(n_29),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_102),
.A2(n_131),
.B1(n_140),
.B2(n_64),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_40),
.B1(n_22),
.B2(n_37),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_119),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_40),
.B1(n_37),
.B2(n_29),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_113),
.B(n_13),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_40),
.B1(n_29),
.B2(n_45),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_50),
.A2(n_40),
.B1(n_45),
.B2(n_36),
.Y(n_119)
);

BUFx4f_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_75),
.B(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_148),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_20),
.B1(n_44),
.B2(n_45),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_52),
.B1(n_63),
.B2(n_60),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_36),
.B1(n_48),
.B2(n_39),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_154),
.B1(n_156),
.B2(n_78),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_36),
.B1(n_48),
.B2(n_39),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_147),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_26),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_97),
.A2(n_48),
.B1(n_26),
.B2(n_46),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_91),
.A2(n_46),
.B1(n_43),
.B2(n_11),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_82),
.B(n_46),
.C(n_88),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_160),
.A2(n_211),
.B(n_172),
.C(n_181),
.Y(n_237)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_164),
.B(n_172),
.Y(n_225)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_168),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx5_ASAP7_75t_SL g262 ( 
.A(n_169),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_171),
.B(n_211),
.Y(n_252)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_110),
.A2(n_124),
.A3(n_121),
.B1(n_147),
.B2(n_116),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_174),
.A2(n_191),
.B1(n_194),
.B2(n_197),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_83),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_178),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_105),
.B(n_82),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_176),
.B(n_204),
.Y(n_249)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_99),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_188),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_180),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_115),
.A2(n_87),
.B1(n_84),
.B2(n_74),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_183),
.A2(n_184),
.B1(n_190),
.B2(n_193),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_55),
.B1(n_69),
.B2(n_51),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_145),
.A2(n_73),
.B1(n_62),
.B2(n_61),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_185),
.Y(n_238)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_111),
.A2(n_57),
.B1(n_54),
.B2(n_46),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_57),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_138),
.A2(n_46),
.B1(n_43),
.B2(n_11),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_127),
.A2(n_43),
.B1(n_7),
.B2(n_13),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_101),
.A2(n_7),
.B1(n_17),
.B2(n_16),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_101),
.A2(n_6),
.B1(n_17),
.B2(n_15),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_127),
.A2(n_43),
.B1(n_6),
.B2(n_13),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_99),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_205),
.Y(n_241)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_109),
.A2(n_43),
.B1(n_6),
.B2(n_14),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_201),
.A2(n_202),
.B1(n_209),
.B2(n_213),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_4),
.B1(n_15),
.B2(n_14),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_14),
.C(n_17),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_139),
.B(n_14),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_117),
.A2(n_125),
.B1(n_151),
.B2(n_108),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_0),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_104),
.Y(n_257)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_217),
.B(n_155),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_119),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_219),
.B1(n_135),
.B2(n_130),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_130),
.A2(n_112),
.B1(n_155),
.B2(n_146),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_120),
.C(n_156),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_254),
.C(n_233),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_228),
.B(n_247),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_176),
.B(n_107),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_204),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_237),
.A2(n_269),
.B(n_215),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_180),
.B1(n_200),
.B2(n_198),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_160),
.A2(n_150),
.B(n_159),
.C(n_146),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_170),
.B(n_159),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_263),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_104),
.C(n_123),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_256),
.B(n_259),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_182),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_163),
.B(n_123),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_182),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_164),
.B(n_165),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_266),
.B(n_212),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_182),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_175),
.A2(n_1),
.B(n_2),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_175),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_270),
.B(n_231),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_222),
.A2(n_161),
.B1(n_178),
.B2(n_237),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_271),
.A2(n_280),
.B1(n_284),
.B2(n_287),
.Y(n_328)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_230),
.A2(n_201),
.B1(n_202),
.B2(n_219),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_275),
.A2(n_282),
.B1(n_303),
.B2(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_278),
.B(n_288),
.Y(n_348)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_222),
.A2(n_209),
.B1(n_194),
.B2(n_193),
.Y(n_280)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_247),
.A2(n_189),
.B1(n_186),
.B2(n_208),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_238),
.A2(n_167),
.B1(n_166),
.B2(n_168),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_297),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_230),
.A2(n_173),
.B1(n_162),
.B2(n_188),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_291),
.A2(n_234),
.B1(n_240),
.B2(n_244),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_214),
.C(n_199),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_293),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_169),
.C(n_179),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_177),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_309),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_268),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_300),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_268),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_315),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_261),
.A2(n_195),
.B1(n_196),
.B2(n_217),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_229),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_305),
.Y(n_323)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_240),
.B1(n_262),
.B2(n_226),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_261),
.A2(n_195),
.B1(n_196),
.B2(n_2),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_2),
.B1(n_3),
.B2(n_212),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_308),
.A2(n_248),
.B1(n_246),
.B2(n_265),
.Y(n_355)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_223),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_263),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_310),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_241),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_311),
.Y(n_341)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_258),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_258),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_238),
.A2(n_212),
.B1(n_250),
.B2(n_242),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_226),
.B1(n_239),
.B2(n_267),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_225),
.B(n_252),
.C(n_253),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_224),
.B(n_232),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_316),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_319),
.A2(n_332),
.B1(n_340),
.B2(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_262),
.B1(n_250),
.B2(n_256),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_255),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_344),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_243),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_335),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_288),
.A2(n_254),
.B(n_236),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_345),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_269),
.B(n_228),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_343),
.B(n_346),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_271),
.A2(n_234),
.B(n_262),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_244),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_277),
.A2(n_235),
.B(n_227),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_270),
.A2(n_235),
.B(n_227),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_354),
.B1(n_289),
.B2(n_300),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_265),
.B(n_251),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_278),
.B(n_231),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_292),
.C(n_293),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_280),
.A2(n_275),
.B1(n_277),
.B2(n_303),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_259),
.B1(n_264),
.B2(n_246),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_355),
.A2(n_276),
.B1(n_283),
.B2(n_279),
.Y(n_357)
);

OAI22x1_ASAP7_75t_L g356 ( 
.A1(n_335),
.A2(n_307),
.B1(n_286),
.B2(n_314),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_357),
.B1(n_380),
.B2(n_383),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_322),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_358),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_370),
.C(n_372),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_325),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_381),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_290),
.B1(n_315),
.B2(n_295),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_364),
.A2(n_365),
.B1(n_368),
.B2(n_369),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_294),
.B1(n_309),
.B2(n_296),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_285),
.B1(n_312),
.B2(n_297),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_248),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_298),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_305),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_322),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_373),
.Y(n_407)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_347),
.Y(n_378)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_324),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_379),
.Y(n_416)
);

OAI22x1_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_281),
.B1(n_272),
.B2(n_273),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_324),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_382),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_353),
.A2(n_274),
.B1(n_304),
.B2(n_306),
.Y(n_383)
);

OAI32xp33_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_251),
.A3(n_344),
.B1(n_350),
.B2(n_333),
.Y(n_384)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_328),
.A2(n_340),
.B1(n_341),
.B2(n_330),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_386),
.A2(n_388),
.B1(n_346),
.B2(n_326),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_352),
.C(n_337),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_348),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_355),
.B1(n_328),
.B2(n_339),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_318),
.B(n_341),
.Y(n_389)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_389),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_348),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_392),
.B(n_409),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_375),
.A2(n_339),
.B1(n_316),
.B2(n_354),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_397),
.A2(n_403),
.B1(n_406),
.B2(n_413),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_389),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_358),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_400),
.B(n_401),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_318),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_390),
.B1(n_405),
.B2(n_415),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_356),
.A2(n_326),
.B1(n_345),
.B2(n_349),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_338),
.B1(n_327),
.B2(n_336),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_338),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_327),
.Y(n_410)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_411),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_371),
.A2(n_334),
.B1(n_336),
.B2(n_323),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_334),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_363),
.C(n_364),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_371),
.A2(n_323),
.B1(n_329),
.B2(n_347),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_418),
.A2(n_383),
.B1(n_403),
.B2(n_369),
.Y(n_424)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_414),
.Y(n_420)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_373),
.Y(n_421)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_418),
.Y(n_456)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_414),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_429),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_424),
.A2(n_377),
.B1(n_412),
.B2(n_404),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_426),
.A2(n_439),
.B1(n_406),
.B2(n_397),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_376),
.B(n_362),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_428),
.A2(n_430),
.B(n_394),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_394),
.A2(n_362),
.B(n_376),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_408),
.C(n_392),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_441),
.C(n_400),
.Y(n_445)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_435),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_407),
.B(n_361),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_434),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_405),
.A2(n_366),
.B1(n_365),
.B2(n_388),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_379),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_436),
.A2(n_440),
.B1(n_443),
.B2(n_395),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_367),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

AOI22x1_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_384),
.B1(n_367),
.B2(n_374),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_363),
.C(n_382),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_449),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_401),
.C(n_417),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_450),
.C(n_445),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_448),
.A2(n_443),
.B1(n_462),
.B2(n_423),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_431),
.C(n_441),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_415),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_457),
.Y(n_473)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_428),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_357),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_412),
.B1(n_404),
.B2(n_385),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_461),
.Y(n_468)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_421),
.A2(n_329),
.B(n_317),
.C(n_321),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_420),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_411),
.B1(n_317),
.B2(n_321),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_425),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_430),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_466),
.B(n_470),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_439),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_447),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_469),
.B(n_438),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_447),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_451),
.B(n_440),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_472),
.B(n_478),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_450),
.B(n_433),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_474),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_479),
.Y(n_487)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_476),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_437),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_460),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_456),
.B(n_439),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_459),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_483),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_476),
.A2(n_449),
.B(n_467),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_481),
.A2(n_458),
.B(n_454),
.Y(n_494)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_477),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_468),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_489),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_490),
.A2(n_471),
.B1(n_453),
.B2(n_435),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_466),
.B(n_448),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_491),
.B(n_492),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_465),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_500),
.C(n_501),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_495),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_484),
.A2(n_473),
.B(n_465),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_452),
.B(n_479),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_499),
.B(n_481),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_446),
.C(n_468),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_496),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_503),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_498),
.B(n_486),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_497),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_509),
.C(n_505),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_490),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_511),
.C(n_509),
.Y(n_512)
);

A2O1A1O1Ixp25_ASAP7_75t_L g511 ( 
.A1(n_508),
.A2(n_482),
.B(n_492),
.C(n_497),
.D(n_483),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_455),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_513),
.A2(n_432),
.B(n_419),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_419),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_463),
.B(n_457),
.Y(n_516)
);


endmodule