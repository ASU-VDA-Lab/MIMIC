module fake_jpeg_20209_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_29),
.B(n_28),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_16),
.B1(n_18),
.B2(n_29),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_47),
.B1(n_31),
.B2(n_38),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_16),
.B1(n_18),
.B2(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_18),
.B1(n_38),
.B2(n_36),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_57),
.B1(n_69),
.B2(n_73),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_35),
.B(n_27),
.C(n_30),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_24),
.B(n_21),
.C(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_66),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_34),
.B1(n_36),
.B2(n_32),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_71),
.B1(n_45),
.B2(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_32),
.B1(n_30),
.B2(n_34),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_67),
.B1(n_45),
.B2(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_28),
.B1(n_19),
.B2(n_22),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_15),
.B1(n_19),
.B2(n_14),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_62),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_44),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_24),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_48),
.C(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_71),
.C(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_68),
.B1(n_24),
.B2(n_14),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_45),
.B1(n_14),
.B2(n_23),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_71),
.B1(n_53),
.B2(n_45),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_57),
.B1(n_62),
.B2(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_58),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_81),
.C(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_106),
.B1(n_87),
.B2(n_83),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_111),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_113),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_70),
.B1(n_53),
.B2(n_45),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_114),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_55),
.B(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_26),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_76),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_21),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_76),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_113),
.B1(n_88),
.B2(n_92),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_130),
.C(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_86),
.C(n_96),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_114),
.C(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_139),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_118),
.B(n_120),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_13),
.B(n_10),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_105),
.B1(n_99),
.B2(n_97),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_138),
.B1(n_88),
.B2(n_1),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_99),
.B1(n_100),
.B2(n_86),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_21),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_125),
.B(n_126),
.C(n_130),
.D(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_151),
.B1(n_132),
.B2(n_134),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_14),
.C(n_23),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_149),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_23),
.B(n_2),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_133),
.B1(n_143),
.B2(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_158),
.Y(n_165)
);

NOR4xp25_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_133),
.C(n_143),
.D(n_136),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_146),
.C(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.C(n_8),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_144),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_163),
.A2(n_153),
.B(n_4),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_8),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_153),
.B(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_165),
.B1(n_10),
.B2(n_5),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_3),
.B(n_4),
.Y(n_174)
);

OAI311xp33_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_170),
.A3(n_171),
.B1(n_6),
.C1(n_7),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_173),
.B(n_5),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_4),
.Y(n_177)
);


endmodule