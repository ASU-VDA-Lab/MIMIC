module fake_aes_4434_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
AND2x4_ASAP7_75t_L g7 ( .A(n_2), .B(n_5), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_3), .Y(n_8) );
BUFx6f_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
NAND2xp33_ASAP7_75t_R g14 ( .A(n_11), .B(n_7), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_13), .B(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_SL g17 ( .A(n_16), .Y(n_17) );
O2A1O1Ixp33_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_14), .B(n_9), .C(n_2), .Y(n_18) );
OAI22x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_8), .B1(n_1), .B2(n_0), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
OAI22xp5_ASAP7_75t_SL g21 ( .A1(n_19), .A2(n_9), .B1(n_0), .B2(n_11), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_20), .B1(n_11), .B2(n_6), .Y(n_22) );
endmodule