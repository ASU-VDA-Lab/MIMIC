module fake_jpeg_11684_n_485 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_485);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_485;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_11),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_58),
.B(n_61),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_16),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_70),
.B(n_87),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_85),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_88),
.Y(n_119)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_48),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_14),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_98),
.Y(n_141)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_26),
.B1(n_30),
.B2(n_47),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_99),
.A2(n_131),
.B1(n_142),
.B2(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_102),
.B(n_105),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_109),
.B(n_110),
.Y(n_175)
);

NAND2x1p5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_30),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_113),
.B(n_68),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_50),
.B(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_116),
.B(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_81),
.B1(n_80),
.B2(n_88),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_82),
.B1(n_55),
.B2(n_66),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_77),
.A2(n_30),
.B1(n_47),
.B2(n_37),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_56),
.B(n_48),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_32),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_51),
.B(n_18),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_87),
.A2(n_47),
.B1(n_24),
.B2(n_37),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_59),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_46),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_144),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_52),
.B(n_46),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_43),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_43),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_155),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_27),
.B(n_33),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_157),
.A2(n_181),
.B(n_121),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_161),
.B1(n_163),
.B2(n_168),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_160),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_102),
.A2(n_57),
.B1(n_60),
.B2(n_23),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_97),
.B1(n_93),
.B2(n_86),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_164),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_166),
.A2(n_190),
.B(n_200),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_64),
.B1(n_25),
.B2(n_33),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_71),
.B1(n_32),
.B2(n_25),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_171),
.B(n_177),
.Y(n_244)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_44),
.B1(n_19),
.B2(n_45),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_178),
.A2(n_184),
.B1(n_198),
.B2(n_207),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_103),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_113),
.A2(n_83),
.B(n_71),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_120),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_201),
.Y(n_217)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_44),
.B1(n_19),
.B2(n_45),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_0),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_195),
.C(n_117),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_15),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_104),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_189),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_105),
.A2(n_15),
.A3(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_194),
.A2(n_137),
.B1(n_150),
.B2(n_127),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_141),
.B(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_126),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_204),
.B1(n_125),
.B2(n_151),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_208),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_130),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_112),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_205),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

BUFx24_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_125),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_124),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_128),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_127),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_210),
.A2(n_215),
.B(n_218),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_140),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_101),
.B1(n_150),
.B2(n_129),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_122),
.C(n_140),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_183),
.C(n_201),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_186),
.B1(n_163),
.B2(n_168),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_181),
.B(n_157),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_200),
.B(n_137),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_222),
.A2(n_223),
.B1(n_235),
.B2(n_164),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_159),
.A2(n_151),
.B1(n_149),
.B2(n_115),
.Y(n_223)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_230),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_155),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_124),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_199),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_114),
.B1(n_149),
.B2(n_115),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_158),
.A2(n_178),
.B1(n_175),
.B2(n_169),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_238),
.A2(n_241),
.B1(n_236),
.B2(n_222),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_107),
.B1(n_108),
.B2(n_114),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_147),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_250),
.B(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_165),
.B(n_122),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_252),
.B(n_210),
.C(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_258),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_165),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_211),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_277),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_213),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_263),
.B(n_269),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_218),
.A2(n_190),
.B1(n_167),
.B2(n_108),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_265),
.A2(n_285),
.B1(n_287),
.B2(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_225),
.A2(n_185),
.B1(n_156),
.B2(n_182),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_186),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_271),
.A2(n_292),
.B(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_206),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_272),
.B(n_273),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_205),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_173),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_280),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_225),
.A2(n_252),
.B(n_215),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_297),
.B(n_271),
.Y(n_316)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_217),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_249),
.B(n_176),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_156),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_284),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_193),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_209),
.A2(n_164),
.B1(n_192),
.B2(n_139),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_204),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_294),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_209),
.A2(n_106),
.B1(n_162),
.B2(n_203),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_106),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_295),
.B1(n_226),
.B2(n_248),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_11),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_236),
.A2(n_11),
.B1(n_12),
.B2(n_238),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_227),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_234),
.A2(n_252),
.B(n_245),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_237),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_259),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_322),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_223),
.B1(n_235),
.B2(n_216),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_324),
.B1(n_326),
.B2(n_287),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_256),
.A2(n_234),
.B1(n_241),
.B2(n_248),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_282),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_315),
.B(n_320),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_329),
.B(n_275),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_214),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_319),
.B(n_335),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_259),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_240),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_295),
.A2(n_226),
.B1(n_254),
.B2(n_251),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_240),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_337),
.Y(n_345)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_256),
.A2(n_246),
.B(n_237),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_220),
.C(n_232),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_332),
.C(n_283),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_262),
.B(n_232),
.C(n_242),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_242),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_336),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_258),
.B(n_251),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_212),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_260),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_314),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_348),
.Y(n_371)
);

XOR2x1_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_297),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_306),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_342),
.A2(n_353),
.B(n_361),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g346 ( 
.A(n_310),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_346),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_314),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_328),
.Y(n_349)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_349),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_301),
.A2(n_264),
.B1(n_265),
.B2(n_291),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_354),
.A2(n_359),
.B1(n_367),
.B2(n_325),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_364),
.C(n_366),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_357),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_296),
.Y(n_358)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_302),
.A2(n_288),
.B1(n_285),
.B2(n_296),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_263),
.B1(n_272),
.B2(n_269),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_360),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_266),
.B(n_294),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_323),
.B(n_329),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_309),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_368),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_266),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_273),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_318),
.A2(n_281),
.B1(n_277),
.B2(n_284),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_280),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_308),
.Y(n_374)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_374),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_362),
.A2(n_326),
.B1(n_300),
.B2(n_301),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_390),
.B1(n_392),
.B2(n_353),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_379),
.A2(n_395),
.B1(n_343),
.B2(n_344),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_331),
.C(n_319),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_389),
.C(n_391),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_338),
.B(n_317),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_386),
.B(n_367),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_317),
.Y(n_388)
);

NAND2xp33_ASAP7_75t_SL g412 ( 
.A(n_388),
.B(n_394),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_366),
.C(n_356),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_362),
.A2(n_308),
.B1(n_323),
.B2(n_330),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_335),
.C(n_313),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_339),
.A2(n_308),
.B1(n_311),
.B2(n_333),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_311),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_354),
.A2(n_303),
.B1(n_304),
.B2(n_268),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_340),
.B(n_307),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_363),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_341),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_398),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_349),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_347),
.C(n_365),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_399),
.B(n_381),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_345),
.C(n_339),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_414),
.C(n_373),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_415),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_361),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_405),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_345),
.Y(n_405)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_382),
.A2(n_359),
.B1(n_343),
.B2(n_344),
.Y(n_409)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_411),
.A2(n_419),
.B1(n_374),
.B2(n_387),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_358),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_416),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_386),
.C(n_382),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_390),
.B(n_368),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_379),
.A2(n_352),
.B1(n_350),
.B2(n_346),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_375),
.B1(n_392),
.B2(n_393),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_373),
.B(n_342),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_385),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_395),
.A2(n_350),
.B1(n_307),
.B2(n_310),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_436),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_393),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_426),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_394),
.B1(n_396),
.B2(n_370),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_372),
.C(n_383),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_387),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_419),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_387),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_429),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_430),
.A2(n_401),
.B1(n_414),
.B2(n_407),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_406),
.B(n_371),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_437),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_434),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_372),
.C(n_383),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_397),
.C(n_400),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_400),
.B(n_388),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_440),
.Y(n_457)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_435),
.C(n_422),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_418),
.C(n_416),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_444),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_426),
.C(n_420),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_431),
.A2(n_370),
.B1(n_412),
.B2(n_415),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_430),
.B1(n_436),
.B2(n_433),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_428),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_377),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_428),
.A2(n_413),
.B(n_377),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_423),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_441),
.B(n_427),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_458),
.Y(n_469)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_463),
.C(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_448),
.B(n_420),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_459),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_423),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_461),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_433),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_447),
.B(n_305),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_462),
.A2(n_384),
.B(n_292),
.Y(n_466)
);

AOI322xp5_ASAP7_75t_L g464 ( 
.A1(n_455),
.A2(n_446),
.A3(n_438),
.B1(n_440),
.B2(n_439),
.C1(n_443),
.C2(n_451),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_465),
.Y(n_474)
);

AOI322xp5_ASAP7_75t_L g465 ( 
.A1(n_457),
.A2(n_449),
.A3(n_442),
.B1(n_444),
.B2(n_384),
.C1(n_305),
.C2(n_278),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_472),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_457),
.A2(n_384),
.B1(n_276),
.B2(n_270),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_467),
.A2(n_276),
.B1(n_463),
.B2(n_454),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_473),
.A2(n_470),
.B1(n_469),
.B2(n_467),
.Y(n_478)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_471),
.A2(n_460),
.B1(n_453),
.B2(n_246),
.C(n_292),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_476),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_292),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_477),
.B(n_470),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_475),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_474),
.B(n_476),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_482),
.Y(n_483)
);

AO22x1_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_480),
.B1(n_246),
.B2(n_212),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_254),
.Y(n_485)
);


endmodule