module fake_ariane_1022_n_2076 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2076);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2076;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_279;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_212;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1865;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_23),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_65),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_115),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_166),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_85),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_14),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_9),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_111),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_8),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_41),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_125),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_140),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_63),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_135),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_91),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_202),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_82),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_100),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_112),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_198),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_156),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_151),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_81),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_7),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_147),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_74),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_189),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_57),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_116),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_65),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_103),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_171),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_37),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_50),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_34),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_44),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_144),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_96),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_59),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_141),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_150),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_131),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_83),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_94),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_15),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_186),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_45),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_181),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_39),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_95),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_184),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_64),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_93),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_87),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_163),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_92),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_172),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_137),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_108),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_109),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_27),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_107),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_152),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_160),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_76),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_178),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_6),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_2),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_50),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_170),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_3),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_25),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_16),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_72),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_53),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_130),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_12),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_22),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_51),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_99),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_36),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_2),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_12),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_5),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_32),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_180),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_192),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_0),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_58),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_70),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_173),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_29),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_59),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_127),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_38),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_15),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_113),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_86),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_196),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_30),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_40),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_124),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_132),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_168),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_201),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_75),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_60),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_73),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_89),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_20),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_48),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_11),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_52),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_183),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_187),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_57),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_29),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_190),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_197),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_118),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_139),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_193),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_55),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_51),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_97),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_78),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_102),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_161),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_10),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_46),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_129),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_199),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_27),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_30),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_128),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_8),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_121),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_16),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_157),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_142),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_73),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_20),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_19),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_88),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_1),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_154),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_105),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_33),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_33),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_79),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_47),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_38),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_44),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_138),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_11),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_10),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_110),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_67),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_167),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_63),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_74),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_136),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_90),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_101),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_98),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_194),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_4),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_48),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_34),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_203),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_224),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_229),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_203),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_204),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_224),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_211),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_204),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_213),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_284),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_213),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_214),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_275),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_214),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_342),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_306),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_209),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_219),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_275),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_365),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_306),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_400),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_262),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_375),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_219),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_294),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_225),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_215),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_225),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_230),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_208),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_327),
.B(n_1),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_208),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_230),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_234),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_227),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_327),
.B(n_3),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_227),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_234),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_281),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_281),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_301),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_334),
.B(n_5),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_317),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_238),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_354),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_264),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_238),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_215),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_239),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_301),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_264),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_283),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_210),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_323),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_239),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_241),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_386),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_220),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_249),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_283),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_381),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_323),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_249),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_366),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_270),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_226),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_270),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_381),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_286),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_231),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_334),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_233),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_286),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_237),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_251),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_296),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_261),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_288),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_265),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_337),
.B(n_6),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_288),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_228),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_274),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_303),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_303),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_276),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_314),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_314),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_228),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_339),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_339),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_355),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_228),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_282),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_287),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_355),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_357),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_228),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_240),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_298),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_302),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_465),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_407),
.B(n_357),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_407),
.B(n_218),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_410),
.B(n_241),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_430),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_417),
.B(n_241),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_418),
.B(n_362),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_424),
.B(n_218),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

CKINVDCx8_ASAP7_75t_R g537 ( 
.A(n_436),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_432),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_432),
.A2(n_290),
.B(n_216),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_435),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_438),
.B(n_258),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_438),
.B(n_241),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_511),
.B(n_241),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_443),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_453),
.B(n_258),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_453),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_458),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_464),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_408),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_482),
.A2(n_206),
.B1(n_223),
.B2(n_222),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_464),
.A2(n_368),
.B(n_362),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_489),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_511),
.B(n_241),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_472),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_472),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_475),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_477),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_480),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_436),
.B(n_361),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_484),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_493),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_490),
.B(n_368),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_493),
.B(n_374),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_496),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_496),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_497),
.B(n_278),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_441),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_440),
.B(n_240),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_445),
.B(n_451),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_500),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_500),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_423),
.B(n_240),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_503),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_562),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_525),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_562),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_562),
.B(n_580),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_576),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_562),
.B(n_580),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_528),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_528),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_523),
.B(n_433),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_552),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_550),
.B(n_457),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_544),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_523),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_548),
.B(n_566),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_552),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_552),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_528),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_580),
.B(n_423),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_580),
.B(n_374),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_525),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_544),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_590),
.B(n_467),
.C(n_462),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_595),
.B(n_457),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_552),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_552),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_552),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_595),
.B(n_548),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_552),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_525),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_552),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_550),
.B(n_461),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_461),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_577),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_544),
.B(n_408),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_525),
.B(n_232),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_525),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_525),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_577),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_544),
.B(n_408),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_544),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_590),
.A2(n_422),
.B1(n_434),
.B2(n_428),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_576),
.B(n_476),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_537),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_576),
.B(n_481),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_530),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_577),
.Y(n_650)
);

INVx4_ASAP7_75t_SL g651 ( 
.A(n_525),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_533),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_577),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_576),
.B(n_483),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_577),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_527),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_544),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_589),
.A2(n_434),
.B1(n_431),
.B2(n_492),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_589),
.A2(n_487),
.B1(n_491),
.B2(n_485),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_564),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_558),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_577),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_565),
.B(n_495),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_558),
.B(n_412),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_558),
.B(n_412),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_SL g668 ( 
.A1(n_537),
.A2(n_446),
.B1(n_450),
.B2(n_449),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_564),
.A2(n_431),
.B1(n_504),
.B2(n_503),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_577),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_565),
.B(n_498),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_527),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_526),
.B(n_459),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_577),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_537),
.B(n_506),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_537),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_527),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_533),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_519),
.B(n_394),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_527),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_564),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_526),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_558),
.B(n_419),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_527),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_598),
.B(n_507),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_527),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_598),
.B(n_513),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_542),
.B(n_409),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_527),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_542),
.B(n_494),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_564),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_542),
.B(n_512),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_527),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_519),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_536),
.B(n_509),
.C(n_508),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_563),
.B(n_361),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_519),
.B(n_394),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_527),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_547),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_547),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_564),
.A2(n_505),
.B1(n_510),
.B2(n_501),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_547),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_536),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_547),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_572),
.B(n_419),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_541),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_547),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_564),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_547),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_572),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_588),
.B(n_416),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_541),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_554),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_563),
.A2(n_469),
.B1(n_478),
.B2(n_470),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_554),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_SL g721 ( 
.A(n_588),
.B(n_277),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_554),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_572),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_588),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_519),
.B(n_529),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_572),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_563),
.A2(n_330),
.B1(n_460),
.B2(n_455),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_518),
.A2(n_545),
.B1(n_555),
.B2(n_535),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_519),
.B(n_399),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_518),
.A2(n_425),
.B1(n_488),
.B2(n_419),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_554),
.Y(n_731)
);

INVx4_ASAP7_75t_SL g732 ( 
.A(n_554),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_598),
.B(n_425),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_554),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_554),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_592),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_554),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_592),
.A2(n_471),
.B1(n_473),
.B2(n_463),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_572),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_591),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_591),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_488),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_591),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_592),
.B(n_421),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_518),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_518),
.B(n_479),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_605),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_602),
.A2(n_574),
.B(n_551),
.C(n_556),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_627),
.B(n_574),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

INVxp33_ASAP7_75t_L g752 ( 
.A(n_607),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_686),
.B(n_574),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_699),
.A2(n_618),
.B1(n_662),
.B2(n_612),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_618),
.A2(n_551),
.B1(n_556),
.B2(n_549),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_616),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_646),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_609),
.B(n_426),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_632),
.B(n_574),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_648),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_649),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_603),
.B(n_574),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_574),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_689),
.B(n_549),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_699),
.B(n_535),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_662),
.B(n_591),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_SL g767 ( 
.A(n_645),
.B(n_427),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_699),
.A2(n_520),
.B1(n_522),
.B2(n_521),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_652),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_670),
.B(n_549),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_609),
.B(n_429),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_662),
.B(n_591),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_610),
.B(n_642),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_746),
.B(n_551),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_747),
.B(n_556),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_618),
.A2(n_559),
.B1(n_567),
.B2(n_557),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_669),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_747),
.B(n_557),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_747),
.B(n_557),
.Y(n_779)
);

BUFx8_ASAP7_75t_L g780 ( 
.A(n_724),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_679),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_623),
.B(n_559),
.Y(n_782)
);

XOR2xp5_ASAP7_75t_L g783 ( 
.A(n_607),
.B(n_413),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_617),
.B(n_559),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_725),
.B(n_567),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_725),
.B(n_567),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_620),
.B(n_568),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_604),
.A2(n_569),
.B(n_570),
.C(n_568),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_610),
.B(n_591),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_724),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_687),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_610),
.B(n_591),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_611),
.Y(n_793)
);

INVx8_ASAP7_75t_L g794 ( 
.A(n_618),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_699),
.A2(n_454),
.B1(n_466),
.B2(n_452),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_611),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_708),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_715),
.B(n_568),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_643),
.B(n_570),
.C(n_569),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_721),
.B(n_222),
.C(n_206),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_618),
.B(n_569),
.Y(n_801)
);

INVxp33_ASAP7_75t_L g802 ( 
.A(n_674),
.Y(n_802)
);

OR2x2_ASAP7_75t_SL g803 ( 
.A(n_716),
.B(n_474),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_642),
.B(n_591),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_682),
.A2(n_539),
.B(n_570),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_618),
.B(n_612),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_612),
.A2(n_520),
.B1(n_522),
.B2(n_521),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_683),
.B(n_486),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_612),
.A2(n_578),
.B1(n_579),
.B2(n_573),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_733),
.B(n_573),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_743),
.B(n_573),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_711),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_717),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_721),
.A2(n_579),
.B1(n_583),
.B2(n_578),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_730),
.B(n_578),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_642),
.B(n_579),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_727),
.A2(n_520),
.B1(n_522),
.B2(n_521),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_583),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_SL g819 ( 
.A(n_645),
.B(n_240),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_663),
.B(n_583),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_680),
.A2(n_593),
.B1(n_594),
.B2(n_586),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_680),
.A2(n_729),
.B1(n_700),
.B2(n_693),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_723),
.B(n_591),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_723),
.B(n_586),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_678),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_599),
.A2(n_539),
.B(n_531),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_716),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_680),
.A2(n_594),
.B1(n_593),
.B2(n_545),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_726),
.B(n_593),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_745),
.Y(n_831)
);

BUFx6f_ASAP7_75t_SL g832 ( 
.A(n_680),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_726),
.B(n_594),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_659),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_728),
.B(n_659),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_697),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_739),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_739),
.B(n_520),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_677),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_601),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_661),
.B(n_517),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_682),
.A2(n_693),
.B(n_713),
.C(n_698),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_702),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_745),
.B(n_535),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_634),
.B(n_641),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_622),
.B(n_517),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_666),
.B(n_522),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_713),
.B(n_524),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_680),
.A2(n_700),
.B1(n_729),
.B2(n_660),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_674),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_734),
.B(n_524),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_667),
.B(n_524),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_684),
.B(n_532),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_710),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_680),
.A2(n_545),
.B1(n_555),
.B2(n_535),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_532),
.Y(n_856)
);

BUFx5_ASAP7_75t_L g857 ( 
.A(n_600),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_692),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_734),
.B(n_532),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_736),
.B(n_545),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_700),
.B(n_534),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_734),
.B(n_534),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_644),
.B(n_517),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_696),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_736),
.B(n_555),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_647),
.B(n_531),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_631),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_696),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_700),
.B(n_534),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_654),
.B(n_676),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_738),
.B(n_531),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_700),
.B(n_729),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_734),
.B(n_534),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_729),
.A2(n_540),
.B1(n_543),
.B2(n_538),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_734),
.B(n_538),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_696),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_729),
.B(n_538),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_729),
.A2(n_585),
.B1(n_555),
.B2(n_582),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_631),
.B(n_585),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_601),
.B(n_538),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_705),
.A2(n_543),
.B1(n_553),
.B2(n_540),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_694),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_665),
.B(n_540),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_703),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_672),
.A2(n_585),
.B1(n_582),
.B2(n_581),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_677),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_628),
.B(n_540),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_628),
.B(n_543),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_L g889 ( 
.A(n_628),
.B(n_543),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_668),
.B(n_209),
.Y(n_890)
);

NAND2x1_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_553),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_695),
.B(n_553),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_703),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_628),
.B(n_553),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_719),
.B(n_585),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_695),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_704),
.B(n_581),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_L g898 ( 
.A(n_690),
.B(n_246),
.C(n_223),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_704),
.B(n_488),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_704),
.B(n_560),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_706),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_706),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_600),
.A2(n_582),
.B(n_581),
.C(n_561),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_628),
.B(n_650),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_722),
.B(n_560),
.Y(n_905)
);

NAND2x1_ASAP7_75t_L g906 ( 
.A(n_722),
.B(n_560),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_737),
.B(n_561),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_737),
.B(n_561),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_619),
.A2(n_575),
.B(n_584),
.C(n_571),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_840),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_759),
.B(n_650),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_871),
.B(n_571),
.Y(n_912)
);

AO21x1_ASAP7_75t_L g913 ( 
.A1(n_759),
.A2(n_401),
.B(n_399),
.Y(n_913)
);

AND2x2_ASAP7_75t_SL g914 ( 
.A(n_754),
.B(n_401),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_871),
.B(n_863),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_790),
.B(n_630),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_794),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_846),
.A2(n_571),
.B(n_584),
.C(n_575),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_757),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_863),
.B(n_630),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_866),
.B(n_575),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_785),
.B(n_650),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_793),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_846),
.A2(n_709),
.B(n_712),
.C(n_707),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_840),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_794),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_827),
.A2(n_636),
.B(n_629),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_764),
.A2(n_584),
.B(n_587),
.C(n_575),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_848),
.A2(n_637),
.B(n_636),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_866),
.B(n_630),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_765),
.B(n_651),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_786),
.B(n_650),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_885),
.B(n_584),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_754),
.A2(n_639),
.B1(n_655),
.B2(n_637),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_773),
.A2(n_655),
.B(n_639),
.Y(n_935)
);

NOR2x1_ASAP7_75t_L g936 ( 
.A(n_839),
.B(n_587),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_780),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_773),
.A2(n_673),
.B(n_658),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_841),
.B(n_587),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_845),
.A2(n_673),
.B(n_658),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_766),
.A2(n_685),
.B(n_681),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_824),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_772),
.A2(n_691),
.B(n_688),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_822),
.B(n_650),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_772),
.A2(n_731),
.B(n_701),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_860),
.B(n_587),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_750),
.A2(n_731),
.B(n_701),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_904),
.A2(n_742),
.B(n_740),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_762),
.B(n_763),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_844),
.B(n_640),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_762),
.A2(n_597),
.B(n_596),
.C(n_250),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_849),
.A2(n_742),
.B1(n_740),
.B2(n_709),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_763),
.B(n_596),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_774),
.B(n_596),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_782),
.B(n_596),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_782),
.B(n_597),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_L g957 ( 
.A(n_828),
.B(n_250),
.C(n_246),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_775),
.B(n_597),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_822),
.B(n_664),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_778),
.B(n_597),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_904),
.A2(n_712),
.B(n_707),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_779),
.B(n_519),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_816),
.A2(n_718),
.B(n_714),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_844),
.B(n_640),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_818),
.A2(n_825),
.B(n_820),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_878),
.B(n_529),
.Y(n_966)
);

INVx11_ASAP7_75t_L g967 ( 
.A(n_780),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_784),
.A2(n_256),
.B(n_263),
.C(n_254),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_805),
.A2(n_842),
.B(n_897),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_809),
.A2(n_539),
.B(n_546),
.C(n_529),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_768),
.B(n_529),
.Y(n_971)
);

AND2x2_ASAP7_75t_SL g972 ( 
.A(n_849),
.B(n_364),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_897),
.A2(n_735),
.B(n_720),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_794),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_865),
.B(n_529),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_835),
.A2(n_903),
.B(n_870),
.C(n_799),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_892),
.A2(n_905),
.B(n_900),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_753),
.A2(n_256),
.B(n_263),
.C(n_254),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_768),
.B(n_529),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_755),
.A2(n_671),
.B1(n_640),
.B2(n_720),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_831),
.A2(n_300),
.B(n_304),
.C(n_268),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_844),
.B(n_882),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_907),
.A2(n_741),
.B(n_735),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_757),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_908),
.A2(n_744),
.B(n_741),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_855),
.B(n_546),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_814),
.B(n_546),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_870),
.A2(n_744),
.B1(n_671),
.B2(n_608),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_760),
.B(n_546),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_761),
.B(n_546),
.Y(n_990)
);

AO21x1_ASAP7_75t_L g991 ( 
.A1(n_810),
.A2(n_811),
.B(n_851),
.Y(n_991)
);

NOR2x1_ASAP7_75t_R g992 ( 
.A(n_886),
.B(n_305),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_847),
.A2(n_614),
.B(n_613),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_800),
.A2(n_546),
.B(n_300),
.C(n_304),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_796),
.B(n_268),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_852),
.A2(n_615),
.B(n_614),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_826),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_776),
.A2(n_671),
.B1(n_624),
.B2(n_625),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_843),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_777),
.B(n_621),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_781),
.B(n_797),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_853),
.A2(n_625),
.B(n_624),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_812),
.B(n_626),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_813),
.B(n_633),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_895),
.B(n_638),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_807),
.B(n_638),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_748),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_789),
.A2(n_657),
.B(n_653),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_832),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_807),
.B(n_653),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_751),
.B(n_657),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_789),
.A2(n_675),
.B(n_664),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_756),
.B(n_769),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_791),
.B(n_675),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_SL g1015 ( 
.A(n_767),
.B(n_839),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_819),
.B(n_664),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_902),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_792),
.A2(n_823),
.B(n_804),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_808),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_896),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_867),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_792),
.A2(n_823),
.B(n_804),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_851),
.A2(n_515),
.B(n_514),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_896),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_850),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_806),
.B(n_664),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_788),
.A2(n_318),
.B(n_380),
.C(n_328),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_864),
.B(n_664),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_868),
.B(n_651),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_829),
.B(n_876),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_857),
.B(n_651),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_883),
.B(n_651),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_787),
.B(n_732),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_802),
.B(n_307),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_830),
.A2(n_656),
.B(n_635),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_758),
.B(n_318),
.C(n_312),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_798),
.B(n_732),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_771),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_899),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_879),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_817),
.A2(n_328),
.B(n_332),
.C(n_345),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_858),
.B(n_765),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_817),
.B(n_732),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_838),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_854),
.B(n_732),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_830),
.A2(n_656),
.B(n_322),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_834),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_765),
.B(n_209),
.Y(n_1048)
);

NOR2x1p5_ASAP7_75t_L g1049 ( 
.A(n_803),
.B(n_872),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_891),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_881),
.B(n_312),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_832),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_833),
.A2(n_909),
.B(n_749),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_836),
.B(n_308),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_884),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_898),
.B(n_332),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_833),
.A2(n_656),
.B(n_207),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_783),
.B(n_209),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_887),
.A2(n_656),
.B(n_212),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_770),
.A2(n_345),
.B1(n_347),
.B2(n_349),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_859),
.A2(n_372),
.B(n_364),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_887),
.A2(n_217),
.B(n_205),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_837),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_857),
.B(n_821),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_881),
.B(n_347),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_894),
.A2(n_515),
.B(n_514),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_856),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_L g1068 ( 
.A(n_795),
.B(n_350),
.C(n_349),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_874),
.B(n_350),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_890),
.B(n_309),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_801),
.A2(n_311),
.B1(n_333),
.B2(n_329),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_894),
.A2(n_235),
.B(n_221),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_874),
.B(n_815),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_752),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_861),
.B(n_360),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_859),
.A2(n_873),
.B(n_862),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_869),
.B(n_360),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_862),
.A2(n_244),
.B(n_242),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_877),
.B(n_367),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_893),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_901),
.B(n_367),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_880),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_857),
.B(n_391),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_873),
.A2(n_247),
.B(n_245),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_875),
.A2(n_252),
.B(n_248),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_875),
.A2(n_257),
.B(n_255),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_906),
.B(n_370),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_857),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_915),
.A2(n_889),
.B(n_888),
.C(n_391),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_912),
.B(n_857),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1013),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_925),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_857),
.B(n_377),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1007),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_931),
.B(n_370),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_920),
.B(n_516),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_972),
.A2(n_380),
.B1(n_388),
.B2(n_405),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_972),
.A2(n_397),
.B1(n_388),
.B2(n_405),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1015),
.B(n_313),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_965),
.A2(n_969),
.B(n_977),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1064),
.A2(n_377),
.B(n_372),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1038),
.B(n_315),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_925),
.Y(n_1103)
);

CKINVDCx6p67_ASAP7_75t_R g1104 ( 
.A(n_923),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1021),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_925),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_920),
.B(n_516),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_917),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1036),
.A2(n_378),
.B(n_382),
.C(n_397),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1064),
.A2(n_243),
.B(n_236),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_921),
.A2(n_930),
.B(n_911),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_982),
.A2(n_379),
.B1(n_406),
.B2(n_344),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_967),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_930),
.A2(n_911),
.B(n_940),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_SL g1115 ( 
.A(n_1070),
.B(n_319),
.C(n_316),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_982),
.B(n_320),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_937),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1040),
.B(n_324),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1025),
.B(n_325),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_R g1120 ( 
.A(n_1009),
.B(n_326),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_919),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_925),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1021),
.B(n_338),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1074),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_927),
.A2(n_253),
.B(n_321),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1019),
.B(n_378),
.Y(n_1126)
);

NOR2xp67_ASAP7_75t_L g1127 ( 
.A(n_1009),
.B(n_516),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_931),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_953),
.A2(n_947),
.B(n_993),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_216),
.B(n_290),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1070),
.B(n_343),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_941),
.A2(n_516),
.B(n_216),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1052),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1034),
.B(n_348),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_914),
.A2(n_390),
.B1(n_373),
.B2(n_398),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_914),
.A2(n_389),
.B1(n_382),
.B2(n_393),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_946),
.B(n_353),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_917),
.B(n_371),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1058),
.B(n_385),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_984),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1052),
.B(n_389),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_976),
.B(n_393),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1001),
.A2(n_278),
.B1(n_293),
.B2(n_395),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1034),
.B(n_392),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1080),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_910),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_950),
.Y(n_1147)
);

INVxp67_ASAP7_75t_SL g1148 ( 
.A(n_1005),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_975),
.B(n_1042),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1042),
.B(n_259),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1055),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_950),
.B(n_260),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1060),
.A2(n_403),
.B1(n_266),
.B2(n_387),
.Y(n_1153)
);

OAI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_1054),
.A2(n_296),
.B(n_216),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1068),
.A2(n_290),
.B1(n_384),
.B2(n_383),
.C(n_376),
.Y(n_1155)
);

AO21x1_ASAP7_75t_L g1156 ( 
.A1(n_1083),
.A2(n_290),
.B(n_402),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_926),
.B(n_267),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1060),
.B(n_9),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1055),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1041),
.A2(n_310),
.B1(n_369),
.B2(n_363),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1073),
.B(n_17),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_926),
.B(n_269),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_964),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1049),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1027),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1048),
.B(n_18),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1044),
.B(n_21),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1081),
.B(n_21),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_SL g1169 ( 
.A1(n_1053),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1027),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_SL g1171 ( 
.A1(n_1083),
.A2(n_402),
.B(n_232),
.C(n_358),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_992),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1082),
.B(n_28),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_995),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_957),
.B(n_31),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1030),
.A2(n_32),
.B(n_35),
.C(n_36),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_964),
.B(n_1041),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_955),
.B(n_35),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_956),
.B(n_37),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1047),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_958),
.B(n_40),
.Y(n_1181)
);

CKINVDCx8_ASAP7_75t_R g1182 ( 
.A(n_1056),
.Y(n_1182)
);

OAI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_986),
.A2(n_299),
.B1(n_359),
.B2(n_356),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1030),
.A2(n_297),
.B1(n_352),
.B2(n_351),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_910),
.B(n_271),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1054),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1039),
.B(n_42),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_L g1188 ( 
.A(n_978),
.B(n_295),
.C(n_346),
.Y(n_1188)
);

INVxp33_ASAP7_75t_SL g1189 ( 
.A(n_1071),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1056),
.B(n_962),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1069),
.A2(n_292),
.B1(n_341),
.B2(n_340),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_968),
.A2(n_913),
.B(n_1051),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1065),
.A2(n_966),
.B1(n_1067),
.B2(n_971),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_999),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_916),
.A2(n_289),
.B1(n_336),
.B2(n_335),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1002),
.A2(n_285),
.B(n_331),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_916),
.B(n_280),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1016),
.B(n_279),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1020),
.B(n_272),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_942),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_960),
.A2(n_990),
.B1(n_989),
.B2(n_970),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1087),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_954),
.B(n_979),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_970),
.A2(n_987),
.B1(n_994),
.B2(n_933),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1075),
.B(n_43),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_963),
.A2(n_291),
.B(n_273),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1077),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_944),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_951),
.A2(n_402),
.B(n_232),
.C(n_47),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_974),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_973),
.A2(n_402),
.B(n_232),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1079),
.B(n_43),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1050),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_997),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_994),
.B(n_46),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1017),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_983),
.A2(n_84),
.B(n_188),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1020),
.B(n_49),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_985),
.A2(n_961),
.B(n_1012),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_944),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_918),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1017),
.Y(n_1222)
);

AO32x2_ASAP7_75t_L g1223 ( 
.A1(n_934),
.A2(n_56),
.A3(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1024),
.B(n_61),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_981),
.A2(n_918),
.B(n_928),
.C(n_932),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1063),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1024),
.B(n_66),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1050),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_922),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1063),
.B(n_69),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_936),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_924),
.A2(n_126),
.B(n_182),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_939),
.B(n_70),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1018),
.A2(n_71),
.B(n_75),
.C(n_76),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1006),
.B(n_71),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1000),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1132),
.A2(n_1076),
.B(n_945),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1111),
.A2(n_1022),
.B(n_952),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_L g1239 ( 
.A1(n_1134),
.A2(n_1004),
.B(n_1003),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1100),
.A2(n_991),
.A3(n_1061),
.B(n_1045),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1156),
.A2(n_1043),
.A3(n_1032),
.B(n_1037),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1211),
.A2(n_1026),
.B(n_922),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1131),
.A2(n_932),
.B(n_959),
.C(n_1046),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1090),
.A2(n_1088),
.B(n_1031),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1094),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1144),
.A2(n_1028),
.B(n_959),
.C(n_1026),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1090),
.A2(n_1129),
.B(n_1201),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1201),
.A2(n_1088),
.B(n_1031),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1180),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_1033),
.A3(n_1010),
.B(n_943),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1186),
.B(n_1011),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1219),
.A2(n_1093),
.B(n_1096),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1136),
.A2(n_988),
.B1(n_980),
.B2(n_998),
.Y(n_1253)
);

OAI22x1_ASAP7_75t_L g1254 ( 
.A1(n_1135),
.A2(n_1023),
.B1(n_1014),
.B2(n_1029),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1096),
.A2(n_935),
.B(n_938),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1174),
.B(n_1072),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1232),
.A2(n_948),
.B(n_1008),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1105),
.B(n_1066),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1204),
.A2(n_1059),
.A3(n_1057),
.B(n_1062),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1207),
.B(n_1086),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1130),
.A2(n_929),
.B(n_1035),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1097),
.A2(n_1050),
.B(n_1084),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1217),
.A2(n_974),
.B(n_1078),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1142),
.A2(n_1085),
.B(n_1050),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1189),
.A2(n_77),
.B(n_80),
.C(n_114),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1202),
.B(n_77),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1107),
.A2(n_119),
.B(n_122),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1091),
.B(n_200),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1107),
.A2(n_123),
.B(n_133),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1204),
.A2(n_134),
.A3(n_143),
.B(n_149),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1115),
.A2(n_153),
.B(n_155),
.C(n_164),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1104),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1147),
.B(n_175),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1125),
.A2(n_177),
.B(n_1191),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1136),
.A2(n_1097),
.B1(n_1098),
.B2(n_1158),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1128),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1171),
.A2(n_1101),
.B(n_1225),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1191),
.A2(n_1142),
.B(n_1161),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1203),
.A2(n_1178),
.B(n_1179),
.Y(n_1279)
);

AOI221x1_ASAP7_75t_L g1280 ( 
.A1(n_1221),
.A2(n_1098),
.B1(n_1234),
.B2(n_1154),
.C(n_1192),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1203),
.A2(n_1178),
.B(n_1179),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1163),
.B(n_1139),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1109),
.A2(n_1192),
.B(n_1212),
.C(n_1205),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1181),
.A2(n_1161),
.B(n_1089),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1181),
.A2(n_1235),
.B(n_1197),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1118),
.B(n_1095),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1113),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1208),
.A2(n_1218),
.B(n_1227),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1124),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1152),
.A2(n_1116),
.B(n_1160),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1150),
.B(n_1182),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_SL g1292 ( 
.A1(n_1169),
.A2(n_1209),
.B(n_1221),
.C(n_1162),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1165),
.A2(n_1170),
.B(n_1176),
.C(n_1175),
.Y(n_1293)
);

NOR4xp25_ASAP7_75t_L g1294 ( 
.A(n_1229),
.B(n_1215),
.C(n_1143),
.D(n_1177),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1172),
.Y(n_1295)
);

AOI221x1_ASAP7_75t_L g1296 ( 
.A1(n_1143),
.A2(n_1160),
.B1(n_1230),
.B2(n_1224),
.C(n_1110),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1149),
.B(n_1099),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1190),
.B(n_1146),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1095),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1220),
.A2(n_1112),
.B1(n_1168),
.B2(n_1164),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1236),
.A2(n_1173),
.B(n_1167),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1128),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1145),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1146),
.B(n_1193),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1120),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1167),
.A2(n_1173),
.B(n_1148),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1233),
.A2(n_1188),
.B(n_1187),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1155),
.A2(n_1199),
.B(n_1184),
.C(n_1166),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1214),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1151),
.A2(n_1159),
.B(n_1140),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1126),
.B(n_1137),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1198),
.A2(n_1185),
.B(n_1206),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1121),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_SL g1314 ( 
.A(n_1226),
.B(n_1195),
.C(n_1102),
.Y(n_1314)
);

AO32x2_ASAP7_75t_L g1315 ( 
.A1(n_1223),
.A2(n_1153),
.A3(n_1231),
.B1(n_1210),
.B2(n_1216),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1141),
.B(n_1128),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1123),
.B(n_1117),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1196),
.A2(n_1108),
.B(n_1213),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1183),
.A2(n_1127),
.B(n_1222),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1141),
.A2(n_1223),
.B(n_1119),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_L g1321 ( 
.A(n_1157),
.B(n_1138),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1194),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1223),
.A2(n_1213),
.A3(n_1103),
.B(n_1106),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1133),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_1133),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1146),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1108),
.A2(n_1228),
.B1(n_1213),
.B2(n_1106),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1108),
.A2(n_1092),
.B(n_1103),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1108),
.A2(n_1092),
.B(n_1103),
.Y(n_1329)
);

NAND2xp33_ASAP7_75t_L g1330 ( 
.A(n_1092),
.B(n_1106),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1122),
.A2(n_915),
.B(n_1131),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1133),
.B(n_1122),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1122),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1094),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1134),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1132),
.A2(n_1219),
.B(n_1129),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1186),
.B(n_915),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1094),
.Y(n_1338)
);

OAI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1134),
.A2(n_915),
.B(n_1144),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1186),
.A2(n_915),
.B1(n_1189),
.B2(n_1144),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1174),
.B(n_844),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1105),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1134),
.A2(n_915),
.B(n_1144),
.C(n_1131),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1094),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1113),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1094),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1128),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1144),
.C(n_1134),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1111),
.A2(n_915),
.B(n_976),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1094),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1100),
.A2(n_991),
.A3(n_1061),
.B(n_1156),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1186),
.B(n_915),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1128),
.B(n_931),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1105),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1134),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1132),
.A2(n_1219),
.B(n_1129),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1134),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1134),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1200),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1094),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1124),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1100),
.A2(n_991),
.A3(n_1061),
.B(n_1156),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1131),
.A2(n_915),
.B1(n_1136),
.B2(n_1098),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1113),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1186),
.A2(n_915),
.B1(n_1189),
.B2(n_1144),
.Y(n_1368)
);

NAND2x2_ASAP7_75t_L g1369 ( 
.A(n_1117),
.B(n_937),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_L g1370 ( 
.A1(n_1131),
.A2(n_1144),
.B(n_1134),
.C(n_915),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1186),
.B(n_915),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1111),
.A2(n_915),
.B(n_976),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1139),
.B(n_844),
.Y(n_1373)
);

AOI221x1_ASAP7_75t_L g1374 ( 
.A1(n_1221),
.A2(n_1098),
.B1(n_1097),
.B2(n_1136),
.C(n_915),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1108),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1104),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1186),
.B(n_915),
.Y(n_1377)
);

BUFx2_ASAP7_75t_R g1378 ( 
.A(n_1113),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1108),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1105),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1105),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_SL g1383 ( 
.A(n_1097),
.B(n_914),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1132),
.A2(n_1219),
.B(n_1129),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_SL g1387 ( 
.A1(n_1142),
.A2(n_915),
.B(n_1225),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1139),
.B(n_844),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1186),
.B(n_915),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1136),
.A2(n_1098),
.B1(n_1097),
.B2(n_915),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1186),
.B(n_915),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1186),
.B(n_915),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1139),
.B(n_844),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1174),
.B(n_844),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1144),
.C(n_1134),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1131),
.B(n_915),
.C(n_1134),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1100),
.A2(n_915),
.B(n_1090),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1128),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1136),
.A2(n_914),
.B1(n_705),
.B2(n_699),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1131),
.A2(n_915),
.B(n_1144),
.C(n_1134),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1094),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1211),
.A2(n_1100),
.B(n_1219),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1376),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1295),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1348),
.A2(n_1401),
.B1(n_1396),
.B2(n_1363),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1383),
.A2(n_1339),
.B1(n_1397),
.B2(n_1290),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1399),
.B(n_1354),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1303),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1367),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1397),
.A2(n_1390),
.B1(n_1355),
.B2(n_1335),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1286),
.B(n_1337),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1324),
.Y(n_1414)
);

CKINVDCx6p67_ASAP7_75t_R g1415 ( 
.A(n_1345),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1245),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1334),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1399),
.B(n_1354),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1289),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1310),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1390),
.A2(n_1357),
.B1(n_1358),
.B2(n_1275),
.Y(n_1421)
);

BUFx2_ASAP7_75t_SL g1422 ( 
.A(n_1287),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1343),
.A2(n_1368),
.B(n_1340),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1305),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1272),
.Y(n_1425)
);

BUFx10_ASAP7_75t_L g1426 ( 
.A(n_1291),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1399),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1274),
.A2(n_1278),
.B1(n_1387),
.B2(n_1307),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1381),
.B(n_1332),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1276),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1275),
.A2(n_1300),
.B1(n_1314),
.B2(n_1311),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1352),
.A2(n_1389),
.B1(n_1371),
.B2(n_1377),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1393),
.A2(n_1282),
.B1(n_1297),
.B2(n_1388),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1373),
.A2(n_1394),
.B1(n_1341),
.B2(n_1395),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1239),
.A2(n_1299),
.B1(n_1372),
.B2(n_1349),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1325),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1338),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1344),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1392),
.A2(n_1308),
.B1(n_1251),
.B2(n_1304),
.Y(n_1439)
);

CKINVDCx11_ASAP7_75t_R g1440 ( 
.A(n_1272),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1361),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1307),
.A2(n_1370),
.B1(n_1331),
.B2(n_1374),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1239),
.A2(n_1372),
.B1(n_1349),
.B2(n_1306),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1273),
.A2(n_1320),
.B1(n_1256),
.B2(n_1266),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1325),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1276),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1346),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1320),
.A2(n_1260),
.B1(n_1301),
.B2(n_1316),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1378),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1253),
.A2(n_1280),
.B1(n_1296),
.B2(n_1258),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1350),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1276),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1279),
.A2(n_1281),
.B1(n_1402),
.B2(n_1360),
.Y(n_1453)
);

BUFx8_ASAP7_75t_L g1454 ( 
.A(n_1302),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1375),
.B(n_1380),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1302),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1302),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1342),
.B(n_1382),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1322),
.B(n_1313),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1319),
.A2(n_1285),
.B1(n_1315),
.B2(n_1268),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1347),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1265),
.A2(n_1293),
.B(n_1253),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1317),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1319),
.A2(n_1315),
.B1(n_1238),
.B2(n_1369),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1238),
.A2(n_1284),
.B1(n_1398),
.B2(n_1391),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1309),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1375),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1380),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1326),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1359),
.A2(n_1321),
.B1(n_1298),
.B2(n_1254),
.Y(n_1472)
);

BUFx10_ASAP7_75t_L g1473 ( 
.A(n_1330),
.Y(n_1473)
);

INVx6_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

BUFx8_ASAP7_75t_L g1475 ( 
.A(n_1315),
.Y(n_1475)
);

INVx3_ASAP7_75t_SL g1476 ( 
.A(n_1333),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1283),
.A2(n_1243),
.B1(n_1248),
.B2(n_1247),
.Y(n_1477)
);

CKINVDCx14_ASAP7_75t_R g1478 ( 
.A(n_1323),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1323),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1323),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1364),
.A2(n_1386),
.B(n_1365),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1294),
.A2(n_1292),
.B1(n_1269),
.B2(n_1267),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1288),
.Y(n_1483)
);

INVx6_ASAP7_75t_L g1484 ( 
.A(n_1328),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1270),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1264),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1329),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1246),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1366),
.A2(n_1384),
.B1(n_1379),
.B2(n_1312),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1250),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1294),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1244),
.B(n_1262),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1261),
.Y(n_1493)
);

CKINVDCx6p67_ASAP7_75t_R g1494 ( 
.A(n_1271),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1250),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1255),
.A2(n_1318),
.B1(n_1277),
.B2(n_1252),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1237),
.A2(n_1263),
.B1(n_1336),
.B2(n_1385),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1403),
.A2(n_1242),
.B1(n_1259),
.B2(n_1362),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1257),
.A2(n_1356),
.B1(n_1259),
.B2(n_1241),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1240),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1351),
.A2(n_1362),
.B1(n_1240),
.B2(n_1259),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1240),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1362),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1241),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1351),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1241),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1325),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1325),
.Y(n_1508)
);

BUFx10_ASAP7_75t_L g1509 ( 
.A(n_1305),
.Y(n_1509)
);

CKINVDCx11_ASAP7_75t_R g1510 ( 
.A(n_1295),
.Y(n_1510)
);

BUFx12f_ASAP7_75t_L g1511 ( 
.A(n_1376),
.Y(n_1511)
);

INVx4_ASAP7_75t_L g1512 ( 
.A(n_1324),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1376),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1324),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1342),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1325),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1361),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1383),
.A2(n_1290),
.B1(n_914),
.B2(n_692),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1345),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1353),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1383),
.A2(n_1290),
.B1(n_914),
.B2(n_692),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1383),
.A2(n_1290),
.B1(n_914),
.B2(n_692),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1340),
.A2(n_1186),
.B1(n_1368),
.B2(n_1397),
.Y(n_1524)
);

INVx5_ASAP7_75t_L g1525 ( 
.A(n_1375),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1361),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1342),
.Y(n_1528)
);

INVx6_ASAP7_75t_L g1529 ( 
.A(n_1399),
.Y(n_1529)
);

BUFx4f_ASAP7_75t_SL g1530 ( 
.A(n_1345),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1399),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1353),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1339),
.B(n_915),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1345),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1345),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1348),
.A2(n_1396),
.B1(n_1401),
.B2(n_1363),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1383),
.A2(n_1290),
.B1(n_914),
.B2(n_692),
.Y(n_1538)
);

CKINVDCx6p67_ASAP7_75t_R g1539 ( 
.A(n_1345),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1342),
.Y(n_1541)
);

BUFx4f_ASAP7_75t_SL g1542 ( 
.A(n_1345),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1339),
.B(n_915),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1383),
.A2(n_1363),
.B1(n_1275),
.B2(n_915),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1547)
);

CKINVDCx6p67_ASAP7_75t_R g1548 ( 
.A(n_1345),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1324),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1286),
.B(n_1337),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1400),
.A2(n_1383),
.B1(n_1339),
.B2(n_1363),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1249),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1342),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1339),
.B(n_915),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1383),
.A2(n_1363),
.B1(n_1275),
.B2(n_915),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1249),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1324),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1361),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1492),
.B(n_1420),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1493),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1516),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1490),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1495),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1481),
.A2(n_1498),
.B(n_1497),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1545),
.B(n_1555),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1545),
.B(n_1555),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1483),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1479),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1480),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1410),
.B(n_1416),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1421),
.B(n_1528),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_SL g1572 ( 
.A(n_1449),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1464),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1525),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1417),
.B(n_1437),
.Y(n_1575)
);

INVx4_ASAP7_75t_SL g1576 ( 
.A(n_1474),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1541),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1496),
.A2(n_1489),
.B(n_1485),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1500),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1438),
.B(n_1447),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1487),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1432),
.B(n_1533),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1554),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1421),
.B(n_1458),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1503),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1451),
.B(n_1552),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1497),
.A2(n_1496),
.B(n_1489),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1519),
.A2(n_1538),
.B1(n_1523),
.B2(n_1522),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1412),
.B(n_1407),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1486),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1423),
.B(n_1524),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1406),
.B(n_1513),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1556),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1501),
.A2(n_1499),
.B(n_1450),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1404),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1478),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1478),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1429),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1484),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1477),
.A2(n_1443),
.B(n_1453),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1459),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1443),
.A2(n_1453),
.B(n_1505),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1502),
.B(n_1525),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1537),
.A2(n_1439),
.B1(n_1475),
.B2(n_1491),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1504),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1405),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1406),
.B(n_1513),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1474),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1527),
.B(n_1536),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1468),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1501),
.A2(n_1450),
.B(n_1467),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1488),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1506),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1467),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1475),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1525),
.Y(n_1617)
);

AO21x2_ASAP7_75t_L g1618 ( 
.A1(n_1462),
.A2(n_1466),
.B(n_1463),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1470),
.Y(n_1619)
);

BUFx4f_ASAP7_75t_SL g1620 ( 
.A(n_1511),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1408),
.A2(n_1428),
.B(n_1412),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1472),
.A2(n_1435),
.B(n_1455),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1435),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1409),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1518),
.B(n_1526),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1409),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1472),
.A2(n_1455),
.B(n_1469),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1418),
.Y(n_1628)
);

AO21x1_ASAP7_75t_L g1629 ( 
.A1(n_1408),
.A2(n_1546),
.B(n_1536),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1448),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1465),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1469),
.A2(n_1418),
.B(n_1527),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1460),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1474),
.Y(n_1634)
);

INVxp67_ASAP7_75t_R g1635 ( 
.A(n_1413),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1430),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1446),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1442),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1452),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1470),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1444),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1454),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1482),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1540),
.A2(n_1543),
.B(n_1551),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1452),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1456),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1540),
.B(n_1546),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1543),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1547),
.B(n_1551),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1547),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1454),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1550),
.B(n_1431),
.Y(n_1652)
);

INVx5_ASAP7_75t_SL g1653 ( 
.A(n_1494),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1476),
.Y(n_1654)
);

OA21x2_ASAP7_75t_L g1655 ( 
.A1(n_1431),
.A2(n_1434),
.B(n_1517),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1427),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1476),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1473),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1558),
.B(n_1441),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1473),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1457),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1427),
.A2(n_1531),
.B(n_1529),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1461),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1425),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1426),
.B(n_1532),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1654),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1594),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1635),
.B(n_1426),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1635),
.B(n_1411),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1565),
.A2(n_1508),
.B(n_1507),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1565),
.A2(n_1471),
.B1(n_1514),
.B2(n_1422),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1602),
.B(n_1557),
.Y(n_1673)
);

BUFx12f_ASAP7_75t_L g1674 ( 
.A(n_1607),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1577),
.B(n_1440),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1561),
.B(n_1414),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1583),
.B(n_1436),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1613),
.B(n_1445),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1580),
.B(n_1414),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1566),
.A2(n_1512),
.B(n_1557),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1613),
.B(n_1445),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1566),
.A2(n_1445),
.B1(n_1511),
.B2(n_1419),
.Y(n_1682)
);

AO21x2_ASAP7_75t_L g1683 ( 
.A1(n_1621),
.A2(n_1532),
.B(n_1521),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1570),
.Y(n_1684)
);

AO32x2_ASAP7_75t_L g1685 ( 
.A1(n_1634),
.A2(n_1424),
.A3(n_1549),
.B1(n_1515),
.B2(n_1510),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1584),
.B(n_1515),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1592),
.A2(n_1629),
.B1(n_1608),
.B2(n_1649),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1570),
.B(n_1415),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1575),
.B(n_1581),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1590),
.A2(n_1542),
.B1(n_1530),
.B2(n_1539),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1575),
.B(n_1548),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1587),
.Y(n_1692)
);

AO32x2_ASAP7_75t_L g1693 ( 
.A1(n_1656),
.A2(n_1530),
.A3(n_1542),
.B1(n_1509),
.B2(n_1534),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1605),
.A2(n_1509),
.B1(n_1520),
.B2(n_1535),
.C(n_1638),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1612),
.A2(n_1629),
.B(n_1623),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1587),
.B(n_1654),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1638),
.B(n_1643),
.C(n_1615),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1589),
.A2(n_1593),
.B1(n_1610),
.B2(n_1643),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1572),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1608),
.A2(n_1647),
.B1(n_1649),
.B2(n_1644),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1623),
.B(n_1615),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1642),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1573),
.B(n_1665),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1611),
.Y(n_1704)
);

BUFx4f_ASAP7_75t_SL g1705 ( 
.A(n_1596),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1605),
.A2(n_1641),
.B(n_1631),
.C(n_1585),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1585),
.B(n_1571),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1569),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1659),
.B(n_1625),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1662),
.B(n_1664),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1612),
.A2(n_1601),
.B(n_1564),
.Y(n_1711)
);

O2A1O1Ixp33_ASAP7_75t_SL g1712 ( 
.A1(n_1658),
.A2(n_1660),
.B(n_1620),
.C(n_1607),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1593),
.A2(n_1610),
.B(n_1647),
.C(n_1633),
.Y(n_1713)
);

AND2x6_ASAP7_75t_L g1714 ( 
.A(n_1609),
.B(n_1604),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1631),
.B(n_1641),
.C(n_1630),
.Y(n_1715)
);

OAI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1630),
.A2(n_1601),
.B(n_1571),
.C(n_1644),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1614),
.B(n_1657),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1559),
.B(n_1612),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1569),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1576),
.B(n_1604),
.Y(n_1720)
);

AO21x2_ASAP7_75t_L g1721 ( 
.A1(n_1606),
.A2(n_1595),
.B(n_1650),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1644),
.A2(n_1603),
.B(n_1648),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1576),
.B(n_1604),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1657),
.B(n_1636),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1657),
.B(n_1646),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1648),
.A2(n_1650),
.B1(n_1652),
.B2(n_1595),
.C(n_1661),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1666),
.B(n_1616),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1614),
.B(n_1652),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1642),
.B(n_1651),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1666),
.B(n_1616),
.Y(n_1730)
);

BUFx2_ASAP7_75t_SL g1731 ( 
.A(n_1651),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1661),
.A2(n_1622),
.B(n_1632),
.C(n_1582),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1637),
.B(n_1639),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1622),
.A2(n_1632),
.B(n_1582),
.C(n_1609),
.Y(n_1734)
);

AO32x2_ASAP7_75t_L g1735 ( 
.A1(n_1656),
.A2(n_1574),
.A3(n_1617),
.B1(n_1595),
.B2(n_1568),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1582),
.A2(n_1609),
.B(n_1598),
.C(n_1597),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1564),
.A2(n_1578),
.B(n_1588),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1607),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1597),
.A2(n_1598),
.B(n_1603),
.C(n_1627),
.Y(n_1739)
);

NAND4xp25_ASAP7_75t_L g1740 ( 
.A(n_1560),
.B(n_1640),
.C(n_1567),
.D(n_1619),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1591),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1644),
.A2(n_1653),
.B1(n_1655),
.B2(n_1578),
.Y(n_1742)
);

NOR2x1_ASAP7_75t_SL g1743 ( 
.A(n_1618),
.B(n_1574),
.Y(n_1743)
);

NAND4xp25_ASAP7_75t_L g1744 ( 
.A(n_1560),
.B(n_1640),
.C(n_1567),
.D(n_1619),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1591),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1696),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1718),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1741),
.B(n_1559),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1667),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1677),
.B(n_1559),
.Y(n_1750)
);

NOR2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1674),
.B(n_1656),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1689),
.B(n_1578),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1694),
.A2(n_1655),
.B1(n_1624),
.B2(n_1628),
.C(n_1626),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1741),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1704),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1707),
.B(n_1578),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1724),
.B(n_1588),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1708),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1719),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1745),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1714),
.B(n_1576),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1668),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1695),
.B(n_1562),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1721),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1684),
.Y(n_1765)
);

CKINVDCx11_ASAP7_75t_R g1766 ( 
.A(n_1738),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1725),
.B(n_1567),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1714),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1692),
.B(n_1727),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1677),
.B(n_1563),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1717),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1714),
.B(n_1600),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1701),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1701),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1730),
.B(n_1568),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1735),
.B(n_1637),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1714),
.B(n_1720),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1705),
.B(n_1653),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1735),
.B(n_1645),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1728),
.B(n_1563),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1698),
.A2(n_1655),
.B1(n_1653),
.B2(n_1599),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1733),
.B(n_1586),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1726),
.B(n_1579),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1726),
.B(n_1711),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1705),
.B(n_1653),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1678),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1687),
.A2(n_1698),
.B1(n_1706),
.B2(n_1713),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1678),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1681),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1720),
.B(n_1600),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1754),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1787),
.A2(n_1697),
.B(n_1694),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1787),
.A2(n_1700),
.B1(n_1715),
.B2(n_1742),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1754),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1770),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1763),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1766),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1784),
.A2(n_1672),
.B(n_1711),
.C(n_1671),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1770),
.B(n_1690),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1784),
.A2(n_1716),
.B(n_1742),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1752),
.B(n_1743),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1757),
.B(n_1737),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1755),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1773),
.B(n_1686),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1757),
.B(n_1737),
.Y(n_1805)
);

OAI33xp33_ASAP7_75t_L g1806 ( 
.A1(n_1783),
.A2(n_1672),
.A3(n_1686),
.B1(n_1690),
.B2(n_1682),
.B3(n_1673),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1764),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1773),
.B(n_1716),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1761),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1748),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1768),
.B(n_1722),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1774),
.B(n_1722),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1783),
.A2(n_1700),
.B1(n_1655),
.B2(n_1683),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1768),
.B(n_1739),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1758),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1776),
.B(n_1732),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1774),
.B(n_1681),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1776),
.B(n_1734),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1781),
.A2(n_1753),
.B1(n_1682),
.B2(n_1680),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1786),
.B(n_1740),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1777),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1758),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1786),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1749),
.Y(n_1824)
);

INVx4_ASAP7_75t_L g1825 ( 
.A(n_1777),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1759),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1747),
.A2(n_1736),
.B(n_1671),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1777),
.Y(n_1828)
);

AOI33xp33_ASAP7_75t_L g1829 ( 
.A1(n_1788),
.A2(n_1679),
.A3(n_1691),
.B1(n_1688),
.B2(n_1702),
.B3(n_1712),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1746),
.A2(n_1653),
.B1(n_1680),
.B2(n_1709),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1756),
.B(n_1744),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1779),
.B(n_1685),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1777),
.Y(n_1833)
);

BUFx8_ASAP7_75t_L g1834 ( 
.A(n_1761),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1761),
.B(n_1723),
.Y(n_1835)
);

NAND2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1828),
.B(n_1663),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1795),
.B(n_1788),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1832),
.B(n_1775),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1812),
.B(n_1780),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1812),
.B(n_1780),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1832),
.B(n_1775),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1832),
.B(n_1769),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1801),
.B(n_1789),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1834),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1807),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1815),
.Y(n_1846)
);

INVxp67_ASAP7_75t_SL g1847 ( 
.A(n_1808),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1815),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1822),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1822),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1828),
.B(n_1769),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1834),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1795),
.B(n_1789),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1828),
.B(n_1767),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1823),
.B(n_1759),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1827),
.B(n_1750),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1808),
.B(n_1771),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1797),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1833),
.B(n_1772),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1823),
.B(n_1760),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1826),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1825),
.B(n_1821),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1807),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1791),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1804),
.B(n_1782),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1797),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1804),
.B(n_1820),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1833),
.B(n_1772),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1807),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1801),
.B(n_1779),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1820),
.B(n_1782),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1825),
.B(n_1772),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1826),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1817),
.B(n_1765),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1803),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1791),
.B(n_1760),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1794),
.B(n_1762),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1803),
.Y(n_1878)
);

OA21x2_ASAP7_75t_SL g1879 ( 
.A1(n_1792),
.A2(n_1685),
.B(n_1790),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1847),
.B(n_1817),
.Y(n_1880)
);

NOR2xp67_ASAP7_75t_L g1881 ( 
.A(n_1844),
.B(n_1825),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1858),
.B(n_1797),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1845),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1864),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1851),
.B(n_1825),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1864),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1847),
.B(n_1799),
.Y(n_1887)
);

OAI21xp33_ASAP7_75t_L g1888 ( 
.A1(n_1867),
.A2(n_1798),
.B(n_1792),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1846),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1867),
.B(n_1831),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1856),
.A2(n_1806),
.B(n_1800),
.Y(n_1891)
);

OAI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1879),
.A2(n_1819),
.B1(n_1800),
.B2(n_1831),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1871),
.B(n_1831),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1851),
.B(n_1825),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1858),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1846),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1858),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1848),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1842),
.B(n_1821),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1848),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1849),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1849),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1844),
.B(n_1821),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1866),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1842),
.B(n_1821),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1844),
.B(n_1835),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1871),
.B(n_1810),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1850),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1866),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1850),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1857),
.B(n_1799),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1838),
.B(n_1801),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1838),
.B(n_1809),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1861),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1866),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1841),
.B(n_1854),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1861),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1852),
.B(n_1835),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1841),
.B(n_1809),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1854),
.B(n_1809),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1857),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1859),
.B(n_1809),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1873),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1839),
.B(n_1810),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1859),
.B(n_1809),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1907),
.B(n_1839),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1889),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1916),
.B(n_1868),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1889),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1891),
.B(n_1843),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1916),
.B(n_1868),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1906),
.B(n_1872),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1907),
.B(n_1840),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1888),
.B(n_1887),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1896),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1911),
.B(n_1843),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1896),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1906),
.B(n_1872),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1898),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1906),
.B(n_1872),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1918),
.B(n_1872),
.Y(n_1941)
);

AOI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1892),
.A2(n_1798),
.B(n_1879),
.C(n_1806),
.Y(n_1942)
);

NAND2x1p5_ASAP7_75t_L g1943 ( 
.A(n_1882),
.B(n_1852),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1890),
.B(n_1840),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1918),
.B(n_1870),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1898),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1900),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1899),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1890),
.B(n_1865),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1900),
.Y(n_1950)
);

XNOR2xp5_ASAP7_75t_L g1951 ( 
.A(n_1921),
.B(n_1751),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1893),
.B(n_1865),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1899),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1901),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1918),
.B(n_1870),
.Y(n_1955)
);

NAND2x1p5_ASAP7_75t_L g1956 ( 
.A(n_1895),
.B(n_1852),
.Y(n_1956)
);

AND2x4_ASAP7_75t_SL g1957 ( 
.A(n_1903),
.B(n_1675),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1893),
.B(n_1874),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1895),
.Y(n_1959)
);

NAND2x1p5_ASAP7_75t_SL g1960 ( 
.A(n_1909),
.B(n_1814),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1909),
.B(n_1862),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1915),
.A2(n_1793),
.B(n_1827),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1942),
.A2(n_1793),
.B1(n_1904),
.B2(n_1881),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1929),
.Y(n_1964)
);

O2A1O1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1934),
.A2(n_1897),
.B(n_1880),
.C(n_1886),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1957),
.Y(n_1966)
);

NOR3xp33_ASAP7_75t_L g1967 ( 
.A(n_1930),
.B(n_1897),
.C(n_1880),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1957),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1929),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1945),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1935),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1956),
.Y(n_1972)
);

AOI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1960),
.A2(n_1816),
.B1(n_1796),
.B2(n_1818),
.C(n_1886),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1962),
.A2(n_1819),
.B1(n_1903),
.B2(n_1814),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1935),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1959),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_1959),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1951),
.A2(n_1884),
.B(n_1816),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1951),
.A2(n_1903),
.B1(n_1814),
.B2(n_1816),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1944),
.B(n_1952),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1956),
.B(n_1699),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1945),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1944),
.B(n_1924),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_SL g1984 ( 
.A(n_1943),
.B(n_1829),
.C(n_1924),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1943),
.A2(n_1860),
.B(n_1855),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1927),
.Y(n_1986)
);

OAI21xp33_ASAP7_75t_SL g1987 ( 
.A1(n_1955),
.A2(n_1905),
.B(n_1912),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1960),
.A2(n_1818),
.B(n_1829),
.C(n_1805),
.Y(n_1988)
);

O2A1O1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1943),
.A2(n_1902),
.B(n_1914),
.C(n_1910),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1952),
.B(n_1908),
.Y(n_1990)
);

OAI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1974),
.A2(n_1949),
.B1(n_1958),
.B2(n_1933),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1977),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1973),
.A2(n_1984),
.B1(n_1963),
.B2(n_1967),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1969),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1965),
.A2(n_1956),
.B(n_1939),
.C(n_1946),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1969),
.Y(n_1996)
);

NAND2xp33_ASAP7_75t_SL g1997 ( 
.A(n_1980),
.B(n_1955),
.Y(n_1997)
);

OAI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1988),
.A2(n_1933),
.B(n_1926),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1970),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1976),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1977),
.B(n_1949),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1990),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_1967),
.A2(n_1958),
.B(n_1926),
.C(n_1954),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_SL g2004 ( 
.A1(n_1979),
.A2(n_1818),
.B1(n_1941),
.B2(n_1940),
.Y(n_2004)
);

A2O1A1Ixp33_ASAP7_75t_L g2005 ( 
.A1(n_1978),
.A2(n_1936),
.B(n_1950),
.C(n_1947),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1976),
.Y(n_2006)
);

OAI32xp33_ASAP7_75t_L g2007 ( 
.A1(n_1987),
.A2(n_1953),
.A3(n_1948),
.B1(n_1937),
.B2(n_1941),
.Y(n_2007)
);

OA21x2_ASAP7_75t_L g2008 ( 
.A1(n_1964),
.A2(n_1883),
.B(n_1961),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1989),
.A2(n_1948),
.B(n_1953),
.C(n_1914),
.Y(n_2009)
);

OAI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1983),
.A2(n_1836),
.B1(n_1813),
.B2(n_1796),
.C(n_1883),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1982),
.B(n_1928),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1971),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_2008),
.Y(n_2013)
);

AOI221xp5_ASAP7_75t_L g2014 ( 
.A1(n_1991),
.A2(n_1975),
.B1(n_1986),
.B2(n_1985),
.C(n_1972),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1998),
.B(n_1966),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1992),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_2000),
.Y(n_2017)
);

AO22x1_ASAP7_75t_L g2018 ( 
.A1(n_2006),
.A2(n_1981),
.B1(n_1968),
.B2(n_1961),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2001),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1991),
.B(n_1928),
.Y(n_2020)
);

OAI31xp33_ASAP7_75t_L g2021 ( 
.A1(n_2005),
.A2(n_1836),
.A3(n_1802),
.B(n_1805),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_2003),
.B(n_1931),
.Y(n_2022)
);

AOI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_1993),
.A2(n_1910),
.B1(n_1902),
.B2(n_1901),
.C(n_1923),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1997),
.Y(n_2024)
);

XNOR2x1_ASAP7_75t_L g2025 ( 
.A(n_2008),
.B(n_1751),
.Y(n_2025)
);

AOI31xp33_ASAP7_75t_L g2026 ( 
.A1(n_2002),
.A2(n_1940),
.A3(n_1938),
.B(n_1932),
.Y(n_2026)
);

NOR4xp25_ASAP7_75t_L g2027 ( 
.A(n_1994),
.B(n_1996),
.C(n_1995),
.D(n_2005),
.Y(n_2027)
);

NOR3x1_ASAP7_75t_L g2028 ( 
.A(n_2018),
.B(n_2011),
.C(n_2012),
.Y(n_2028)
);

NOR2xp67_ASAP7_75t_L g2029 ( 
.A(n_2017),
.B(n_1999),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2013),
.Y(n_2030)
);

OAI211xp5_ASAP7_75t_L g2031 ( 
.A1(n_2027),
.A2(n_2007),
.B(n_2009),
.C(n_2004),
.Y(n_2031)
);

NAND4xp75_ASAP7_75t_L g2032 ( 
.A(n_2015),
.B(n_2008),
.C(n_1999),
.D(n_1938),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2027),
.B(n_1931),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_2021),
.B(n_1961),
.Y(n_2034)
);

NAND3xp33_ASAP7_75t_SL g2035 ( 
.A(n_2014),
.B(n_2010),
.C(n_1932),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2016),
.Y(n_2036)
);

NAND3xp33_ASAP7_75t_SL g2037 ( 
.A(n_2021),
.B(n_1836),
.C(n_1905),
.Y(n_2037)
);

INVxp67_ASAP7_75t_L g2038 ( 
.A(n_2020),
.Y(n_2038)
);

NAND4xp25_ASAP7_75t_L g2039 ( 
.A(n_2023),
.B(n_1729),
.C(n_1703),
.D(n_1785),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_2033),
.A2(n_2025),
.B1(n_2022),
.B2(n_2019),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2029),
.B(n_2024),
.Y(n_2041)
);

NAND4xp25_ASAP7_75t_SL g2042 ( 
.A(n_2031),
.B(n_2026),
.C(n_1885),
.D(n_1894),
.Y(n_2042)
);

O2A1O1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_2038),
.A2(n_2030),
.B(n_2035),
.C(n_2036),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2037),
.A2(n_1917),
.B1(n_1802),
.B2(n_1805),
.C(n_1870),
.Y(n_2044)
);

OAI21xp33_ASAP7_75t_L g2045 ( 
.A1(n_2034),
.A2(n_1894),
.B(n_1885),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2032),
.A2(n_1802),
.B1(n_1813),
.B2(n_1710),
.C(n_1863),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_2041),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2040),
.A2(n_2028),
.B1(n_1912),
.B2(n_1925),
.Y(n_2048)
);

NOR3xp33_ASAP7_75t_L g2049 ( 
.A(n_2043),
.B(n_2039),
.C(n_1778),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_2046),
.A2(n_1863),
.B1(n_1869),
.B2(n_1845),
.C(n_1811),
.Y(n_2050)
);

AOI211xp5_ASAP7_75t_SL g2051 ( 
.A1(n_2045),
.A2(n_1920),
.B(n_1922),
.C(n_1925),
.Y(n_2051)
);

O2A1O1Ixp33_ASAP7_75t_L g2052 ( 
.A1(n_2042),
.A2(n_1836),
.B(n_1860),
.C(n_1855),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_2044),
.A2(n_1845),
.B1(n_1863),
.B2(n_1869),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_2041),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2054),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_L g2056 ( 
.A(n_2047),
.B(n_2048),
.C(n_2052),
.Y(n_2056)
);

AO22x2_ASAP7_75t_L g2057 ( 
.A1(n_2049),
.A2(n_1913),
.B1(n_1919),
.B2(n_1922),
.Y(n_2057)
);

NAND4xp75_ASAP7_75t_L g2058 ( 
.A(n_2050),
.B(n_1919),
.C(n_1913),
.D(n_1920),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_2051),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2053),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2055),
.B(n_1862),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_SL g2062 ( 
.A(n_2060),
.B(n_1830),
.C(n_1685),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_2059),
.A2(n_1877),
.B(n_1876),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_2061),
.Y(n_2064)
);

OAI22x1_ASAP7_75t_L g2065 ( 
.A1(n_2064),
.A2(n_2056),
.B1(n_2057),
.B2(n_2062),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2065),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_2065),
.A2(n_2057),
.B1(n_2063),
.B2(n_2058),
.Y(n_2067)
);

OAI22x1_ASAP7_75t_L g2068 ( 
.A1(n_2066),
.A2(n_2067),
.B1(n_1862),
.B2(n_1676),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2066),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_2069),
.Y(n_2070)
);

OAI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_2068),
.A2(n_1853),
.B(n_1837),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2070),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2072),
.A2(n_2071),
.B(n_1853),
.Y(n_2073)
);

OAI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2073),
.A2(n_1874),
.B1(n_1875),
.B2(n_1878),
.Y(n_2074)
);

OAI221xp5_ASAP7_75t_R g2075 ( 
.A1(n_2074),
.A2(n_1693),
.B1(n_1731),
.B2(n_1862),
.C(n_1824),
.Y(n_2075)
);

AOI211xp5_ASAP7_75t_L g2076 ( 
.A1(n_2075),
.A2(n_1669),
.B(n_1670),
.C(n_1830),
.Y(n_2076)
);


endmodule