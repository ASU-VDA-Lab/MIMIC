module fake_netlist_6_1558_n_1783 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1783);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1783;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_31),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_45),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_92),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_45),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_7),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_3),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_115),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_29),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_19),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_43),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_93),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_65),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_55),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_75),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_100),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_72),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_31),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_10),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_95),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_112),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_3),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_136),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_29),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_38),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_6),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_10),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_19),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_9),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_67),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_54),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_27),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_20),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_18),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_56),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_85),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_48),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_51),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_36),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_50),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_40),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_79),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_37),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_44),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_130),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_52),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_94),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_120),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_39),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_5),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_154),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_140),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_41),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_150),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_44),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_8),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_80),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_78),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_143),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_119),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_73),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_145),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_81),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_83),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_109),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_144),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_6),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_121),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_89),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_149),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_53),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_137),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_15),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_99),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_74),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_14),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_23),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_4),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_60),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_8),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_30),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_14),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_12),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_116),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_108),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_141),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_32),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_22),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_24),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_9),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_61),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_124),
.Y(n_307)
);

CKINVDCx11_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_35),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_195),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_157),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_176),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_308),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_157),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_156),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_216),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_160),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_161),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_160),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_171),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_173),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_163),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_170),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_166),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_174),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_219),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_166),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_231),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_248),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_169),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_181),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_181),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_186),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_186),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_170),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_218),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_305),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_195),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_196),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_196),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_158),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_158),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_210),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_179),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_210),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_226),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_159),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_226),
.Y(n_356)
);

BUFx2_ASAP7_75t_SL g357 ( 
.A(n_297),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_162),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_232),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_225),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_159),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_232),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_274),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_305),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_182),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_277),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_164),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_244),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_283),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_283),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_183),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_184),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_188),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_199),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_202),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_290),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_291),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_291),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_203),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_165),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_315),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_384),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_297),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_205),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

BUFx8_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_342),
.A2(n_221),
.B1(n_201),
.B2(n_178),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_R g400 ( 
.A(n_313),
.B(n_168),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_323),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_195),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_324),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_325),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_361),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_357),
.B(n_209),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_331),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_165),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_345),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_311),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_180),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_311),
.Y(n_421)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_254),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_355),
.B(n_227),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_322),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_352),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_314),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_312),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_314),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_316),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

CKINVDCx11_ASAP7_75t_R g432 ( 
.A(n_375),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_317),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_327),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_334),
.A2(n_271),
.B1(n_220),
.B2(n_252),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_366),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_328),
.A2(n_197),
.B1(n_286),
.B2(n_304),
.Y(n_437)
);

NAND2x1_ASAP7_75t_L g438 ( 
.A(n_330),
.B(n_195),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_330),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_317),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_321),
.B(n_187),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_321),
.B(n_254),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_329),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_318),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_318),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_333),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_332),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_336),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_336),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

NOR2x1p5_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_293),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_383),
.Y(n_456)
);

NOR3xp33_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_370),
.C(n_266),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_427),
.C(n_417),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_415),
.B(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_400),
.B(n_335),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_393),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_408),
.B(n_172),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_187),
.Y(n_465)
);

NOR2x1p5_ASAP7_75t_L g466 ( 
.A(n_409),
.B(n_293),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_348),
.B1(n_200),
.B2(n_309),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_393),
.B(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_419),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_177),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_390),
.A2(n_302),
.B1(n_300),
.B2(n_304),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_412),
.B(n_172),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_430),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

AND2x2_ASAP7_75t_SL g478 ( 
.A(n_445),
.B(n_272),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_445),
.B(n_272),
.Y(n_481)
);

BUFx8_ASAP7_75t_SL g482 ( 
.A(n_424),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_419),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_236),
.B1(n_239),
.B2(n_242),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_431),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_390),
.A2(n_418),
.B1(n_422),
.B2(n_427),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_423),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_423),
.B(n_185),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_441),
.B(n_319),
.Y(n_495)
);

INVx8_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_410),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_389),
.A2(n_441),
.B1(n_442),
.B2(n_414),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_441),
.B(n_195),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_442),
.B(n_215),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_399),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_391),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_396),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_436),
.B(n_447),
.Y(n_514)
);

AND3x2_ASAP7_75t_L g515 ( 
.A(n_447),
.B(n_299),
.C(n_276),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_418),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_440),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_442),
.B(n_237),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_397),
.A2(n_259),
.B1(n_225),
.B2(n_306),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_442),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_438),
.A2(n_191),
.B(n_190),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_404),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_443),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_414),
.B(n_319),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

BUFx6f_ASAP7_75t_SL g531 ( 
.A(n_389),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_440),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_407),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_398),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_402),
.B(n_238),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_450),
.B(n_172),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_450),
.B(n_397),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_438),
.A2(n_191),
.B(n_190),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_389),
.B(n_193),
.C(n_189),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_446),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_394),
.B(n_299),
.C(n_276),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_389),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_413),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_397),
.B(n_306),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_398),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_403),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_413),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_420),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_420),
.Y(n_557)
);

CKINVDCx6p67_ASAP7_75t_R g558 ( 
.A(n_432),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_386),
.B(n_292),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_386),
.B(n_406),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_414),
.B(n_434),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_416),
.Y(n_562)
);

INVxp33_ASAP7_75t_SL g563 ( 
.A(n_399),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_416),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_434),
.A2(n_300),
.B1(n_302),
.B2(n_240),
.Y(n_565)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_385),
.A2(n_198),
.B(n_192),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_439),
.B(n_194),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_397),
.B(n_306),
.Y(n_568)
);

BUFx6f_ASAP7_75t_SL g569 ( 
.A(n_439),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_394),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_416),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_448),
.B(n_245),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_448),
.A2(n_235),
.B1(n_222),
.B2(n_303),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_451),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_449),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_386),
.B(n_251),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_421),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_403),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_449),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_452),
.A2(n_192),
.B1(n_198),
.B2(n_204),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_386),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_452),
.B(n_208),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_421),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_421),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_453),
.B(n_255),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_406),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_426),
.B(n_240),
.C(n_298),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_426),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_406),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_429),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_429),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_406),
.B(n_256),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_429),
.B(n_213),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_433),
.B(n_214),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_385),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_385),
.Y(n_598)
);

AND3x2_ASAP7_75t_L g599 ( 
.A(n_433),
.B(n_241),
.C(n_298),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_388),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_433),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_388),
.B(n_258),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_444),
.B(n_260),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_546),
.B(n_523),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_463),
.B(n_388),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_478),
.B(n_262),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_263),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_516),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_468),
.B(n_392),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_478),
.A2(n_267),
.B1(n_264),
.B2(n_307),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_478),
.A2(n_224),
.B1(n_265),
.B2(n_278),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_562),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_579),
.B(n_561),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_579),
.B(n_392),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_495),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_523),
.Y(n_617)
);

AND2x4_ASAP7_75t_SL g618 ( 
.A(n_476),
.B(n_259),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_516),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_481),
.A2(n_458),
.B1(n_490),
.B2(n_494),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_481),
.B(n_223),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_561),
.B(n_392),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_481),
.B(n_273),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_395),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_533),
.B(n_279),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_228),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_541),
.B(n_281),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_533),
.B(n_282),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_533),
.B(n_287),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_593),
.B(n_501),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_482),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_471),
.A2(n_233),
.B1(n_265),
.B2(n_278),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_495),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_L g635 ( 
.A(n_457),
.B(n_294),
.C(n_229),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_506),
.B(n_288),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_529),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_395),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_521),
.B(n_234),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_395),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_567),
.B(n_462),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_511),
.B(n_405),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_522),
.B(n_206),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_511),
.B(n_405),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_602),
.A2(n_403),
.B(n_405),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_512),
.B(n_207),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_529),
.B(n_337),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_512),
.B(n_211),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_570),
.B(n_538),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_518),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_518),
.A2(n_212),
.B1(n_217),
.B2(n_224),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_564),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_519),
.B(n_211),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_476),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_514),
.B(n_444),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_455),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_476),
.B(n_259),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_519),
.B(n_212),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_467),
.B(n_476),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_520),
.A2(n_217),
.B1(n_241),
.B2(n_270),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_595),
.B(n_233),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_459),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_596),
.B(n_465),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_537),
.B(n_243),
.Y(n_666)
);

O2A1O1Ixp5_ASAP7_75t_L g667 ( 
.A1(n_524),
.A2(n_270),
.B(n_444),
.C(n_339),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_455),
.Y(n_668)
);

OAI221xp5_ASAP7_75t_L g669 ( 
.A1(n_565),
.A2(n_339),
.B1(n_382),
.B2(n_381),
.C(n_380),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_464),
.B(n_58),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_576),
.A2(n_403),
.B(n_340),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_465),
.B(n_246),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_527),
.B(n_403),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_527),
.B(n_402),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_466),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_534),
.A2(n_289),
.B1(n_247),
.B2(n_249),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_534),
.B(n_402),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_517),
.B(n_250),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_547),
.B(n_253),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_547),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_549),
.B(n_402),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_582),
.B(n_259),
.Y(n_683)
);

HB1xp67_ASAP7_75t_SL g684 ( 
.A(n_570),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_549),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_555),
.B(n_337),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_571),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_555),
.B(n_257),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_556),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_465),
.B(n_338),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_556),
.A2(n_382),
.B1(n_381),
.B2(n_380),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_557),
.B(n_338),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_456),
.A2(n_261),
.B1(n_268),
.B2(n_269),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_465),
.B(n_275),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_496),
.B(n_280),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_496),
.B(n_284),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_557),
.B(n_340),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_517),
.B(n_285),
.Y(n_699)
);

BUFx5_ASAP7_75t_L g700 ( 
.A(n_489),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_530),
.B(n_295),
.Y(n_701)
);

BUFx6f_ASAP7_75t_SL g702 ( 
.A(n_558),
.Y(n_702)
);

AND2x4_ASAP7_75t_SL g703 ( 
.A(n_558),
.B(n_341),
.Y(n_703)
);

BUFx5_ASAP7_75t_L g704 ( 
.A(n_489),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_509),
.B(n_341),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_571),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_530),
.A2(n_376),
.B(n_372),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_376),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_577),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_372),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_574),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_584),
.B(n_371),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_583),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_584),
.B(n_296),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_532),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_589),
.B(n_371),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_509),
.B(n_369),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_485),
.B(n_369),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_589),
.B(n_367),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_466),
.A2(n_301),
.B1(n_364),
.B2(n_363),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_532),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_563),
.A2(n_367),
.B1(n_364),
.B2(n_363),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_551),
.B(n_362),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_559),
.B(n_362),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_473),
.B(n_1),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_485),
.B(n_359),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_573),
.B(n_359),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_568),
.B(n_356),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_540),
.B(n_356),
.Y(n_731)
);

AND2x6_ASAP7_75t_SL g732 ( 
.A(n_563),
.B(n_354),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_540),
.B(n_354),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_496),
.B(n_353),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_580),
.A2(n_353),
.B1(n_351),
.B2(n_347),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_496),
.B(n_351),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_542),
.B(n_347),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_585),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_572),
.B(n_586),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_585),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_531),
.A2(n_59),
.B1(n_142),
.B2(n_139),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_569),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_542),
.B(n_155),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_503),
.A2(n_4),
.B(n_7),
.C(n_13),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_543),
.B(n_138),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_543),
.B(n_133),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_545),
.B(n_550),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_545),
.B(n_125),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_496),
.B(n_13),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_550),
.B(n_122),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_581),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_513),
.B(n_117),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_544),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_587),
.B(n_113),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_587),
.B(n_105),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_590),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_513),
.B(n_17),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_590),
.Y(n_759)
);

AOI221xp5_ASAP7_75t_L g760 ( 
.A1(n_592),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_591),
.B(n_97),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_597),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_24),
.C(n_25),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_601),
.Y(n_764)
);

OA22x2_ASAP7_75t_L g765 ( 
.A1(n_515),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_591),
.B(n_62),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_594),
.B(n_96),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_597),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_454),
.B(n_91),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_454),
.B(n_90),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_601),
.Y(n_771)
);

INVxp33_ASAP7_75t_L g772 ( 
.A(n_588),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_598),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_460),
.B(n_88),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_599),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_650),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_SL g777 ( 
.A1(n_649),
.A2(n_712),
.B1(n_727),
.B2(n_612),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_616),
.B(n_483),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_614),
.B(n_502),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_659),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_620),
.B(n_513),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_604),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_654),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_634),
.B(n_483),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_662),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_771),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_771),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_609),
.B(n_513),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_609),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_710),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_690),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_690),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_619),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_684),
.Y(n_794)
);

CKINVDCx11_ASAP7_75t_R g795 ( 
.A(n_732),
.Y(n_795)
);

BUFx4f_ASAP7_75t_SL g796 ( 
.A(n_632),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_605),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_681),
.Y(n_798)
);

INVxp33_ASAP7_75t_SL g799 ( 
.A(n_692),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_619),
.B(n_513),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_665),
.A2(n_560),
.B(n_525),
.Y(n_801)
);

NAND2x2_ASAP7_75t_L g802 ( 
.A(n_656),
.B(n_566),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_750),
.B(n_569),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_685),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_717),
.Y(n_805)
);

AND2x6_ASAP7_75t_L g806 ( 
.A(n_631),
.B(n_488),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_621),
.A2(n_531),
.B1(n_569),
.B2(n_480),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_689),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_641),
.B(n_531),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_612),
.B(n_492),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_723),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_621),
.B(n_480),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_705),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_637),
.B(n_472),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_690),
.B(n_513),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_617),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_606),
.B(n_492),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_719),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_622),
.B(n_497),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_633),
.A2(n_588),
.B1(n_598),
.B2(n_600),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_726),
.B(n_497),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_627),
.B(n_472),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_613),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_762),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_768),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_773),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_605),
.B(n_525),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_638),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_720),
.A2(n_460),
.B1(n_469),
.B2(n_498),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_684),
.Y(n_830)
);

OR2x2_ASAP7_75t_SL g831 ( 
.A(n_635),
.B(n_507),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_647),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_SL g833 ( 
.A(n_643),
.B(n_600),
.C(n_502),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_626),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_640),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_604),
.A2(n_623),
.B1(n_608),
.B2(n_639),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_647),
.B(n_469),
.Y(n_837)
);

OR2x2_ASAP7_75t_SL g838 ( 
.A(n_763),
.B(n_484),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_667),
.A2(n_498),
.B(n_499),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_711),
.B(n_499),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_657),
.B(n_479),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_683),
.B(n_536),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_627),
.B(n_578),
.Y(n_843)
);

BUFx12f_ASAP7_75t_L g844 ( 
.A(n_754),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_711),
.B(n_477),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_605),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_660),
.B(n_578),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_772),
.A2(n_639),
.B(n_727),
.C(n_666),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_623),
.A2(n_477),
.B1(n_474),
.B2(n_475),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_664),
.A2(n_525),
.B1(n_479),
.B2(n_508),
.Y(n_850)
);

AND3x1_ASAP7_75t_L g851 ( 
.A(n_666),
.B(n_475),
.C(n_508),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_642),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_728),
.B(n_578),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_644),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_690),
.B(n_474),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_655),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_690),
.B(n_505),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_724),
.B(n_505),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_624),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_607),
.A2(n_487),
.B1(n_488),
.B2(n_493),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_605),
.B(n_611),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_731),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_625),
.A2(n_487),
.B(n_493),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_663),
.A2(n_504),
.B1(n_507),
.B2(n_553),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_703),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_SL g866 ( 
.A(n_677),
.B(n_28),
.C(n_30),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_775),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_651),
.A2(n_504),
.B(n_553),
.C(n_552),
.Y(n_868)
);

AND2x2_ASAP7_75t_SL g869 ( 
.A(n_618),
.B(n_500),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_738),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_610),
.B(n_729),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_680),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_740),
.A2(n_535),
.B1(n_486),
.B2(n_553),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_633),
.A2(n_535),
.B1(n_486),
.B2(n_552),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_742),
.B(n_535),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_733),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_673),
.B(n_28),
.Y(n_877)
);

BUFx12f_ASAP7_75t_L g878 ( 
.A(n_668),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_733),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_615),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_718),
.B(n_461),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_721),
.B(n_461),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_680),
.B(n_688),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_748),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_702),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_686),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_710),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_688),
.B(n_670),
.Y(n_888)
);

AND2x6_ASAP7_75t_SL g889 ( 
.A(n_649),
.B(n_32),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_676),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_725),
.B(n_486),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_646),
.A2(n_552),
.B(n_461),
.C(n_566),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_710),
.Y(n_893)
);

NOR2x1p5_ASAP7_75t_L g894 ( 
.A(n_702),
.B(n_539),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_679),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_693),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_698),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_750),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_710),
.B(n_525),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_708),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_737),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_737),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_649),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_725),
.Y(n_904)
);

NOR2x1p5_ASAP7_75t_L g905 ( 
.A(n_713),
.B(n_539),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_743),
.B(n_526),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_674),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_SL g908 ( 
.A(n_694),
.B(n_33),
.C(n_34),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_724),
.B(n_525),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_628),
.B(n_525),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_652),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_743),
.B(n_752),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_671),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_722),
.B(n_554),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_687),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_700),
.B(n_554),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_695),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_648),
.B(n_554),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_706),
.Y(n_919)
);

AO22x1_ASAP7_75t_L g920 ( 
.A1(n_653),
.A2(n_658),
.B1(n_765),
.B2(n_752),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_752),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_679),
.A2(n_554),
.B1(n_548),
.B2(n_500),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_709),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_700),
.B(n_554),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_752),
.B(n_526),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_700),
.B(n_548),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_730),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_716),
.B(n_548),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_667),
.A2(n_548),
.B(n_500),
.Y(n_929)
);

NOR2x1p5_ASAP7_75t_L g930 ( 
.A(n_767),
.B(n_548),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_699),
.B(n_701),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_765),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_700),
.B(n_500),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_737),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_661),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_700),
.B(n_500),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_700),
.B(n_66),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_704),
.B(n_68),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_704),
.B(n_86),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_714),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_735),
.A2(n_87),
.B(n_76),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_669),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_699),
.B(n_38),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_715),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_704),
.B(n_69),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_704),
.B(n_739),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_704),
.B(n_39),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_704),
.B(n_46),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_734),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_636),
.B(n_47),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_741),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_701),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_745),
.B(n_47),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_757),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_758),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_769),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_770),
.B(n_50),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_753),
.B(n_678),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_759),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_764),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_707),
.B(n_661),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_675),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_682),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_755),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_SL g965 ( 
.A1(n_883),
.A2(n_753),
.B(n_629),
.C(n_630),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_815),
.A2(n_924),
.B(n_916),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_848),
.A2(n_760),
.B(n_629),
.C(n_630),
.Y(n_967)
);

OA21x2_ASAP7_75t_L g968 ( 
.A1(n_839),
.A2(n_672),
.B(n_774),
.Y(n_968)
);

AOI21x1_ASAP7_75t_L g969 ( 
.A1(n_863),
.A2(n_625),
.B(n_766),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_805),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_871),
.A2(n_761),
.B1(n_756),
.B2(n_746),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_789),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_872),
.B(n_696),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_812),
.A2(n_697),
.B(n_751),
.C(n_744),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_937),
.A2(n_645),
.B(n_747),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_776),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_878),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_783),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_908),
.A2(n_749),
.B(n_691),
.C(n_736),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_790),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_SL g981 ( 
.A(n_777),
.B(n_691),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_871),
.B(n_736),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_859),
.B(n_886),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_842),
.A2(n_917),
.B1(n_809),
.B2(n_895),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_829),
.A2(n_836),
.B1(n_822),
.B2(n_810),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_782),
.B(n_799),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_896),
.B(n_897),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_793),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_780),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_900),
.B(n_884),
.Y(n_991)
);

OAI22x1_ASAP7_75t_L g992 ( 
.A1(n_903),
.A2(n_917),
.B1(n_830),
.B2(n_818),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_916),
.A2(n_933),
.B(n_926),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_790),
.Y(n_994)
);

BUFx6f_ASAP7_75t_SL g995 ( 
.A(n_865),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_950),
.A2(n_888),
.B(n_952),
.C(n_877),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_912),
.B(n_890),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_926),
.A2(n_936),
.B(n_933),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_936),
.A2(n_946),
.B(n_861),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_SL g1000 ( 
.A(n_927),
.B(n_935),
.C(n_885),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_947),
.A2(n_948),
.B(n_866),
.C(n_856),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_862),
.B(n_870),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_844),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_961),
.A2(n_931),
.B(n_847),
.C(n_942),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_832),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_785),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_794),
.B(n_867),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_790),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_828),
.B(n_835),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_932),
.B(n_943),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_912),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_798),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_893),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_957),
.A2(n_858),
.B1(n_837),
.B2(n_802),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_816),
.B(n_955),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_804),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_837),
.B(n_841),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_893),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_811),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_791),
.B(n_792),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_810),
.A2(n_961),
.B1(n_807),
.B2(n_782),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_893),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_819),
.A2(n_817),
.B(n_792),
.Y(n_1023)
);

O2A1O1Ixp5_ASAP7_75t_L g1024 ( 
.A1(n_843),
.A2(n_914),
.B(n_781),
.C(n_920),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_808),
.B(n_898),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_853),
.A2(n_957),
.B(n_928),
.C(n_854),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_904),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_786),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_795),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_918),
.A2(n_821),
.B(n_938),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_821),
.A2(n_945),
.B(n_939),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_852),
.B(n_880),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_947),
.A2(n_948),
.B(n_953),
.C(n_955),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_833),
.A2(n_964),
.B(n_879),
.C(n_876),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_960),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_779),
.B(n_907),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_787),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_921),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_850),
.A2(n_791),
.B1(n_792),
.B2(n_840),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_887),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_778),
.B(n_784),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_869),
.B(n_921),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_891),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_SL g1044 ( 
.A(n_934),
.B(n_894),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_791),
.B(n_792),
.Y(n_1045)
);

OAI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_824),
.A2(n_826),
.B(n_825),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_778),
.B(n_784),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_779),
.B(n_962),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_938),
.A2(n_945),
.B(n_881),
.Y(n_1049)
);

CKINVDCx11_ASAP7_75t_R g1050 ( 
.A(n_889),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_814),
.A2(n_891),
.B1(n_806),
.B2(n_840),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_814),
.B(n_845),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_823),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_901),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_953),
.A2(n_845),
.B(n_909),
.C(n_911),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_801),
.A2(n_925),
.B(n_855),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_803),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_803),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_963),
.B(n_882),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_887),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_913),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_901),
.B(n_902),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_963),
.B(n_803),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_953),
.A2(n_923),
.B(n_919),
.C(n_954),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_901),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_831),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_925),
.A2(n_855),
.B(n_857),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_834),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_901),
.B(n_902),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_881),
.B(n_882),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_929),
.A2(n_958),
.B(n_892),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_846),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_846),
.B(n_934),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_838),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_929),
.A2(n_958),
.B(n_857),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_915),
.B(n_951),
.Y(n_1076)
);

OAI21xp33_ASAP7_75t_SL g1077 ( 
.A1(n_874),
.A2(n_905),
.B(n_930),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_902),
.A2(n_797),
.B1(n_958),
.B2(n_873),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_944),
.B(n_959),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_902),
.B(n_956),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_940),
.B(n_949),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_839),
.A2(n_868),
.B(n_849),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_910),
.A2(n_956),
.B(n_851),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_906),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_806),
.B(n_956),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_906),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_806),
.B(n_820),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_806),
.B(n_820),
.Y(n_1088)
);

BUFx4f_ASAP7_75t_L g1089 ( 
.A(n_906),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_899),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_860),
.A2(n_941),
.B(n_922),
.C(n_864),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_899),
.B(n_788),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_800),
.B(n_827),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_875),
.A2(n_812),
.B(n_665),
.Y(n_1094)
);

O2A1O1Ixp5_ASAP7_75t_L g1095 ( 
.A1(n_875),
.A2(n_883),
.B(n_888),
.C(n_848),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_875),
.B(n_871),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_875),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_912),
.B(n_890),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_789),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_848),
.A2(n_871),
.B1(n_829),
.B2(n_883),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_848),
.A2(n_883),
.B(n_872),
.C(n_621),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_805),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_789),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_848),
.A2(n_871),
.B1(n_829),
.B2(n_883),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_871),
.B(n_463),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_SL g1106 ( 
.A1(n_883),
.A2(n_612),
.B(n_961),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_803),
.B(n_844),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_872),
.B(n_478),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_883),
.A2(n_621),
.B1(n_872),
.B2(n_777),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_783),
.Y(n_1110)
);

BUFx8_ASAP7_75t_L g1111 ( 
.A(n_844),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_813),
.B(n_705),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1056),
.A2(n_998),
.B(n_993),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_966),
.A2(n_999),
.B(n_1082),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1116)
);

AOI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_1101),
.A2(n_1104),
.B(n_1100),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1108),
.A2(n_1105),
.B(n_1033),
.C(n_1001),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1036),
.B(n_1009),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1067),
.A2(n_969),
.B(n_975),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1009),
.B(n_988),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_988),
.A2(n_1109),
.B1(n_991),
.B2(n_984),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1065),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_991),
.B(n_1002),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_976),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_1024),
.A2(n_1095),
.B(n_1094),
.C(n_973),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_984),
.B(n_1002),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1075),
.A2(n_1083),
.B(n_1085),
.Y(n_1129)
);

INVx4_ASAP7_75t_SL g1130 ( 
.A(n_1038),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1075),
.A2(n_1083),
.B(n_1085),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_990),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1071),
.A2(n_986),
.A3(n_1021),
.B(n_1087),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1023),
.A2(n_965),
.B(n_1059),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1011),
.B(n_997),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1059),
.A2(n_1071),
.B(n_1070),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1070),
.A2(n_1087),
.B(n_1088),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1032),
.B(n_1048),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_1004),
.A2(n_1026),
.B(n_1034),
.C(n_1096),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1032),
.B(n_1048),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1088),
.A2(n_1078),
.B(n_1097),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_974),
.A2(n_971),
.B(n_1091),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1039),
.A2(n_1055),
.B(n_1020),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_967),
.A2(n_1106),
.B(n_1096),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_985),
.B(n_1112),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_996),
.A2(n_979),
.B(n_1064),
.C(n_981),
.Y(n_1146)
);

NAND3x1_ASAP7_75t_L g1147 ( 
.A(n_1007),
.B(n_1010),
.C(n_1063),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1077),
.A2(n_983),
.B(n_1051),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_983),
.B(n_1052),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_1046),
.A2(n_1014),
.B(n_1084),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_968),
.A2(n_1045),
.B(n_1020),
.Y(n_1151)
);

OAI22x1_ASAP7_75t_L g1152 ( 
.A1(n_1074),
.A2(n_1015),
.B1(n_1058),
.B2(n_1057),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1066),
.A2(n_1047),
.B(n_1041),
.C(n_1076),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1017),
.B(n_1006),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1080),
.A2(n_968),
.B(n_1092),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1072),
.A2(n_1069),
.B(n_1062),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1012),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1081),
.A2(n_1093),
.B(n_1089),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1016),
.B(n_1079),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1061),
.Y(n_1160)
);

NAND2x1_ASAP7_75t_L g1161 ( 
.A(n_1065),
.B(n_1040),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_978),
.B(n_1110),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_SL g1163 ( 
.A1(n_1042),
.A2(n_1054),
.B(n_1038),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_SL g1164 ( 
.A1(n_1025),
.A2(n_1098),
.B(n_997),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1072),
.A2(n_1040),
.B(n_1090),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_982),
.Y(n_1166)
);

AO21x1_ASAP7_75t_L g1167 ( 
.A1(n_1044),
.A2(n_1073),
.B(n_1102),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1028),
.A2(n_1037),
.B(n_970),
.Y(n_1168)
);

AOI31xp67_ASAP7_75t_L g1169 ( 
.A1(n_1019),
.A2(n_1053),
.A3(n_1068),
.B(n_987),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1035),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1054),
.A2(n_1038),
.B(n_1060),
.Y(n_1171)
);

AO21x2_ASAP7_75t_L g1172 ( 
.A1(n_1000),
.A2(n_1089),
.B(n_1086),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_972),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_980),
.A2(n_1022),
.B(n_1005),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_980),
.A2(n_1022),
.B(n_1018),
.C(n_1013),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1054),
.Y(n_1176)
);

AO32x2_ASAP7_75t_L g1177 ( 
.A1(n_1013),
.A2(n_1018),
.A3(n_1060),
.B1(n_1103),
.B2(n_992),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1043),
.A2(n_994),
.B(n_1008),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1043),
.B(n_994),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_989),
.B(n_1099),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_994),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1008),
.A2(n_1043),
.A3(n_1107),
.B(n_995),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1008),
.A2(n_995),
.B(n_1107),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1107),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1027),
.B(n_977),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_SL g1186 ( 
.A1(n_1050),
.A2(n_1111),
.B(n_1003),
.C(n_1029),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1111),
.A2(n_1031),
.B(n_1049),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_SL g1188 ( 
.A(n_978),
.B(n_478),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1071),
.A2(n_1031),
.B(n_1049),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1109),
.B(n_848),
.C(n_883),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1112),
.B(n_705),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1071),
.A2(n_1031),
.A3(n_1049),
.B(n_986),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1101),
.A2(n_848),
.B(n_967),
.C(n_620),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1105),
.B(n_872),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1038),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1101),
.A2(n_848),
.B(n_967),
.C(n_620),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1011),
.B(n_997),
.Y(n_1201)
);

AOI31xp67_ASAP7_75t_L g1202 ( 
.A1(n_1087),
.A2(n_888),
.A3(n_836),
.B(n_1088),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1203)
);

AOI221x1_ASAP7_75t_L g1204 ( 
.A1(n_1094),
.A2(n_1071),
.B1(n_848),
.B2(n_986),
.C(n_1100),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1065),
.B(n_1054),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1106),
.A2(n_1004),
.B(n_1071),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_978),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1056),
.A2(n_998),
.B(n_993),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_976),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_978),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_982),
.Y(n_1213)
);

BUFx2_ASAP7_75t_SL g1214 ( 
.A(n_982),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1029),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1105),
.A2(n_612),
.B1(n_988),
.B2(n_1109),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1071),
.A2(n_1031),
.B(n_1049),
.Y(n_1219)
);

NOR3xp33_ASAP7_75t_SL g1220 ( 
.A(n_981),
.B(n_903),
.C(n_400),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1111),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1056),
.A2(n_998),
.B(n_993),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1101),
.A2(n_848),
.B(n_967),
.C(n_620),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_1064),
.A2(n_1096),
.B(n_1033),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1112),
.B(n_705),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1071),
.A2(n_1031),
.B(n_1049),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_982),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1056),
.A2(n_998),
.B(n_993),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1038),
.Y(n_1233)
);

O2A1O1Ixp5_ASAP7_75t_SL g1234 ( 
.A1(n_1021),
.A2(n_663),
.B(n_883),
.C(n_888),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1109),
.B(n_848),
.C(n_462),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_972),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1105),
.B(n_872),
.Y(n_1237)
);

NAND2xp33_ASAP7_75t_L g1238 ( 
.A(n_1038),
.B(n_848),
.Y(n_1238)
);

NAND2x1p5_ASAP7_75t_L g1239 ( 
.A(n_1065),
.B(n_1054),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1109),
.B(n_848),
.C(n_883),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1056),
.A2(n_998),
.B(n_993),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1010),
.B(n_664),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1031),
.A2(n_1049),
.B(n_1030),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_982),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1109),
.A2(n_664),
.B(n_683),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1105),
.A2(n_612),
.B1(n_988),
.B2(n_1109),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1112),
.B(n_705),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_976),
.Y(n_1249)
);

NAND3x1_ASAP7_75t_L g1250 ( 
.A(n_1109),
.B(n_683),
.C(n_399),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1056),
.A2(n_998),
.B(n_993),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_SL g1252 ( 
.A(n_1109),
.B(n_848),
.C(n_462),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1065),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1126),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1246),
.A2(n_1146),
.B(n_1252),
.C(n_1235),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1120),
.A2(n_1114),
.B(n_1113),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1184),
.B(n_1182),
.Y(n_1257)
);

AO32x2_ASAP7_75t_L g1258 ( 
.A1(n_1122),
.A2(n_1218),
.A3(n_1247),
.B1(n_1204),
.B2(n_1202),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1208),
.Y(n_1259)
);

AO21x2_ASAP7_75t_L g1260 ( 
.A1(n_1187),
.A2(n_1117),
.B(n_1142),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1195),
.A2(n_1225),
.B(n_1200),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1132),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_1221),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1246),
.B(n_1243),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1207),
.A2(n_1229),
.B(n_1224),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1182),
.B(n_1183),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1210),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1249),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1190),
.A2(n_1240),
.B(n_1118),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1197),
.A2(n_1223),
.A3(n_1241),
.B(n_1216),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1244),
.A2(n_1241),
.B(n_1227),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1144),
.A2(n_1167),
.A3(n_1247),
.B(n_1218),
.Y(n_1272)
);

NAND2x1_ASAP7_75t_L g1273 ( 
.A(n_1124),
.B(n_1253),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1128),
.A2(n_1121),
.B1(n_1125),
.B2(n_1119),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1151),
.A2(n_1122),
.B(n_1149),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1157),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1198),
.B(n_1237),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1182),
.B(n_1135),
.Y(n_1278)
);

BUFx2_ASAP7_75t_R g1279 ( 
.A(n_1212),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1199),
.Y(n_1280)
);

CKINVDCx12_ASAP7_75t_R g1281 ( 
.A(n_1192),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1199),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1236),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1121),
.B(n_1125),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1160),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1209),
.A2(n_1232),
.B(n_1251),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1173),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1149),
.A2(n_1131),
.B(n_1129),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1159),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1220),
.B(n_1228),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1119),
.B(n_1116),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1116),
.B(n_1191),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1155),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1248),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1134),
.A2(n_1242),
.B(n_1222),
.Y(n_1295)
);

AO21x1_ASAP7_75t_L g1296 ( 
.A1(n_1188),
.A2(n_1238),
.B(n_1158),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1136),
.A2(n_1141),
.B(n_1143),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1154),
.B(n_1145),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1188),
.A2(n_1148),
.B1(n_1211),
.B2(n_1196),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1148),
.A2(n_1217),
.B1(n_1203),
.B2(n_1211),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1153),
.B(n_1201),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1159),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1127),
.A2(n_1137),
.B(n_1165),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1154),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1152),
.A2(n_1234),
.A3(n_1226),
.B(n_1203),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1168),
.A2(n_1226),
.B(n_1217),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1215),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1213),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1169),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1156),
.A2(n_1230),
.B(n_1219),
.Y(n_1311)
);

AND2x6_ASAP7_75t_L g1312 ( 
.A(n_1138),
.B(n_1140),
.Y(n_1312)
);

CKINVDCx11_ASAP7_75t_R g1313 ( 
.A(n_1166),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1189),
.A2(n_1230),
.B(n_1219),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1214),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1158),
.C(n_1250),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1135),
.B(n_1201),
.Y(n_1317)
);

AOI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1150),
.A2(n_1189),
.B(n_1161),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1193),
.A2(n_1174),
.B(n_1133),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1170),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1205),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_SL g1322 ( 
.A1(n_1150),
.A2(n_1178),
.B(n_1179),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1164),
.A2(n_1175),
.B(n_1147),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1176),
.B(n_1130),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1193),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1124),
.A2(n_1253),
.B(n_1239),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1231),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1193),
.A2(n_1133),
.B(n_1139),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1180),
.B(n_1179),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1205),
.A2(n_1239),
.B(n_1176),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1181),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1162),
.A2(n_1233),
.B1(n_1199),
.B2(n_1213),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1177),
.A2(n_1172),
.B(n_1130),
.Y(n_1333)
);

AND2x4_ASAP7_75t_SL g1334 ( 
.A(n_1233),
.B(n_1185),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1245),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1130),
.B(n_1233),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1177),
.A2(n_1120),
.B(n_1114),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1186),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1187),
.A2(n_1117),
.B(n_1142),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1126),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1128),
.B(n_1198),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1120),
.A2(n_1114),
.B(n_1113),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1115),
.A2(n_1194),
.B(n_1123),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1128),
.A2(n_612),
.B(n_1246),
.C(n_1094),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1204),
.A2(n_1142),
.B(n_1206),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1126),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1126),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1236),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1120),
.A2(n_1114),
.B(n_1113),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1236),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1187),
.B(n_1183),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1215),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1115),
.A2(n_1194),
.B(n_1123),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1236),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1126),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1192),
.B(n_1228),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1236),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1126),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1204),
.A2(n_1142),
.B(n_1206),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1204),
.A2(n_1142),
.B(n_1206),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1243),
.B(n_1010),
.Y(n_1361)
);

AO221x2_ASAP7_75t_L g1362 ( 
.A1(n_1246),
.A2(n_1240),
.B1(n_1190),
.B2(n_935),
.C(n_777),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1236),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1128),
.A2(n_612),
.B(n_1246),
.C(n_1094),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1190),
.A2(n_981),
.B1(n_883),
.B2(n_1240),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1190),
.A2(n_981),
.B1(n_883),
.B2(n_1240),
.Y(n_1366)
);

INVx2_ASAP7_75t_R g1367 ( 
.A(n_1187),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1184),
.B(n_1086),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_SL g1369 ( 
.A(n_1246),
.B(n_848),
.C(n_462),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1128),
.B(n_1198),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1208),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1126),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1128),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_1215),
.Y(n_1374)
);

NAND2x1_ASAP7_75t_L g1375 ( 
.A(n_1124),
.B(n_1253),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1246),
.A2(n_848),
.B(n_883),
.C(n_1146),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1126),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1126),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1236),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1243),
.B(n_1010),
.Y(n_1380)
);

AOI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_1190),
.A2(n_883),
.B(n_1101),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1126),
.Y(n_1382)
);

INVx5_ASAP7_75t_L g1383 ( 
.A(n_1199),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1337),
.A2(n_1314),
.B(n_1311),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1356),
.B(n_1294),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1298),
.B(n_1316),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1287),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1316),
.B(n_1348),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1341),
.A2(n_1370),
.B1(n_1373),
.B2(n_1365),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1320),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1309),
.Y(n_1391)
);

OA22x2_ASAP7_75t_L g1392 ( 
.A1(n_1269),
.A2(n_1261),
.B1(n_1305),
.B2(n_1277),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1292),
.B(n_1299),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1337),
.A2(n_1314),
.B(n_1311),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1319),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1274),
.A2(n_1364),
.B(n_1344),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1265),
.A2(n_1353),
.B(n_1343),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1350),
.B(n_1264),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1291),
.B(n_1284),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1309),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1304),
.A2(n_1297),
.B(n_1310),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1290),
.B(n_1361),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1283),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1301),
.B(n_1289),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1301),
.B(n_1303),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1327),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1380),
.B(n_1264),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1300),
.B(n_1354),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1300),
.B(n_1357),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1366),
.A2(n_1344),
.B1(n_1364),
.B2(n_1315),
.Y(n_1411)
);

O2A1O1Ixp5_ASAP7_75t_L g1412 ( 
.A1(n_1296),
.A2(n_1275),
.B(n_1381),
.C(n_1288),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1379),
.B(n_1363),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1329),
.B(n_1302),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1259),
.Y(n_1415)
);

O2A1O1Ixp5_ASAP7_75t_L g1416 ( 
.A1(n_1325),
.A2(n_1318),
.B(n_1293),
.C(n_1331),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1315),
.A2(n_1329),
.B1(n_1255),
.B2(n_1376),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1276),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1319),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1312),
.B(n_1346),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1362),
.B(n_1368),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1312),
.B(n_1347),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1369),
.A2(n_1362),
.B(n_1332),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1319),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1362),
.A2(n_1345),
.B(n_1359),
.Y(n_1425)
);

NAND2x1_ASAP7_75t_L g1426 ( 
.A(n_1351),
.B(n_1322),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1338),
.A2(n_1317),
.B1(n_1334),
.B2(n_1335),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1368),
.B(n_1355),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1345),
.A2(n_1359),
.B(n_1360),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_SL g1430 ( 
.A1(n_1266),
.A2(n_1257),
.B(n_1278),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1368),
.B(n_1355),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1312),
.B(n_1358),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1306),
.B(n_1378),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1378),
.B(n_1382),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1260),
.A2(n_1339),
.B(n_1285),
.C(n_1377),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1281),
.B(n_1259),
.Y(n_1436)
);

O2A1O1Ixp5_ASAP7_75t_L g1437 ( 
.A1(n_1325),
.A2(n_1293),
.B(n_1258),
.C(n_1268),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1271),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1254),
.B(n_1267),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1312),
.B(n_1340),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1260),
.A2(n_1372),
.B(n_1262),
.C(n_1351),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1312),
.B(n_1306),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1334),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1321),
.B(n_1383),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1327),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1307),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1321),
.B(n_1336),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1324),
.A2(n_1367),
.B(n_1258),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1351),
.A2(n_1360),
.B1(n_1279),
.B2(n_1383),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1313),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1333),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1328),
.A2(n_1367),
.B(n_1371),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1383),
.A2(n_1321),
.B1(n_1371),
.B2(n_1375),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_SL g1454 ( 
.A(n_1352),
.Y(n_1454)
);

O2A1O1Ixp5_ASAP7_75t_L g1455 ( 
.A1(n_1293),
.A2(n_1258),
.B(n_1273),
.C(n_1272),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1328),
.A2(n_1281),
.B(n_1295),
.C(n_1272),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1280),
.B(n_1282),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1295),
.A2(n_1323),
.B(n_1313),
.C(n_1333),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1280),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1280),
.A2(n_1282),
.B(n_1308),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1330),
.A2(n_1326),
.B(n_1286),
.C(n_1342),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1383),
.A2(n_1263),
.B1(n_1282),
.B2(n_1308),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1282),
.B(n_1270),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1330),
.B(n_1270),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1256),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1256),
.B(n_1349),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1374),
.A2(n_1128),
.B(n_1373),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1356),
.B(n_1294),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1356),
.B(n_1294),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1373),
.B(n_1341),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1373),
.B(n_1341),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1464),
.B(n_1429),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1384),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1426),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1395),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1394),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1419),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1394),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1419),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1411),
.A2(n_1410),
.B1(n_1389),
.B2(n_1417),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1401),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1424),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1404),
.B(n_1405),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1396),
.B(n_1397),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1451),
.B(n_1425),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1442),
.B(n_1433),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1437),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1465),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1466),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1463),
.B(n_1438),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1392),
.B(n_1386),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1448),
.A2(n_1412),
.B(n_1416),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1456),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1418),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1392),
.A2(n_1471),
.B1(n_1470),
.B2(n_1402),
.Y(n_1497)
);

AO21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1420),
.A2(n_1432),
.B(n_1422),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1440),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1435),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1452),
.B(n_1408),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1441),
.B(n_1467),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1393),
.B(n_1399),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1439),
.A2(n_1388),
.B(n_1409),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1407),
.B(n_1414),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1458),
.B(n_1421),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1387),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1458),
.B(n_1434),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1449),
.A2(n_1390),
.B(n_1431),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1398),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1423),
.B(n_1428),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1475),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1484),
.B(n_1385),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1476),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1494),
.A2(n_1444),
.B(n_1427),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1474),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.Y(n_1519)
);

OR2x2_ASAP7_75t_SL g1520 ( 
.A(n_1505),
.B(n_1469),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1487),
.B(n_1468),
.Y(n_1521)
);

AOI222xp33_ASAP7_75t_L g1522 ( 
.A1(n_1481),
.A2(n_1454),
.B1(n_1450),
.B2(n_1406),
.C1(n_1436),
.C2(n_1445),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1403),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1487),
.B(n_1413),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1484),
.B(n_1459),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1473),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1487),
.B(n_1453),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1457),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1473),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1473),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1479),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1483),
.B(n_1462),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1483),
.B(n_1443),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1484),
.B(n_1391),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1490),
.B(n_1430),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1498),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1496),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1511),
.B(n_1508),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1496),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1537),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1515),
.A2(n_1493),
.B1(n_1481),
.B2(n_1497),
.C(n_1500),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1524),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1537),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1526),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1515),
.A2(n_1493),
.B1(n_1497),
.B2(n_1500),
.C(n_1495),
.Y(n_1546)
);

OAI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1522),
.A2(n_1485),
.B1(n_1503),
.B2(n_1500),
.C(n_1512),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_R g1548 ( 
.A(n_1534),
.B(n_1415),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1526),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1518),
.A2(n_1488),
.B(n_1492),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1513),
.A2(n_1485),
.B1(n_1507),
.B2(n_1500),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1521),
.A2(n_1503),
.B1(n_1485),
.B2(n_1512),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1518),
.A2(n_1488),
.B(n_1477),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1503),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1539),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1525),
.B(n_1511),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1539),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1519),
.A2(n_1492),
.B(n_1482),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1527),
.A2(n_1485),
.B1(n_1502),
.B2(n_1512),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1522),
.A2(n_1485),
.B1(n_1507),
.B2(n_1509),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1514),
.B(n_1472),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1519),
.A2(n_1492),
.B(n_1482),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1514),
.B(n_1472),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1520),
.B(n_1538),
.Y(n_1564)
);

OAI33xp33_ASAP7_75t_L g1565 ( 
.A1(n_1524),
.A2(n_1504),
.A3(n_1495),
.B1(n_1491),
.B2(n_1478),
.B3(n_1480),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1538),
.A2(n_1485),
.B(n_1460),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1511),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1529),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1525),
.B(n_1499),
.Y(n_1571)
);

NAND4xp25_ASAP7_75t_SL g1572 ( 
.A(n_1527),
.B(n_1507),
.C(n_1502),
.D(n_1504),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1536),
.A2(n_1495),
.B1(n_1504),
.B2(n_1507),
.C(n_1501),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1517),
.B(n_1505),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1514),
.B(n_1472),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1520),
.A2(n_1485),
.B1(n_1502),
.B2(n_1510),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1530),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1540),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1545),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1542),
.B(n_1485),
.C(n_1501),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1546),
.B(n_1536),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1545),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1561),
.B(n_1531),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1569),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1523),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1570),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1554),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1516),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1531),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1556),
.B(n_1523),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1558),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1576),
.A2(n_1485),
.B(n_1501),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1573),
.B(n_1523),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1574),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1541),
.B(n_1544),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1577),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1563),
.B(n_1531),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1550),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1550),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1531),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1551),
.B(n_1560),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1555),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1584),
.B(n_1563),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1588),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1590),
.B(n_1564),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1581),
.B(n_1548),
.C(n_1547),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1584),
.B(n_1575),
.Y(n_1613)
);

NOR3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1581),
.B(n_1552),
.C(n_1572),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1588),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1575),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1591),
.B(n_1568),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

CKINVDCx16_ASAP7_75t_R g1619 ( 
.A(n_1589),
.Y(n_1619)
);

AND2x2_ASAP7_75t_SL g1620 ( 
.A(n_1595),
.B(n_1505),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1582),
.B(n_1595),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1568),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1605),
.B(n_1566),
.C(n_1531),
.Y(n_1623)
);

INVxp67_ASAP7_75t_SL g1624 ( 
.A(n_1582),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1589),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1608),
.B(n_1557),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1579),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1591),
.B(n_1513),
.Y(n_1629)
);

OAI31xp33_ASAP7_75t_L g1630 ( 
.A1(n_1605),
.A2(n_1559),
.A3(n_1502),
.B(n_1486),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1579),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1608),
.B(n_1578),
.Y(n_1632)
);

AOI221x1_ASAP7_75t_L g1633 ( 
.A1(n_1594),
.A2(n_1400),
.B1(n_1567),
.B2(n_1571),
.C(n_1489),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1513),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1583),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1580),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1594),
.B(n_1521),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1580),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1586),
.Y(n_1640)
);

OAI33xp33_ASAP7_75t_L g1641 ( 
.A1(n_1590),
.A2(n_1524),
.A3(n_1521),
.B1(n_1533),
.B2(n_1491),
.B3(n_1528),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1587),
.B(n_1528),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1586),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1579),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1587),
.B(n_1528),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1585),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1585),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1597),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1580),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1592),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1619),
.B(n_1592),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1625),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1627),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1619),
.B(n_1597),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1506),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1629),
.B(n_1600),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1612),
.A2(n_1603),
.B(n_1601),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1631),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1625),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1631),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1618),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1618),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1618),
.Y(n_1664)
);

OAI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1623),
.A2(n_1527),
.B1(n_1607),
.B2(n_1532),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1644),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1611),
.B(n_1608),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1635),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1644),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1614),
.B(n_1506),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1648),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1640),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1646),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1646),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1630),
.B(n_1506),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1611),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1647),
.Y(n_1678)
);

NAND2x1p5_ASAP7_75t_L g1679 ( 
.A(n_1638),
.B(n_1505),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1647),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1620),
.B(n_1506),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1610),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1600),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1668),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1652),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1660),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1677),
.B(n_1622),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1656),
.B(n_1609),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1679),
.A2(n_1615),
.B(n_1610),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1656),
.B(n_1620),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1683),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1623),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1651),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1622),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1673),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1653),
.Y(n_1698)
);

NOR2xp67_ASAP7_75t_SL g1699 ( 
.A(n_1672),
.B(n_1400),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1658),
.A2(n_1620),
.B1(n_1642),
.B2(n_1645),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1683),
.B(n_1609),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1657),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1667),
.B(n_1676),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1667),
.Y(n_1704)
);

NOR2x1_ASAP7_75t_L g1705 ( 
.A(n_1682),
.B(n_1615),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1658),
.A2(n_1641),
.B1(n_1607),
.B2(n_1565),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1684),
.B(n_1634),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1662),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1657),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1697),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1670),
.Y(n_1711)
);

AOI222xp33_ASAP7_75t_L g1712 ( 
.A1(n_1700),
.A2(n_1665),
.B1(n_1681),
.B2(n_1682),
.C1(n_1655),
.C2(n_1607),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1685),
.B(n_1613),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1693),
.A2(n_1699),
.B1(n_1694),
.B2(n_1697),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1688),
.B(n_1642),
.Y(n_1715)
);

AOI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1686),
.A2(n_1679),
.B1(n_1680),
.B2(n_1678),
.C(n_1675),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1705),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1707),
.B(n_1679),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1704),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1686),
.B(n_1659),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_L g1723 ( 
.A(n_1699),
.B(n_1633),
.C(n_1659),
.Y(n_1723)
);

OAI322xp33_ASAP7_75t_L g1724 ( 
.A1(n_1685),
.A2(n_1680),
.A3(n_1678),
.B1(n_1675),
.B2(n_1674),
.C1(n_1661),
.C2(n_1669),
.Y(n_1724)
);

OAI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1706),
.A2(n_1596),
.B1(n_1669),
.B2(n_1674),
.C(n_1666),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1690),
.A2(n_1633),
.B(n_1661),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1689),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1692),
.B(n_1613),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1725),
.A2(n_1712),
.B1(n_1711),
.B2(n_1717),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1722),
.Y(n_1730)
);

OR3x1_ASAP7_75t_L g1731 ( 
.A(n_1710),
.B(n_1698),
.C(n_1695),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1720),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1713),
.B(n_1692),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1719),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1721),
.B(n_1701),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1727),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1724),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1714),
.B(n_1688),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1713),
.B(n_1701),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1737),
.A2(n_1714),
.B1(n_1728),
.B2(n_1723),
.Y(n_1740)
);

NOR3xp33_ASAP7_75t_L g1741 ( 
.A(n_1738),
.B(n_1724),
.C(n_1716),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1738),
.A2(n_1726),
.B(n_1718),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1730),
.A2(n_1735),
.B(n_1736),
.C(n_1734),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1739),
.A2(n_1704),
.B(n_1715),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1733),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1729),
.B(n_1691),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1731),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1729),
.A2(n_1732),
.B1(n_1709),
.B2(n_1702),
.C(n_1698),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1738),
.A2(n_1696),
.B1(n_1703),
.B2(n_1691),
.C(n_1702),
.Y(n_1749)
);

AOI222xp33_ASAP7_75t_L g1750 ( 
.A1(n_1746),
.A2(n_1709),
.B1(n_1695),
.B2(n_1690),
.C1(n_1708),
.C2(n_1666),
.Y(n_1750)
);

AOI322xp5_ASAP7_75t_L g1751 ( 
.A1(n_1741),
.A2(n_1601),
.A3(n_1603),
.B1(n_1708),
.B2(n_1602),
.C1(n_1606),
.C2(n_1593),
.Y(n_1751)
);

AO22x1_ASAP7_75t_L g1752 ( 
.A1(n_1747),
.A2(n_1664),
.B1(n_1663),
.B2(n_1671),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1745),
.Y(n_1753)
);

AOI222xp33_ASAP7_75t_L g1754 ( 
.A1(n_1748),
.A2(n_1671),
.B1(n_1664),
.B2(n_1663),
.C1(n_1662),
.C2(n_1637),
.Y(n_1754)
);

AO22x2_ASAP7_75t_L g1755 ( 
.A1(n_1742),
.A2(n_1696),
.B1(n_1703),
.B2(n_1649),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1755),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1753),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1750),
.B(n_1744),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1752),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1754),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1751),
.B(n_1749),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1740),
.B1(n_1743),
.B2(n_1636),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1758),
.A2(n_1604),
.B(n_1649),
.C(n_1639),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1756),
.B(n_1760),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1757),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1759),
.A2(n_1617),
.B(n_1649),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1762),
.B(n_1759),
.C(n_1639),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1764),
.B(n_1645),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1765),
.B(n_1639),
.C(n_1637),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1767),
.B(n_1763),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1770),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1768),
.B1(n_1766),
.B2(n_1769),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1771),
.B(n_1596),
.C(n_1617),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1772),
.A2(n_1626),
.B(n_1632),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1773),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1628),
.B1(n_1636),
.B2(n_1634),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1774),
.A2(n_1636),
.B1(n_1628),
.B2(n_1607),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1636),
.B1(n_1628),
.B2(n_1596),
.Y(n_1778)
);

OAI222xp33_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1776),
.B1(n_1596),
.B2(n_1602),
.C1(n_1593),
.C2(n_1606),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1779),
.B(n_1616),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_R g1781 ( 
.A1(n_1780),
.A2(n_1628),
.B1(n_1598),
.B2(n_1586),
.C(n_1602),
.Y(n_1781)
);

AOI31xp33_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1626),
.A3(n_1632),
.B(n_1616),
.Y(n_1782)
);

AOI211xp5_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_1606),
.B(n_1593),
.C(n_1599),
.Y(n_1783)
);


endmodule