module fake_jpeg_12358_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_0),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_57),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_86),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_91),
.B1(n_57),
.B2(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_52),
.B1(n_64),
.B2(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_70),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_77),
.B1(n_64),
.B2(n_60),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_72),
.B1(n_71),
.B2(n_74),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_1),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_113),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_79),
.C(n_59),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_114),
.Y(n_144)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_78),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_74),
.B1(n_60),
.B2(n_54),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_124),
.B1(n_63),
.B2(n_2),
.Y(n_127)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_65),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_66),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_126),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_15),
.B1(n_17),
.B2(n_21),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_137),
.Y(n_155)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_6),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_26),
.B(n_27),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_146),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_151),
.B1(n_161),
.B2(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_156),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_140),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_164),
.C(n_165),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_132),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_142),
.B(n_29),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B(n_173),
.C(n_37),
.D(n_42),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_28),
.C(n_31),
.Y(n_171)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_180),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_160),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_182),
.C(n_176),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_163),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_166),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_179),
.C(n_181),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_174),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_190),
.A2(n_174),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_47),
.Y(n_193)
);


endmodule