module fake_jpeg_19392_n_377 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_377);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_377;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_54),
.B(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_68),
.Y(n_101)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_8),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_70),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_25),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_84),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_87),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_44),
.B1(n_25),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_88),
.A2(n_92),
.B1(n_109),
.B2(n_112),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_25),
.B1(n_42),
.B2(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_100),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_57),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_49),
.B(n_34),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_39),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_39),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_120),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_52),
.B(n_21),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_47),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_20),
.B1(n_26),
.B2(n_41),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_50),
.B1(n_63),
.B2(n_60),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_38),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_38),
.C(n_20),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_132),
.B(n_71),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_66),
.A2(n_20),
.B1(n_26),
.B2(n_41),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_28),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_133),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_43),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_78),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_26),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_166),
.Y(n_184)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g139 ( 
.A(n_89),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_141),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_27),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_142),
.A2(n_89),
.B(n_113),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_144),
.B(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_147),
.A2(n_155),
.B1(n_159),
.B2(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_84),
.A2(n_53),
.B1(n_73),
.B2(n_27),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_149),
.A2(n_150),
.B1(n_157),
.B2(n_161),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_72),
.B1(n_58),
.B2(n_43),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_128),
.B1(n_83),
.B2(n_93),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_110),
.B1(n_127),
.B2(n_111),
.Y(n_180)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_156),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_28),
.B1(n_35),
.B2(n_42),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_71),
.B1(n_9),
.B2(n_10),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_106),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_2),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_82),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_88),
.A2(n_7),
.B1(n_11),
.B2(n_13),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_175),
.B1(n_132),
.B2(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_172),
.Y(n_185)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_90),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_11),
.B1(n_16),
.B2(n_6),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_117),
.A2(n_16),
.B1(n_2),
.B2(n_4),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_116),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_180),
.A2(n_182),
.B1(n_187),
.B2(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_140),
.B1(n_163),
.B2(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_132),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_211),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_127),
.B1(n_97),
.B2(n_124),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_157),
.C(n_150),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_197),
.B1(n_207),
.B2(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_166),
.B1(n_161),
.B2(n_142),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_97),
.B1(n_91),
.B2(n_117),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_144),
.B(n_94),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_206),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_138),
.A2(n_129),
.B1(n_95),
.B2(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_104),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_160),
.A2(n_85),
.B(n_4),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_96),
.B1(n_122),
.B2(n_119),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_228),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_143),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_220),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_152),
.B1(n_172),
.B2(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_134),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_152),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_135),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_226),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_195),
.A2(n_141),
.B1(n_135),
.B2(n_162),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_122),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_151),
.B1(n_156),
.B2(n_171),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_192),
.B1(n_180),
.B2(n_200),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_137),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_231),
.B(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_158),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_153),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_123),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_123),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_113),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_119),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_208),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_192),
.B(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_220),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_266),
.B1(n_219),
.B2(n_226),
.Y(n_279)
);

NOR4xp25_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_209),
.C(n_193),
.D(n_212),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_236),
.B(n_193),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_203),
.C(n_202),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_271),
.C(n_217),
.Y(n_283)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_234),
.B1(n_223),
.B2(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_270),
.B(n_238),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_198),
.C(n_178),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_249),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_284),
.B(n_263),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_231),
.B1(n_243),
.B2(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_286),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_218),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_280),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_219),
.B1(n_230),
.B2(n_210),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_210),
.B1(n_222),
.B2(n_196),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_289),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_216),
.B(n_233),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_216),
.C(n_228),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_255),
.C(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_227),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_293),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_245),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_290),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_248),
.A2(n_246),
.B1(n_242),
.B2(n_240),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_250),
.B1(n_259),
.B2(n_269),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_251),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_215),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_250),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_215),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_269),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_301),
.C(n_302),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_298),
.A2(n_287),
.B1(n_279),
.B2(n_291),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_255),
.C(n_258),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_258),
.C(n_264),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_247),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_286),
.B(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_247),
.C(n_272),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_303),
.C(n_301),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_254),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_324),
.B(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_326),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_312),
.C(n_300),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_297),
.A2(n_284),
.B1(n_293),
.B2(n_280),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_322),
.A2(n_328),
.B1(n_309),
.B2(n_306),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_290),
.C(n_247),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_329),
.Y(n_332)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

AOI321xp33_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_292),
.A3(n_288),
.B1(n_281),
.B2(n_273),
.C(n_253),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_330),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_299),
.A2(n_292),
.B1(n_288),
.B2(n_281),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_273),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_319),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_334),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_337),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_302),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_317),
.A2(n_323),
.B1(n_315),
.B2(n_318),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_241),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_340),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_322),
.A2(n_314),
.B1(n_296),
.B2(n_306),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_313),
.C(n_314),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_342),
.B(n_343),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_254),
.C(n_267),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_328),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_354),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_335),
.A2(n_270),
.B1(n_260),
.B2(n_265),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_348),
.A2(n_353),
.B1(n_338),
.B2(n_201),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_316),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_352),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_331),
.A2(n_316),
.B(n_261),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_351),
.B(n_343),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_260),
.B1(n_253),
.B2(n_251),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_239),
.B1(n_235),
.B2(n_200),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_356),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_337),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_358),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_347),
.A2(n_200),
.B1(n_205),
.B2(n_201),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_359),
.A2(n_360),
.B(n_362),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_346),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_342),
.Y(n_363)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_344),
.C(n_349),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_366),
.A2(n_368),
.B(n_369),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_336),
.C(n_352),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_350),
.C(n_181),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_361),
.C(n_359),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_370),
.B(n_372),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_364),
.B(n_205),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_188),
.C(n_185),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_191),
.B(n_188),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_371),
.B(n_191),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_376),
.B(n_375),
.Y(n_377)
);


endmodule