module fake_netlist_6_4883_n_1972 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_44, n_1972);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_44;

output n_1972;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_68;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_77;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_78;
wire n_1380;
wire n_442;
wire n_480;
wire n_142;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_62;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_65;
wire n_230;
wire n_461;
wire n_873;
wire n_141;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_71;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_112;
wire n_1280;
wire n_713;
wire n_1400;
wire n_126;
wire n_1467;
wire n_58;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_166;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_92;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_102;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_121;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_61;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_117;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_134;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_136;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_88;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_55;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_91;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_63;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_125;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_131;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_59;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_108;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_86;
wire n_104;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_72;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_79;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_147;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_118;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_107;
wire n_1228;
wire n_417;
wire n_446;
wire n_89;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_69;
wire n_293;
wire n_53;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_98;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_66;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_100;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_124;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_123;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_128;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_146;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_113;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_90;
wire n_54;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_99;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_120;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_106;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_140;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_67;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_73;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_101;
wire n_167;
wire n_1356;
wire n_1589;
wire n_127;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_133;
wire n_1320;
wire n_96;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_137;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_122;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_70;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_97;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_80;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_83;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_105;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_76;
wire n_548;
wire n_1782;
wire n_94;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_139;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_138;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_85;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_75;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_110;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_57;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_52;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_84;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_114;
wire n_300;
wire n_222;
wire n_747;
wire n_74;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_111;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1785;
wire n_1848;
wire n_56;
wire n_763;
wire n_1114;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_119;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_129;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_109;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_82;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_93;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_103;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_132;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_130;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_116;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_95;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_115;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_87;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_81;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_64;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_135;
wire n_165;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_60;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_51;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

BUFx2_ASAP7_75t_R g74 ( 
.A(n_9),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_13),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_26),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_3),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_31),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_31),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_7),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_4),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_36),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_77),
.B(n_92),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_68),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_100),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVxp33_ASAP7_75t_SL g138 ( 
.A(n_120),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_57),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_57),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_112),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_112),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_67),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_136),
.B(n_134),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_R g167 ( 
.A(n_139),
.B(n_115),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_R g168 ( 
.A(n_137),
.B(n_115),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_113),
.Y(n_176)
);

AO21x2_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_145),
.B(n_149),
.Y(n_177)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_137),
.B(n_68),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_139),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_R g189 ( 
.A(n_147),
.B(n_106),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_113),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_147),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

CKINVDCx6p67_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_145),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_145),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_145),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_126),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_146),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_R g215 ( 
.A(n_135),
.B(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_126),
.B1(n_131),
.B2(n_146),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_67),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_110),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

AND3x4_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_74),
.C(n_65),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_110),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_119),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_119),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_126),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_91),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_177),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_167),
.B(n_135),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_152),
.B(n_70),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_153),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_157),
.B(n_186),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_157),
.B(n_150),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_156),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_177),
.B(n_126),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_157),
.B(n_150),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_167),
.B(n_135),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_126),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_160),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_157),
.B(n_150),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g260 ( 
.A(n_213),
.Y(n_260)
);

CKINVDCx6p67_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_157),
.B(n_150),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_215),
.B(n_178),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_159),
.B(n_91),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_215),
.B(n_135),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_150),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_131),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_163),
.B(n_126),
.C(n_136),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_168),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_159),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_161),
.B(n_70),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_162),
.B(n_126),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_173),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_187),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_187),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_166),
.B(n_131),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_198),
.B(n_187),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_182),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_198),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_182),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_204),
.A2(n_126),
.B1(n_131),
.B2(n_146),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_186),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_212),
.B(n_164),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_173),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_212),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_155),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_186),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_155),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_214),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_176),
.A2(n_77),
.B(n_75),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_189),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_191),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_186),
.B(n_150),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_176),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_192),
.B(n_131),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_191),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_216),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_158),
.B(n_108),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_192),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_170),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_164),
.B(n_131),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_192),
.B(n_131),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_192),
.Y(n_318)
);

OR2x6_ASAP7_75t_L g319 ( 
.A(n_158),
.B(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_197),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_183),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_197),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g323 ( 
.A(n_197),
.B(n_131),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_197),
.B(n_131),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_197),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_171),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_179),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_220),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_224),
.B(n_185),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_254),
.B(n_68),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_180),
.Y(n_332)
);

AOI221xp5_ASAP7_75t_L g333 ( 
.A1(n_238),
.A2(n_56),
.B1(n_66),
.B2(n_75),
.C(n_80),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_220),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_265),
.A2(n_195),
.B1(n_188),
.B2(n_254),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_184),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_190),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_194),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_233),
.A2(n_131),
.B1(n_146),
.B2(n_149),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_220),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_196),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_150),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_271),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_287),
.A2(n_131),
.B1(n_146),
.B2(n_100),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_227),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_254),
.A2(n_65),
.B1(n_135),
.B2(n_100),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_227),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_SL g351 ( 
.A(n_254),
.B(n_66),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_150),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_254),
.B(n_135),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_287),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_287),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_287),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_122),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_260),
.B(n_135),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_291),
.B(n_134),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_291),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_289),
.A2(n_131),
.B1(n_146),
.B2(n_100),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_227),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_288),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_260),
.B(n_135),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_272),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_291),
.B(n_134),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_298),
.B(n_134),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_134),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_223),
.B(n_53),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_226),
.B(n_54),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_298),
.B(n_134),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_260),
.B(n_135),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_217),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_272),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_217),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_219),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_273),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_273),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_219),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_311),
.B(n_148),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_233),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_276),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_298),
.B(n_148),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_222),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_260),
.B(n_135),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_228),
.B(n_55),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_222),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_230),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_281),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_224),
.B(n_77),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_281),
.A2(n_149),
.B(n_148),
.C(n_136),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_279),
.B(n_148),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_236),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_279),
.B(n_148),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_283),
.B(n_149),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_283),
.B(n_149),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_233),
.A2(n_146),
.B1(n_144),
.B2(n_141),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_267),
.A2(n_121),
.B(n_124),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_L g401 ( 
.A(n_295),
.B(n_100),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_292),
.B(n_141),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_292),
.B(n_141),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_289),
.B(n_141),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_236),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_233),
.A2(n_146),
.B1(n_144),
.B2(n_141),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_289),
.B(n_141),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_221),
.B(n_58),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_289),
.B(n_141),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_237),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_278),
.A2(n_234),
.B1(n_232),
.B2(n_312),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_282),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_260),
.B(n_135),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_232),
.B(n_141),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_310),
.B(n_144),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_310),
.B(n_144),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_224),
.B(n_135),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_224),
.B(n_253),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_295),
.B(n_80),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_296),
.A2(n_146),
.B1(n_144),
.B2(n_113),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_237),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_239),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_296),
.A2(n_146),
.B1(n_144),
.B2(n_114),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_253),
.B(n_121),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_255),
.B(n_59),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_253),
.B(n_121),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_312),
.B(n_60),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_234),
.B(n_144),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_239),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_346),
.B(n_240),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_342),
.B(n_427),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_368),
.B(n_253),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_368),
.B(n_302),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_247),
.B(n_241),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_392),
.A2(n_242),
.B(n_267),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_302),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_369),
.B(n_278),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

OR2x6_ASAP7_75t_L g440 ( 
.A(n_354),
.B(n_305),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_389),
.B(n_297),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_411),
.A2(n_320),
.B(n_317),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_370),
.B(n_313),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_408),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_392),
.A2(n_267),
.B(n_318),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_338),
.B(n_313),
.Y(n_446)
);

CKINVDCx8_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_393),
.A2(n_275),
.B(n_246),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_304),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_267),
.B(n_318),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_339),
.B(n_313),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_390),
.B(n_322),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_360),
.B(n_322),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_318),
.B(n_325),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_363),
.A2(n_318),
.B(n_325),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_360),
.B(n_322),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_363),
.A2(n_325),
.B(n_248),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_326),
.A2(n_296),
.B1(n_295),
.B2(n_317),
.Y(n_460)
);

O2A1O1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_411),
.A2(n_327),
.B(n_337),
.C(n_263),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_330),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_368),
.B(n_302),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_231),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_332),
.B(n_231),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_330),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_420),
.A2(n_275),
.B(n_251),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_363),
.A2(n_257),
.B(n_243),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_425),
.B(n_244),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_391),
.B(n_302),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g472 ( 
.A1(n_404),
.A2(n_320),
.B(n_407),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_335),
.B(n_305),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_354),
.B(n_321),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_330),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_366),
.B(n_246),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_363),
.A2(n_270),
.B(n_262),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_355),
.B(n_245),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_375),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_363),
.A2(n_307),
.B(n_424),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_330),
.Y(n_481)
);

BUFx4f_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_366),
.B(n_251),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_329),
.B(n_261),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_355),
.B(n_268),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_363),
.A2(n_295),
.B(n_269),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_356),
.A2(n_295),
.B1(n_381),
.B2(n_368),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_426),
.A2(n_295),
.B(n_300),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_333),
.A2(n_303),
.B(n_268),
.C(n_247),
.Y(n_490)
);

O2A1O1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_365),
.A2(n_303),
.B(n_256),
.C(n_241),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_336),
.B(n_245),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_L g493 ( 
.A1(n_345),
.A2(n_218),
.B(n_294),
.Y(n_493)
);

BUFx12f_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_428),
.A2(n_300),
.B(n_235),
.Y(n_495)
);

BUFx12f_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_376),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_409),
.A2(n_300),
.B(n_250),
.Y(n_498)
);

INVx11_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

O2A1O1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_365),
.A2(n_266),
.B(n_252),
.C(n_256),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_356),
.B(n_261),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_336),
.B(n_225),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_344),
.B(n_225),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_359),
.A2(n_300),
.B(n_264),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_344),
.B(n_245),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_359),
.A2(n_300),
.B(n_264),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_420),
.A2(n_324),
.B(n_316),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_357),
.A2(n_300),
.B(n_264),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_343),
.A2(n_264),
.B(n_316),
.Y(n_509)
);

A2O1A1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_374),
.A2(n_268),
.B(n_249),
.C(n_259),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_419),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_352),
.A2(n_264),
.B(n_324),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_423),
.A2(n_309),
.B(n_268),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_381),
.B(n_264),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_347),
.B(n_309),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_380),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_367),
.A2(n_319),
.B(n_323),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_347),
.B(n_225),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_381),
.B(n_229),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_380),
.B(n_249),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_395),
.B(n_252),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_381),
.A2(n_319),
.B1(n_323),
.B2(n_258),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_419),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_423),
.B(n_323),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_395),
.B(n_258),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_421),
.B(n_285),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_371),
.A2(n_319),
.B(n_290),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_422),
.B(n_259),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_329),
.B(n_285),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_396),
.B(n_398),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_L g533 ( 
.A1(n_374),
.A2(n_266),
.B(n_319),
.C(n_89),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_385),
.B(n_285),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_396),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_382),
.A2(n_274),
.B(n_319),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_348),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_384),
.A2(n_293),
.B(n_290),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_351),
.A2(n_284),
.B(n_286),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_417),
.A2(n_293),
.B(n_290),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_398),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_385),
.A2(n_429),
.B1(n_388),
.B2(n_405),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_382),
.A2(n_399),
.B(n_406),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_402),
.A2(n_293),
.B(n_290),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_403),
.A2(n_293),
.B(n_290),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_388),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_405),
.B(n_410),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_353),
.A2(n_293),
.B(n_290),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_R g549 ( 
.A(n_410),
.B(n_229),
.Y(n_549)
);

AO21x1_ASAP7_75t_L g550 ( 
.A1(n_401),
.A2(n_377),
.B(n_378),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_429),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_377),
.B(n_229),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_348),
.Y(n_553)
);

CKINVDCx10_ASAP7_75t_R g554 ( 
.A(n_340),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_416),
.A2(n_293),
.B(n_285),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_378),
.B(n_379),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_379),
.B(n_315),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_383),
.B(n_229),
.Y(n_558)
);

AO21x1_ASAP7_75t_L g559 ( 
.A1(n_383),
.A2(n_284),
.B(n_286),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_358),
.A2(n_285),
.B(n_121),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_546),
.Y(n_561)
);

AND3x1_ASAP7_75t_L g562 ( 
.A(n_502),
.B(n_87),
.C(n_92),
.Y(n_562)
);

O2A1O1Ixp33_ASAP7_75t_SL g563 ( 
.A1(n_444),
.A2(n_341),
.B(n_334),
.C(n_328),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_535),
.B(n_364),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_450),
.A2(n_413),
.B(n_372),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_431),
.A2(n_532),
.B1(n_438),
.B2(n_503),
.Y(n_566)
);

O2A1O1Ixp5_ASAP7_75t_L g567 ( 
.A1(n_442),
.A2(n_386),
.B(n_397),
.C(n_394),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_476),
.B(n_328),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_455),
.A2(n_445),
.B(n_443),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_434),
.Y(n_570)
);

NOR3xp33_ASAP7_75t_SL g571 ( 
.A(n_502),
.B(n_85),
.C(n_62),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_430),
.Y(n_572)
);

A2O1A1Ixp33_ASAP7_75t_L g573 ( 
.A1(n_513),
.A2(n_341),
.B(n_334),
.C(n_350),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_466),
.B(n_350),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_434),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_470),
.A2(n_315),
.B1(n_406),
.B2(n_399),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_454),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_436),
.A2(n_487),
.B(n_461),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_456),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_485),
.B(n_314),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_441),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_SL g582 ( 
.A1(n_490),
.A2(n_362),
.B(n_340),
.C(n_89),
.Y(n_582)
);

O2A1O1Ixp5_ASAP7_75t_L g583 ( 
.A1(n_550),
.A2(n_362),
.B(n_400),
.C(n_284),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_483),
.B(n_314),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_446),
.B(n_314),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_451),
.A2(n_517),
.B(n_528),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_457),
.A2(n_285),
.B(n_286),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_498),
.A2(n_349),
.B(n_121),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_508),
.A2(n_121),
.B(n_124),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_473),
.B(n_361),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_464),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_437),
.B(n_331),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_L g594 ( 
.A1(n_503),
.A2(n_76),
.B(n_63),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_441),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_518),
.A2(n_99),
.B(n_87),
.C(n_65),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_535),
.A2(n_314),
.B1(n_315),
.B2(n_78),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_518),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_456),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_495),
.A2(n_128),
.B(n_124),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_504),
.A2(n_128),
.B(n_124),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_465),
.B(n_315),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_535),
.B(n_315),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_552),
.B(n_315),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_474),
.Y(n_606)
);

O2A1O1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_531),
.A2(n_99),
.B(n_114),
.C(n_116),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_447),
.B(n_315),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_456),
.Y(n_609)
);

CKINVDCx14_ASAP7_75t_R g610 ( 
.A(n_474),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_541),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_549),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_439),
.Y(n_613)
);

OAI22x1_ASAP7_75t_SL g614 ( 
.A1(n_554),
.A2(n_73),
.B1(n_101),
.B2(n_98),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_541),
.B(n_315),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_541),
.B(n_331),
.Y(n_616)
);

AOI21x1_ASAP7_75t_L g617 ( 
.A1(n_472),
.A2(n_114),
.B(n_116),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_439),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_541),
.B(n_331),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_468),
.B(n_331),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_452),
.B(n_331),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_484),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_551),
.A2(n_552),
.B1(n_507),
.B2(n_547),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_558),
.B(n_331),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_484),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_61),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_506),
.A2(n_128),
.B(n_121),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_475),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_SL g629 ( 
.A(n_549),
.B(n_519),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_555),
.A2(n_331),
.B(n_144),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_475),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_460),
.B(n_100),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_437),
.B(n_274),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_440),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_497),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_469),
.A2(n_128),
.B(n_121),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_477),
.A2(n_128),
.B(n_121),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_462),
.B(n_140),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_437),
.B(n_274),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_478),
.B(n_274),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_524),
.A2(n_69),
.B1(n_97),
.B2(n_72),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_497),
.B(n_274),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_516),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_435),
.A2(n_116),
.B(n_118),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_490),
.A2(n_93),
.B(n_81),
.C(n_82),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_501),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_475),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_531),
.A2(n_118),
.B(n_79),
.C(n_94),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_516),
.B(n_274),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_459),
.A2(n_128),
.B(n_121),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_526),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_475),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_526),
.B(n_274),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_448),
.B(n_274),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_530),
.B(n_100),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_481),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_SL g658 ( 
.A1(n_533),
.A2(n_118),
.B(n_129),
.C(n_130),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_440),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_530),
.B(n_96),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_524),
.A2(n_433),
.B(n_463),
.C(n_510),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_520),
.B(n_288),
.Y(n_662)
);

CKINVDCx6p67_ASAP7_75t_R g663 ( 
.A(n_494),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_553),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_481),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_489),
.A2(n_124),
.B(n_121),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_553),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_521),
.B(n_288),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_537),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_432),
.A2(n_124),
.B(n_121),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_525),
.B(n_288),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_543),
.A2(n_100),
.B1(n_146),
.B2(n_84),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_493),
.A2(n_146),
.B1(n_83),
.B2(n_86),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_501),
.Y(n_675)
);

BUFx4f_ASAP7_75t_L g676 ( 
.A(n_481),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_449),
.B(n_90),
.C(n_95),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_SL g678 ( 
.A1(n_536),
.A2(n_480),
.B(n_540),
.C(n_548),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_433),
.A2(n_132),
.B(n_130),
.C(n_129),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_529),
.B(n_288),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_556),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_440),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_556),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_530),
.B(n_143),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_478),
.B(n_288),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_432),
.A2(n_121),
.B(n_124),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_542),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_557),
.B(n_143),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_478),
.B(n_288),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_481),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_486),
.A2(n_288),
.B1(n_143),
.B2(n_142),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_515),
.B(n_146),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_462),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_463),
.B(n_0),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_522),
.B(n_143),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_509),
.A2(n_121),
.B(n_124),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_514),
.B(n_0),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_492),
.B(n_146),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_514),
.B(n_146),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_505),
.B(n_146),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_598),
.B(n_467),
.Y(n_701)
);

AO32x2_ASAP7_75t_L g702 ( 
.A1(n_623),
.A2(n_523),
.A3(n_511),
.B1(n_488),
.B2(n_559),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_561),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_645),
.A2(n_630),
.B(n_578),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_595),
.B(n_471),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_572),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_566),
.B(n_471),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_610),
.A2(n_496),
.B1(n_494),
.B2(n_482),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_693),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_569),
.A2(n_510),
.B(n_512),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_534),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_586),
.A2(n_545),
.B(n_544),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_678),
.A2(n_538),
.B(n_458),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_566),
.B(n_467),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_646),
.A2(n_560),
.B(n_500),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_599),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_678),
.A2(n_453),
.B(n_491),
.Y(n_717)
);

O2A1O1Ixp5_ASAP7_75t_SL g718 ( 
.A1(n_632),
.A2(n_534),
.B(n_527),
.C(n_539),
.Y(n_718)
);

AO31x2_ASAP7_75t_L g719 ( 
.A1(n_573),
.A2(n_527),
.A3(n_482),
.B(n_499),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_570),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_583),
.A2(n_496),
.B(n_130),
.Y(n_721)
);

NAND3x1_ASAP7_75t_L g722 ( 
.A(n_677),
.B(n_1),
.C(n_2),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_577),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_617),
.A2(n_130),
.B(n_129),
.Y(n_724)
);

AOI22x1_ASAP7_75t_L g725 ( 
.A1(n_675),
.A2(n_130),
.B1(n_129),
.B2(n_132),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_590),
.B(n_146),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_591),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_693),
.Y(n_728)
);

AOI211x1_ASAP7_75t_L g729 ( 
.A1(n_594),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_729)
);

NOR2x1_ASAP7_75t_SL g730 ( 
.A(n_564),
.B(n_143),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_592),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_626),
.B(n_146),
.Y(n_732)
);

BUFx2_ASAP7_75t_R g733 ( 
.A(n_606),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_646),
.A2(n_584),
.B(n_567),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_571),
.B(n_143),
.C(n_142),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_562),
.B(n_146),
.Y(n_736)
);

OAI21x1_ASAP7_75t_SL g737 ( 
.A1(n_661),
.A2(n_8),
.B(n_9),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_596),
.B(n_143),
.C(n_142),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_660),
.B(n_146),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_660),
.B(n_610),
.Y(n_740)
);

BUFx12f_ASAP7_75t_L g741 ( 
.A(n_659),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_565),
.A2(n_563),
.B(n_573),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_647),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_570),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_585),
.A2(n_649),
.B(n_632),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_694),
.B(n_146),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_634),
.B(n_10),
.Y(n_747)
);

NAND3x1_ASAP7_75t_L g748 ( 
.A(n_694),
.B(n_12),
.C(n_14),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_599),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_146),
.Y(n_750)
);

AOI221xp5_ASAP7_75t_L g751 ( 
.A1(n_641),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.C(n_19),
.Y(n_751)
);

AO31x2_ASAP7_75t_L g752 ( 
.A1(n_687),
.A2(n_130),
.A3(n_129),
.B(n_132),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_563),
.A2(n_121),
.B(n_124),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_682),
.B(n_15),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_582),
.A2(n_121),
.B(n_124),
.Y(n_755)
);

AO22x2_ASAP7_75t_L g756 ( 
.A1(n_585),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_593),
.B(n_146),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_620),
.A2(n_130),
.A3(n_129),
.B(n_132),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_587),
.A2(n_129),
.B(n_130),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_580),
.B(n_143),
.Y(n_760)
);

OAI21x1_ASAP7_75t_L g761 ( 
.A1(n_588),
.A2(n_132),
.B(n_133),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_681),
.B(n_20),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_636),
.A2(n_132),
.B(n_133),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_611),
.B(n_23),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_683),
.B(n_24),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_622),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_SL g767 ( 
.A1(n_574),
.A2(n_133),
.B(n_127),
.C(n_125),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_593),
.B(n_132),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_568),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_697),
.B(n_24),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_576),
.A2(n_604),
.B1(n_564),
.B2(n_615),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_693),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_697),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_635),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_593),
.B(n_132),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_575),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_637),
.A2(n_132),
.B(n_133),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_674),
.B(n_29),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_652),
.B(n_29),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_693),
.Y(n_780)
);

AOI21xp33_ASAP7_75t_L g781 ( 
.A1(n_674),
.A2(n_32),
.B(n_33),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_564),
.A2(n_143),
.B1(n_142),
.B2(n_140),
.Y(n_782)
);

NOR2x1_ASAP7_75t_SL g783 ( 
.A(n_599),
.B(n_143),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_601),
.A2(n_133),
.B(n_127),
.Y(n_784)
);

NAND2x1_ASAP7_75t_L g785 ( 
.A(n_644),
.B(n_665),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_603),
.A2(n_143),
.B1(n_142),
.B2(n_140),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_582),
.A2(n_121),
.B(n_128),
.Y(n_787)
);

OAI21xp33_ASAP7_75t_L g788 ( 
.A1(n_673),
.A2(n_35),
.B(n_36),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_SL g789 ( 
.A(n_673),
.B(n_35),
.C(n_37),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_599),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_37),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_655),
.A2(n_143),
.B1(n_142),
.B2(n_140),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_631),
.B(n_38),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_613),
.B(n_38),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_651),
.A2(n_133),
.B(n_125),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_692),
.B(n_40),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_618),
.B(n_42),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_663),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_696),
.A2(n_133),
.B(n_127),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_605),
.A2(n_121),
.B(n_124),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_589),
.A2(n_133),
.B(n_125),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_667),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_644),
.Y(n_803)
);

AO31x2_ASAP7_75t_L g804 ( 
.A1(n_691),
.A2(n_43),
.A3(n_45),
.B(n_143),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_605),
.A2(n_574),
.B(n_684),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_618),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_625),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_625),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_676),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_643),
.B(n_143),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_631),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_643),
.Y(n_812)
);

BUFx12f_ASAP7_75t_L g813 ( 
.A(n_579),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_664),
.Y(n_814)
);

AOI21x1_ASAP7_75t_SL g815 ( 
.A1(n_624),
.A2(n_143),
.B(n_142),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_695),
.A2(n_143),
.B(n_142),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_684),
.A2(n_124),
.B(n_128),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_676),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_602),
.A2(n_133),
.B(n_125),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_664),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_662),
.A2(n_672),
.B(n_668),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_699),
.B(n_143),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_579),
.Y(n_823)
);

OA21x2_ASAP7_75t_L g824 ( 
.A1(n_695),
.A2(n_143),
.B(n_142),
.Y(n_824)
);

AO21x2_ASAP7_75t_L g825 ( 
.A1(n_658),
.A2(n_143),
.B(n_142),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_669),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_671),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_633),
.A2(n_140),
.B1(n_142),
.B2(n_133),
.Y(n_828)
);

NAND2x1_ASAP7_75t_L g829 ( 
.A(n_742),
.B(n_690),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_776),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_752),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_806),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_788),
.A2(n_629),
.B(n_597),
.C(n_621),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_756),
.B(n_609),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_752),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_704),
.A2(n_627),
.B(n_666),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_823),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_748),
.A2(n_614),
.B1(n_640),
.B2(n_639),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_720),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_752),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_820),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_769),
.B(n_700),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_769),
.B(n_698),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_719),
.B(n_656),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_710),
.A2(n_656),
.B(n_670),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_742),
.A2(n_680),
.B(n_688),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_717),
.A2(n_688),
.B(n_616),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_740),
.B(n_619),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_717),
.A2(n_686),
.B(n_689),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_820),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_758),
.Y(n_851)
);

OAI21x1_ASAP7_75t_SL g852 ( 
.A1(n_737),
.A2(n_607),
.B(n_685),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_749),
.B(n_690),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_710),
.A2(n_679),
.B(n_654),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_713),
.B(n_665),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_L g856 ( 
.A(n_713),
.B(n_609),
.Y(n_856)
);

OA21x2_ASAP7_75t_L g857 ( 
.A1(n_712),
.A2(n_734),
.B(n_715),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_773),
.A2(n_658),
.B(n_650),
.C(n_642),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_712),
.A2(n_721),
.B(n_753),
.Y(n_859)
);

OAI221xp5_ASAP7_75t_L g860 ( 
.A1(n_770),
.A2(n_773),
.B1(n_743),
.B2(n_751),
.C(n_781),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_752),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_766),
.Y(n_862)
);

AOI221xp5_ASAP7_75t_SL g863 ( 
.A1(n_798),
.A2(n_600),
.B1(n_628),
.B2(n_609),
.C(n_657),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_SL g864 ( 
.A(n_749),
.B(n_600),
.Y(n_864)
);

NOR2x1_ASAP7_75t_SL g865 ( 
.A(n_749),
.B(n_600),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_SL g866 ( 
.A1(n_798),
.A2(n_640),
.B(n_638),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_706),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_789),
.B(n_640),
.C(n_648),
.Y(n_868)
);

OA21x2_ASAP7_75t_L g869 ( 
.A1(n_745),
.A2(n_608),
.B(n_657),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_774),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_805),
.A2(n_821),
.B(n_707),
.Y(n_871)
);

AO21x2_ASAP7_75t_L g872 ( 
.A1(n_821),
.A2(n_608),
.B(n_657),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_802),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_753),
.A2(n_579),
.B(n_628),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_720),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_815),
.A2(n_638),
.B(n_133),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_815),
.A2(n_133),
.B(n_657),
.Y(n_877)
);

CKINVDCx11_ASAP7_75t_R g878 ( 
.A(n_741),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_805),
.B(n_579),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_789),
.A2(n_653),
.B(n_648),
.C(n_127),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_771),
.A2(n_628),
.A3(n_609),
.B(n_600),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_708),
.B(n_628),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_778),
.A2(n_653),
.B1(n_140),
.B2(n_142),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_705),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_718),
.A2(n_125),
.B(n_127),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_711),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_711),
.B(n_140),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_701),
.B(n_140),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_756),
.B(n_140),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_723),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_759),
.A2(n_125),
.B(n_127),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_762),
.B(n_140),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_727),
.Y(n_893)
);

OA21x2_ASAP7_75t_L g894 ( 
.A1(n_714),
.A2(n_140),
.B(n_142),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_749),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_758),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_731),
.A2(n_765),
.B(n_703),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_807),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_767),
.A2(n_125),
.B(n_127),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_755),
.A2(n_140),
.B(n_142),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_724),
.A2(n_125),
.B(n_127),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_755),
.A2(n_125),
.B(n_127),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_823),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_756),
.B(n_124),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_744),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_733),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_758),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_808),
.Y(n_908)
);

AOI21x1_ASAP7_75t_L g909 ( 
.A1(n_782),
.A2(n_140),
.B(n_142),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_796),
.B(n_125),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_702),
.B(n_140),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_823),
.Y(n_912)
);

BUFx12f_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_811),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_806),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_787),
.A2(n_125),
.B(n_127),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_812),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_809),
.B(n_125),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_726),
.B(n_140),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_747),
.Y(n_920)
);

OAI21x1_ASAP7_75t_L g921 ( 
.A1(n_787),
.A2(n_127),
.B(n_140),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_804),
.B(n_719),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_826),
.A2(n_140),
.B(n_142),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_814),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_761),
.A2(n_127),
.B(n_140),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_790),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_790),
.A2(n_124),
.B(n_128),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_754),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_823),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_748),
.A2(n_140),
.B(n_142),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_790),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_702),
.B(n_142),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_818),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_763),
.A2(n_142),
.B(n_124),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_702),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_777),
.A2(n_124),
.B(n_128),
.Y(n_936)
);

AO31x2_ASAP7_75t_L g937 ( 
.A1(n_702),
.A2(n_730),
.A3(n_827),
.B(n_800),
.Y(n_937)
);

BUFx8_ASAP7_75t_L g938 ( 
.A(n_809),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_732),
.A2(n_124),
.B1(n_128),
.B2(n_736),
.Y(n_939)
);

AO31x2_ASAP7_75t_L g940 ( 
.A1(n_800),
.A2(n_746),
.A3(n_791),
.B(n_794),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_862),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_884),
.B(n_729),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_839),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_859),
.A2(n_725),
.B(n_795),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_862),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_830),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_881),
.B(n_719),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_859),
.A2(n_784),
.B(n_819),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_839),
.Y(n_949)
);

OA21x2_ASAP7_75t_L g950 ( 
.A1(n_836),
.A2(n_861),
.B(n_835),
.Y(n_950)
);

OA21x2_ASAP7_75t_L g951 ( 
.A1(n_836),
.A2(n_861),
.B(n_835),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_870),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_845),
.A2(n_816),
.B(n_799),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_842),
.B(n_764),
.Y(n_954)
);

OA21x2_ASAP7_75t_L g955 ( 
.A1(n_831),
.A2(n_801),
.B(n_739),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_922),
.B(n_804),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_867),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_870),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_860),
.A2(n_793),
.B(n_722),
.C(n_750),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_833),
.A2(n_760),
.B(n_735),
.Y(n_960)
);

OA21x2_ASAP7_75t_L g961 ( 
.A1(n_831),
.A2(n_760),
.B(n_738),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_831),
.A2(n_783),
.A3(n_792),
.B(n_786),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_869),
.B(n_790),
.Y(n_963)
);

OA21x2_ASAP7_75t_L g964 ( 
.A1(n_835),
.A2(n_840),
.B(n_845),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_873),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_843),
.B(n_797),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_839),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_881),
.B(n_719),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_857),
.A2(n_822),
.B(n_757),
.Y(n_969)
);

AO21x2_ASAP7_75t_L g970 ( 
.A1(n_856),
.A2(n_855),
.B(n_840),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_838),
.A2(n_793),
.B1(n_757),
.B2(n_779),
.Y(n_971)
);

AO31x2_ASAP7_75t_L g972 ( 
.A1(n_840),
.A2(n_828),
.A3(n_804),
.B(n_817),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_866),
.A2(n_793),
.B(n_809),
.C(n_757),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_848),
.B(n_804),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_906),
.Y(n_975)
);

AOI21x1_ASAP7_75t_L g976 ( 
.A1(n_829),
.A2(n_785),
.B(n_810),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_933),
.B(n_818),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_854),
.A2(n_803),
.B(n_817),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_881),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_897),
.B(n_772),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_897),
.B(n_772),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_854),
.A2(n_803),
.B(n_780),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_873),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_881),
.B(n_758),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_829),
.A2(n_709),
.B(n_728),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_920),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_907),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_857),
.A2(n_775),
.B(n_768),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_838),
.A2(n_775),
.B1(n_768),
.B2(n_809),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_907),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_875),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_890),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_881),
.B(n_780),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_905),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_897),
.B(n_709),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_857),
.A2(n_716),
.B(n_824),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_849),
.A2(n_728),
.B(n_824),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_889),
.A2(n_775),
.B(n_768),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_893),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_889),
.A2(n_904),
.B1(n_868),
.B2(n_886),
.Y(n_1001)
);

AO22x2_ASAP7_75t_L g1002 ( 
.A1(n_922),
.A2(n_935),
.B1(n_834),
.B2(n_844),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_866),
.A2(n_716),
.B(n_813),
.C(n_824),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_893),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_841),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_898),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_898),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_879),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_879),
.Y(n_1009)
);

AO21x2_ASAP7_75t_L g1010 ( 
.A1(n_856),
.A2(n_825),
.B(n_813),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_841),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_881),
.B(n_825),
.Y(n_1012)
);

INVxp67_ASAP7_75t_SL g1013 ( 
.A(n_850),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_849),
.A2(n_124),
.B(n_128),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_904),
.A2(n_124),
.B1(n_128),
.B2(n_886),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_850),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_857),
.A2(n_128),
.B(n_858),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_928),
.B(n_128),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_908),
.Y(n_1020)
);

OA21x2_ASAP7_75t_L g1021 ( 
.A1(n_935),
.A2(n_128),
.B(n_907),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_851),
.A2(n_128),
.B(n_896),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_904),
.A2(n_128),
.B1(n_886),
.B2(n_852),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_908),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_834),
.B(n_128),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_869),
.B(n_864),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_917),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_917),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_869),
.A2(n_872),
.B(n_865),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_886),
.B(n_914),
.Y(n_1030)
);

AO21x2_ASAP7_75t_L g1031 ( 
.A1(n_855),
.A2(n_874),
.B(n_852),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_911),
.A2(n_932),
.B(n_844),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_924),
.A2(n_832),
.A3(n_915),
.B(n_865),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_924),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_879),
.Y(n_1035)
);

OA21x2_ASAP7_75t_L g1036 ( 
.A1(n_911),
.A2(n_932),
.B(n_844),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_879),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_832),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_940),
.B(n_875),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_915),
.A2(n_904),
.A3(n_851),
.B(n_896),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_871),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_863),
.A2(n_904),
.B1(n_882),
.B2(n_933),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_875),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1002),
.B(n_871),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_941),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_941),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_988),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1002),
.B(n_871),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_988),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_1041),
.A2(n_896),
.B(n_851),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_988),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_991),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_945),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_991),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_957),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_960),
.A2(n_959),
.B(n_973),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1002),
.B(n_871),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_1041),
.A2(n_851),
.B(n_896),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_945),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_952),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1008),
.B(n_844),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_952),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_991),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_958),
.Y(n_1065)
);

NAND2x1_ASAP7_75t_L g1066 ( 
.A(n_1029),
.B(n_869),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_1026),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_980),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_1025),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1008),
.B(n_926),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_997),
.A2(n_944),
.B(n_978),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_993),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_993),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1039),
.B(n_940),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_963),
.B(n_882),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1006),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_974),
.B(n_887),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1002),
.B(n_937),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_1031),
.A2(n_996),
.B(n_981),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1006),
.Y(n_1080)
);

OA21x2_ASAP7_75t_L g1081 ( 
.A1(n_979),
.A2(n_998),
.B(n_982),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_956),
.B(n_940),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1007),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_947),
.B(n_937),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_958),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_947),
.B(n_937),
.Y(n_1086)
);

BUFx4f_ASAP7_75t_SL g1087 ( 
.A(n_975),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_994),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_944),
.A2(n_847),
.B(n_923),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_965),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_965),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_1033),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1008),
.B(n_926),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1007),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1013),
.B(n_940),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_963),
.B(n_931),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_971),
.A2(n_931),
.B1(n_926),
.B2(n_895),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1020),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_983),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1026),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_983),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1020),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_985),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_985),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_963),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1000),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1004),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1004),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1024),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_968),
.B(n_937),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_968),
.B(n_937),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1024),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1027),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1026),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1038),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1033),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1027),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1033),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_978),
.A2(n_847),
.B(n_923),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_994),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1038),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_956),
.B(n_940),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1005),
.B(n_1011),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_1031),
.A2(n_874),
.B(n_872),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1028),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_979),
.B(n_937),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1028),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1034),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1034),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_984),
.B(n_1032),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_994),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1033),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1033),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1009),
.B(n_931),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_984),
.B(n_940),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_984),
.B(n_846),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_984),
.B(n_846),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1005),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1011),
.B(n_1017),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1017),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_982),
.A2(n_909),
.B(n_846),
.Y(n_1142)
);

BUFx4f_ASAP7_75t_L g1143 ( 
.A(n_961),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1033),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_994),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_964),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_964),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_964),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1032),
.B(n_846),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_964),
.Y(n_1150)
);

OA21x2_ASAP7_75t_L g1151 ( 
.A1(n_998),
.A2(n_885),
.B(n_902),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1032),
.B(n_894),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_946),
.B(n_894),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1014),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_950),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1014),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_966),
.B(n_894),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1009),
.B(n_1035),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1032),
.B(n_894),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1037),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1037),
.Y(n_1161)
);

OAI221xp5_ASAP7_75t_L g1162 ( 
.A1(n_1056),
.A2(n_971),
.B1(n_990),
.B2(n_1042),
.C(n_954),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1071),
.A2(n_986),
.B(n_1009),
.Y(n_1163)
);

OAI211xp5_ASAP7_75t_L g1164 ( 
.A1(n_1056),
.A2(n_1001),
.B(n_1042),
.C(n_990),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1077),
.A2(n_999),
.B1(n_987),
.B2(n_969),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1139),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1105),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1105),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1156),
.Y(n_1169)
);

OR2x2_ASAP7_75t_SL g1170 ( 
.A(n_1145),
.B(n_1030),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1105),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1077),
.A2(n_1003),
.B1(n_999),
.B2(n_942),
.Y(n_1172)
);

AND2x4_ASAP7_75t_SL g1173 ( 
.A(n_1075),
.B(n_949),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1139),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1155),
.A2(n_986),
.B(n_1018),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1097),
.A2(n_977),
.B1(n_1075),
.B2(n_1069),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1143),
.A2(n_989),
.B(n_872),
.Y(n_1177)
);

AOI211xp5_ASAP7_75t_L g1178 ( 
.A1(n_1097),
.A2(n_995),
.B(n_1019),
.C(n_1025),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1121),
.B(n_1035),
.Y(n_1179)
);

AOI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1068),
.A2(n_1023),
.B1(n_880),
.B2(n_949),
.C(n_967),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1070),
.B(n_1035),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1121),
.B(n_1035),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1143),
.A2(n_1031),
.B(n_892),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1075),
.A2(n_1016),
.B1(n_895),
.B2(n_931),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1121),
.B(n_1132),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1055),
.A2(n_913),
.B1(n_878),
.B2(n_910),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1055),
.A2(n_1087),
.B1(n_1069),
.B2(n_913),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1069),
.A2(n_931),
.B1(n_895),
.B2(n_992),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1068),
.A2(n_910),
.B1(n_967),
.B2(n_992),
.C(n_943),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1075),
.A2(n_1043),
.B1(n_992),
.B2(n_943),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1075),
.A2(n_1043),
.B1(n_943),
.B2(n_853),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1157),
.A2(n_1043),
.B(n_888),
.Y(n_1192)
);

OAI211xp5_ASAP7_75t_L g1193 ( 
.A1(n_1044),
.A2(n_918),
.B(n_930),
.C(n_939),
.Y(n_1193)
);

AOI322xp5_ASAP7_75t_L g1194 ( 
.A1(n_1078),
.A2(n_1012),
.A3(n_919),
.B1(n_883),
.B2(n_929),
.C1(n_912),
.C2(n_903),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1087),
.A2(n_955),
.B1(n_1012),
.B2(n_961),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1154),
.Y(n_1196)
);

AOI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1044),
.A2(n_1012),
.B1(n_903),
.B2(n_929),
.C(n_912),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1069),
.A2(n_1036),
.B1(n_938),
.B2(n_1012),
.Y(n_1198)
);

AOI221xp5_ASAP7_75t_L g1199 ( 
.A1(n_1044),
.A2(n_837),
.B1(n_929),
.B2(n_912),
.C(n_903),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1075),
.A2(n_1096),
.B1(n_1082),
.B2(n_1123),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1157),
.A2(n_955),
.B1(n_961),
.B2(n_938),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1153),
.B(n_1040),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1105),
.Y(n_1203)
);

AOI221xp5_ASAP7_75t_L g1204 ( 
.A1(n_1048),
.A2(n_837),
.B1(n_929),
.B2(n_912),
.C(n_903),
.Y(n_1204)
);

AOI322xp5_ASAP7_75t_L g1205 ( 
.A1(n_1078),
.A2(n_837),
.A3(n_929),
.B1(n_912),
.B2(n_903),
.C1(n_1036),
.C2(n_1040),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1078),
.A2(n_955),
.B1(n_961),
.B2(n_938),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1048),
.A2(n_955),
.B1(n_938),
.B2(n_1036),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1156),
.Y(n_1208)
);

AOI222xp33_ASAP7_75t_L g1209 ( 
.A1(n_1048),
.A2(n_864),
.B1(n_837),
.B2(n_1015),
.C1(n_953),
.C2(n_877),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1058),
.A2(n_1036),
.B1(n_874),
.B2(n_900),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1121),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1071),
.A2(n_950),
.B(n_951),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1143),
.B(n_837),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1075),
.A2(n_853),
.B1(n_976),
.B2(n_1021),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1160),
.B(n_1082),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1096),
.A2(n_853),
.B1(n_1021),
.B2(n_951),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_1010),
.B1(n_970),
.B2(n_948),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1160),
.Y(n_1218)
);

OAI211xp5_ASAP7_75t_L g1219 ( 
.A1(n_1058),
.A2(n_976),
.B(n_951),
.C(n_950),
.Y(n_1219)
);

OAI221xp5_ASAP7_75t_L g1220 ( 
.A1(n_1067),
.A2(n_950),
.B1(n_951),
.B2(n_1021),
.C(n_927),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1141),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1153),
.B(n_1124),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1108),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1154),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1141),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1058),
.A2(n_1123),
.B1(n_1082),
.B2(n_1143),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1095),
.A2(n_970),
.B1(n_1010),
.B2(n_900),
.C(n_1040),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1123),
.A2(n_1143),
.B1(n_1095),
.B2(n_1084),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1045),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1108),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1070),
.A2(n_1010),
.B1(n_970),
.B2(n_948),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1070),
.B(n_1040),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1084),
.A2(n_900),
.B1(n_948),
.B2(n_1021),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1154),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1084),
.A2(n_948),
.B1(n_953),
.B2(n_1015),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1045),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1046),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1086),
.A2(n_1112),
.B1(n_1111),
.B2(n_1074),
.Y(n_1238)
);

OAI211xp5_ASAP7_75t_L g1239 ( 
.A1(n_1066),
.A2(n_909),
.B(n_1022),
.C(n_877),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1066),
.A2(n_1022),
.B(n_885),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1124),
.B(n_1040),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1096),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1046),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1096),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1053),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1086),
.A2(n_876),
.B1(n_916),
.B2(n_902),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1096),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1086),
.A2(n_876),
.B1(n_916),
.B2(n_921),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1070),
.B(n_1040),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1053),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1071),
.A2(n_921),
.B(n_891),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1096),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1111),
.A2(n_899),
.B1(n_891),
.B2(n_901),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1070),
.B(n_972),
.Y(n_1254)
);

OAI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1067),
.A2(n_972),
.B1(n_962),
.B2(n_899),
.C(n_901),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1093),
.B(n_972),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1108),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1108),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1128),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1060),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1136),
.A2(n_1111),
.B1(n_1112),
.B2(n_1127),
.C(n_1074),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1096),
.A2(n_972),
.B1(n_962),
.B2(n_925),
.Y(n_1262)
);

AOI33xp33_ASAP7_75t_L g1263 ( 
.A1(n_1112),
.A2(n_972),
.A3(n_962),
.B1(n_925),
.B2(n_934),
.B3(n_936),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1106),
.B(n_972),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1074),
.A2(n_934),
.B1(n_936),
.B2(n_962),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1136),
.A2(n_962),
.B1(n_1161),
.B2(n_1154),
.Y(n_1266)
);

OR2x6_ASAP7_75t_L g1267 ( 
.A(n_1106),
.B(n_962),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1093),
.A2(n_1158),
.B1(n_1057),
.B2(n_1062),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1093),
.A2(n_1158),
.B1(n_1057),
.B2(n_1062),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1066),
.A2(n_1125),
.B(n_1135),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1161),
.B(n_1136),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1093),
.B(n_1057),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1128),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1050),
.A2(n_1059),
.B(n_1142),
.Y(n_1274)
);

OAI221xp5_ASAP7_75t_L g1275 ( 
.A1(n_1067),
.A2(n_1100),
.B1(n_1115),
.B2(n_1106),
.C(n_1135),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1135),
.A2(n_1161),
.B1(n_1106),
.B2(n_1093),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1161),
.A2(n_1093),
.B1(n_1127),
.B2(n_1125),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1140),
.B(n_1079),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1131),
.A2(n_1115),
.B(n_1100),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1060),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1057),
.B(n_1158),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1128),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1140),
.B(n_1079),
.Y(n_1283)
);

OAI211xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1145),
.A2(n_1107),
.B(n_1091),
.C(n_1090),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1061),
.Y(n_1285)
);

AOI221xp5_ASAP7_75t_L g1286 ( 
.A1(n_1127),
.A2(n_1131),
.B1(n_1115),
.B2(n_1100),
.C(n_1067),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1061),
.Y(n_1287)
);

OAI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1100),
.A2(n_1115),
.B1(n_1106),
.B2(n_1135),
.C(n_1132),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_L g1289 ( 
.A(n_1092),
.B(n_1117),
.C(n_1144),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1135),
.A2(n_1062),
.B1(n_1158),
.B2(n_1057),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1202),
.B(n_1079),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1222),
.B(n_1079),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1166),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1174),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1162),
.A2(n_1062),
.B1(n_1158),
.B2(n_1057),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1221),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1167),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1167),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1244),
.B(n_1132),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1225),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1165),
.B(n_1079),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1168),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1244),
.B(n_1132),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1165),
.B(n_1063),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1229),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1185),
.B(n_1088),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1168),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1185),
.B(n_1088),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1236),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1237),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1172),
.B(n_1158),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1267),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1245),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1215),
.B(n_1122),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1250),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1185),
.B(n_1088),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1272),
.B(n_1088),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1244),
.B(n_1088),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1260),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1280),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1281),
.B(n_1131),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1228),
.B(n_1109),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1228),
.B(n_1109),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1171),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1171),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1241),
.B(n_1122),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1285),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1169),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1238),
.B(n_1122),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1259),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1273),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1282),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1181),
.B(n_1268),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1287),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1176),
.A2(n_1062),
.B1(n_1135),
.B2(n_1138),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1269),
.B(n_1062),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1238),
.B(n_1116),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1226),
.A2(n_1135),
.B1(n_1138),
.B2(n_1137),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1211),
.B(n_1179),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1211),
.B(n_1137),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1203),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1179),
.B(n_1137),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1242),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1208),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1226),
.A2(n_1138),
.B1(n_1152),
.B2(n_1125),
.Y(n_1347)
);

INVx5_ASAP7_75t_L g1348 ( 
.A(n_1267),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1179),
.B(n_1116),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1223),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1182),
.B(n_1116),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1223),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1230),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1164),
.A2(n_1152),
.B1(n_1125),
.B2(n_1149),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1230),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1182),
.B(n_1116),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1242),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1182),
.B(n_1232),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1249),
.B(n_1242),
.Y(n_1359)
);

NAND4xp25_ASAP7_75t_L g1360 ( 
.A(n_1178),
.B(n_1149),
.C(n_1134),
.D(n_1159),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1213),
.B(n_1242),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1247),
.B(n_1122),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1257),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1257),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1192),
.B(n_1104),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1258),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1247),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1261),
.B(n_1104),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1218),
.B(n_1103),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1258),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1247),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1278),
.B(n_1128),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1247),
.B(n_1073),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1252),
.B(n_1119),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1284),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1271),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1194),
.B(n_1283),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1170),
.B(n_1129),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1254),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1183),
.B(n_1103),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1196),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1234),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1252),
.B(n_1102),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1252),
.B(n_1102),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1289),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1277),
.B(n_1129),
.Y(n_1386)
);

NOR2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1252),
.B(n_1149),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1189),
.B(n_1099),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1177),
.B(n_1099),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1256),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1277),
.B(n_1129),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1173),
.B(n_1133),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1286),
.B(n_1101),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1358),
.B(n_1279),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1330),
.B(n_1290),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1293),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1293),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1375),
.B(n_1205),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1304),
.B(n_1187),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1378),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1354),
.B(n_1187),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1358),
.B(n_1173),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1359),
.B(n_1224),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1359),
.B(n_1276),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1347),
.A2(n_1186),
.B1(n_1200),
.B2(n_1266),
.C(n_1207),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1340),
.B(n_1213),
.Y(n_1406)
);

AND2x4_ASAP7_75t_SL g1407 ( 
.A(n_1381),
.B(n_1267),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_SL g1408 ( 
.A(n_1378),
.B(n_1190),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_SL g1409 ( 
.A(n_1360),
.B(n_1275),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1330),
.B(n_1129),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1340),
.B(n_1188),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1375),
.B(n_1180),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1294),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1295),
.B(n_1191),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1296),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1338),
.B(n_1264),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1338),
.B(n_1264),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1388),
.B(n_1186),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1349),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1385),
.B(n_1288),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1377),
.B(n_1266),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1296),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1300),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1300),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1305),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1393),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1305),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1313),
.B(n_1119),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1309),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1346),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1385),
.B(n_1197),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1309),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1310),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1310),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1368),
.B(n_1199),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1312),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1323),
.B(n_1072),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1324),
.B(n_1072),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1312),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1345),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1349),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1345),
.B(n_1198),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1351),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1351),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1380),
.B(n_1072),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_SL g1448 ( 
.A(n_1357),
.B(n_1184),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1335),
.B(n_1204),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1356),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1357),
.B(n_1207),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1316),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1311),
.B(n_1193),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1389),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1335),
.B(n_1201),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1313),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1316),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1313),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1371),
.B(n_1195),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1301),
.B(n_1201),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1365),
.B(n_1195),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1329),
.B(n_1063),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1356),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1297),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1376),
.B(n_1065),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1320),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1371),
.B(n_1206),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_SL g1469 ( 
.A(n_1313),
.B(n_1348),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1297),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1320),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1321),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1299),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1334),
.B(n_1206),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1334),
.B(n_1217),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1361),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1376),
.B(n_1065),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1367),
.B(n_1231),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1321),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1382),
.B(n_1085),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1313),
.B(n_1270),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1328),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1313),
.B(n_1119),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1367),
.B(n_1175),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1298),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_L g1486 ( 
.A(n_1348),
.B(n_1219),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1367),
.B(n_1175),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1299),
.B(n_1175),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1400),
.B(n_1386),
.Y(n_1489)
);

NOR3xp33_ASAP7_75t_L g1490 ( 
.A(n_1401),
.B(n_1292),
.C(n_1382),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1422),
.A2(n_1339),
.B1(n_1336),
.B2(n_1386),
.Y(n_1491)
);

NOR3xp33_ASAP7_75t_L g1492 ( 
.A(n_1405),
.B(n_1291),
.C(n_1391),
.Y(n_1492)
);

NAND4xp25_ASAP7_75t_L g1493 ( 
.A(n_1412),
.B(n_1391),
.C(n_1291),
.D(n_1227),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1397),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1457),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1441),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1469),
.A2(n_1319),
.B(n_1331),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1399),
.A2(n_1387),
.B1(n_1303),
.B2(n_1299),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1400),
.B(n_1327),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1409),
.A2(n_1448),
.B1(n_1398),
.B2(n_1436),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1441),
.Y(n_1501)
);

OAI31xp33_ASAP7_75t_L g1502 ( 
.A1(n_1419),
.A2(n_1387),
.A3(n_1361),
.B(n_1216),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_SL g1503 ( 
.A(n_1427),
.B(n_1361),
.C(n_1337),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1484),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1394),
.B(n_1299),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1394),
.B(n_1303),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1457),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1454),
.A2(n_1303),
.B1(n_1348),
.B2(n_1337),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1431),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1455),
.B(n_1362),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1457),
.B(n_1303),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1461),
.B(n_1348),
.C(n_1333),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1473),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1432),
.A2(n_1319),
.B(n_1348),
.Y(n_1514)
);

OA332x1_ASAP7_75t_L g1515 ( 
.A1(n_1408),
.A2(n_1214),
.A3(n_1262),
.B1(n_1348),
.B2(n_1327),
.B3(n_1372),
.C1(n_1379),
.C2(n_1390),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1408),
.B(n_1306),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1411),
.B(n_1402),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1374),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1487),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1487),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1411),
.B(n_1306),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1443),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1410),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1462),
.A2(n_1390),
.B1(n_1379),
.B2(n_1369),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1402),
.B(n_1308),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1438),
.B(n_1372),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1406),
.B(n_1308),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1406),
.B(n_1317),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1414),
.A2(n_1374),
.B1(n_1317),
.B2(n_1344),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1486),
.A2(n_1333),
.B(n_1331),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1397),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1438),
.B(n_1332),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1413),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1413),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1404),
.B(n_1344),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1439),
.B(n_1332),
.Y(n_1537)
);

OAI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1421),
.A2(n_1328),
.B1(n_1362),
.B2(n_1384),
.C(n_1373),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1423),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1396),
.B(n_1298),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1423),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1424),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1404),
.B(n_1443),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_SL g1544 ( 
.A1(n_1478),
.A2(n_1383),
.B(n_1373),
.C(n_1384),
.Y(n_1544)
);

AOI33xp33_ASAP7_75t_L g1545 ( 
.A1(n_1475),
.A2(n_1383),
.A3(n_1210),
.B1(n_1355),
.B2(n_1341),
.B3(n_1353),
.Y(n_1545)
);

AOI33xp33_ASAP7_75t_L g1546 ( 
.A1(n_1475),
.A2(n_1210),
.A3(n_1341),
.B1(n_1363),
.B2(n_1353),
.B3(n_1355),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1424),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1459),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1456),
.A2(n_1352),
.B1(n_1350),
.B2(n_1363),
.C(n_1374),
.Y(n_1549)
);

OAI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1421),
.A2(n_1350),
.B1(n_1352),
.B2(n_1370),
.C(n_1302),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1473),
.B(n_1322),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1410),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1459),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1459),
.B(n_1374),
.Y(n_1554)
);

AOI222xp33_ASAP7_75t_L g1555 ( 
.A1(n_1449),
.A2(n_1152),
.B1(n_1220),
.B2(n_1117),
.C1(n_1144),
.C2(n_1092),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1407),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1468),
.B(n_1322),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1420),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1476),
.B(n_1392),
.Y(n_1559)
);

OAI33xp33_ASAP7_75t_L g1560 ( 
.A1(n_1425),
.A2(n_1315),
.A3(n_1325),
.B1(n_1370),
.B2(n_1343),
.B3(n_1302),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1474),
.A2(n_1392),
.B1(n_1342),
.B2(n_1209),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1415),
.B(n_1307),
.Y(n_1562)
);

NOR3xp33_ASAP7_75t_L g1563 ( 
.A(n_1476),
.B(n_1163),
.C(n_1239),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1543),
.B(n_1468),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1535),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1496),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1523),
.B(n_1474),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1501),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1425),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1543),
.B(n_1452),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1501),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1523),
.B(n_1439),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1509),
.B(n_1460),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1501),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1517),
.B(n_1460),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1517),
.B(n_1452),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1557),
.B(n_1403),
.Y(n_1577)
);

NAND2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_SL g1579 ( 
.A(n_1502),
.B(n_1511),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1494),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1511),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1557),
.B(n_1403),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1478),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1495),
.B(n_1417),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1513),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1507),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1513),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1556),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1511),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1536),
.B(n_1420),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1522),
.B(n_1442),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1514),
.A2(n_1485),
.B(n_1465),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1494),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1532),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1553),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1553),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1522),
.B(n_1442),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1489),
.B(n_1447),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1500),
.B(n_1444),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1512),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1489),
.B(n_1447),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1505),
.B(n_1444),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1532),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1490),
.B(n_1446),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1534),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1505),
.B(n_1450),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1558),
.B(n_1426),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1506),
.B(n_1450),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1506),
.B(n_1464),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1558),
.B(n_1426),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1530),
.B(n_1464),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1512),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1548),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1526),
.B(n_1407),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1495),
.B(n_1463),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1526),
.B(n_1395),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1558),
.B(n_1428),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1519),
.B(n_1428),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1528),
.B(n_1395),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1533),
.B(n_1430),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1534),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1519),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1533),
.B(n_1430),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1548),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1539),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1528),
.B(n_1529),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1546),
.B(n_1416),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1539),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1529),
.B(n_1516),
.Y(n_1630)
);

INVx5_ASAP7_75t_L g1631 ( 
.A(n_1495),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1600),
.B(n_1495),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1566),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1564),
.B(n_1544),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1568),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1576),
.B(n_1556),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1564),
.B(n_1545),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1568),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1567),
.B(n_1510),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1570),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1575),
.B(n_1493),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1596),
.B(n_1548),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1630),
.B(n_1516),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1596),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1579),
.A2(n_1491),
.B1(n_1493),
.B2(n_1502),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1596),
.B(n_1548),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1491),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1614),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1568),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1605),
.B(n_1499),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1554),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1614),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_SL g1657 ( 
.A(n_1615),
.B(n_1519),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1571),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1571),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1574),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1604),
.B(n_1499),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1503),
.Y(n_1663)
);

NAND2x1_ASAP7_75t_L g1664 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1589),
.B(n_1549),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1574),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1612),
.B(n_1572),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1572),
.B(n_1498),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1586),
.B(n_1560),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1595),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1599),
.B(n_1561),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1595),
.Y(n_1673)
);

OR2x6_ASAP7_75t_L g1674 ( 
.A(n_1581),
.B(n_1514),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1581),
.B(n_1595),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1580),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1551),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1580),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1627),
.B(n_1551),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1593),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1582),
.B(n_1554),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1625),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1628),
.B(n_1525),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1582),
.B(n_1559),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1593),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1620),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1623),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1594),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1594),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1583),
.B(n_1559),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1592),
.A2(n_1563),
.B(n_1508),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1631),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1620),
.B(n_1537),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1603),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1617),
.B(n_1537),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1617),
.B(n_1417),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1583),
.B(n_1559),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1633),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1670),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1648),
.A2(n_1615),
.B1(n_1602),
.B2(n_1607),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1645),
.B(n_1585),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1647),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1694),
.B(n_1584),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1648),
.A2(n_1602),
.B1(n_1607),
.B2(n_1610),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1650),
.A2(n_1687),
.B1(n_1672),
.B2(n_1684),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1647),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1683),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1683),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1671),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1673),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1657),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1684),
.A2(n_1610),
.B1(n_1597),
.B2(n_1591),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1635),
.B(n_1565),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1669),
.B(n_1565),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1670),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1670),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1696),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1677),
.B(n_1680),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1639),
.A2(n_1623),
.B1(n_1418),
.B2(n_1578),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1669),
.B(n_1585),
.Y(n_1723)
);

AOI32xp33_ASAP7_75t_L g1724 ( 
.A1(n_1665),
.A2(n_1597),
.A3(n_1616),
.B1(n_1592),
.B2(n_1590),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1675),
.B(n_1688),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1664),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1675),
.B(n_1585),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1687),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1637),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1634),
.B(n_1590),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1640),
.Y(n_1731)
);

NAND2x1_ASAP7_75t_L g1732 ( 
.A(n_1649),
.B(n_1584),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1638),
.A2(n_1531),
.B1(n_1555),
.B2(n_1584),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1653),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1649),
.B(n_1587),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1644),
.A2(n_1418),
.B1(n_1578),
.B2(n_1515),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1658),
.Y(n_1738)
);

NAND2xp33_ASAP7_75t_SL g1739 ( 
.A(n_1638),
.B(n_1587),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1659),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1660),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1632),
.A2(n_1606),
.B1(n_1629),
.B2(n_1626),
.C(n_1603),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1667),
.A2(n_1578),
.B1(n_1587),
.B2(n_1631),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1652),
.B(n_1606),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1649),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1666),
.Y(n_1746)
);

OAI22xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1674),
.A2(n_1631),
.B1(n_1569),
.B2(n_1619),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1652),
.Y(n_1748)
);

INVx4_ASAP7_75t_L g1749 ( 
.A(n_1700),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1703),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1728),
.B(n_1641),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1655),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1708),
.B(n_1716),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1709),
.Y(n_1754)
);

AOI32xp33_ASAP7_75t_L g1755 ( 
.A1(n_1737),
.A2(n_1655),
.A3(n_1682),
.B1(n_1679),
.B2(n_1662),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1736),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1710),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1736),
.B(n_1656),
.Y(n_1758)
);

NAND2xp67_ASAP7_75t_L g1759 ( 
.A(n_1745),
.B(n_1656),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1702),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1732),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1733),
.A2(n_1654),
.B1(n_1651),
.B2(n_1636),
.Y(n_1762)
);

AOI222xp33_ASAP7_75t_L g1763 ( 
.A1(n_1716),
.A2(n_1692),
.B1(n_1632),
.B2(n_1695),
.C1(n_1678),
.C2(n_1676),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1723),
.B(n_1661),
.Y(n_1764)
);

NOR2x1_ASAP7_75t_L g1765 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1735),
.Y(n_1766)
);

AOI32xp33_ASAP7_75t_L g1767 ( 
.A1(n_1722),
.A2(n_1662),
.A3(n_1679),
.B1(n_1682),
.B2(n_1691),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1707),
.A2(n_1674),
.B(n_1668),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1723),
.A2(n_1631),
.B(n_1663),
.C(n_1693),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1730),
.Y(n_1771)
);

AND2x4_ASAP7_75t_SL g1772 ( 
.A(n_1726),
.B(n_1691),
.Y(n_1772)
);

OAI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1724),
.A2(n_1693),
.B1(n_1690),
.B2(n_1689),
.C(n_1686),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1748),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1707),
.A2(n_1681),
.B(n_1642),
.C(n_1531),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1704),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1705),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1720),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1744),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1747),
.A2(n_1698),
.B(n_1685),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_L g1781 ( 
.A(n_1701),
.B(n_1698),
.C(n_1685),
.D(n_1697),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1713),
.A2(n_1646),
.B1(n_1531),
.B2(n_1555),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1706),
.A2(n_1646),
.B(n_1598),
.Y(n_1783)
);

XOR2x2_ASAP7_75t_L g1784 ( 
.A(n_1714),
.B(n_1721),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1699),
.B(n_1622),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1727),
.B(n_1622),
.Y(n_1786)
);

OAI211xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1742),
.A2(n_1626),
.B(n_1629),
.C(n_1601),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1744),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1715),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1715),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1763),
.B(n_1727),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1763),
.A2(n_1739),
.B1(n_1725),
.B2(n_1743),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1756),
.B(n_1725),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1758),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1759),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1751),
.B(n_1711),
.Y(n_1796)
);

AOI311xp33_ASAP7_75t_L g1797 ( 
.A1(n_1762),
.A2(n_1742),
.A3(n_1743),
.B(n_1712),
.C(n_1741),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1752),
.B(n_1729),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1758),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1772),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1771),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1775),
.A2(n_1631),
.B(n_1734),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1768),
.A2(n_1631),
.B(n_1740),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1749),
.Y(n_1805)
);

OAI32xp33_ASAP7_75t_L g1806 ( 
.A1(n_1782),
.A2(n_1746),
.A3(n_1738),
.B1(n_1624),
.B2(n_1621),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1764),
.B(n_1598),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1765),
.Y(n_1808)
);

OAI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1764),
.A2(n_1601),
.B1(n_1624),
.B2(n_1621),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1760),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1773),
.A2(n_1550),
.B1(n_1618),
.B2(n_1611),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1750),
.Y(n_1813)
);

NAND2x1p5_ASAP7_75t_L g1814 ( 
.A(n_1761),
.B(n_1569),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1768),
.B(n_1619),
.C(n_1569),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_SL g1816 ( 
.A(n_1773),
.B(n_1753),
.C(n_1767),
.Y(n_1816)
);

AOI32xp33_ASAP7_75t_L g1817 ( 
.A1(n_1762),
.A2(n_1619),
.A3(n_1569),
.B1(n_1542),
.B2(n_1547),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1755),
.B(n_1619),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1785),
.Y(n_1819)
);

XNOR2x2_ASAP7_75t_L g1820 ( 
.A(n_1753),
.B(n_1608),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1776),
.A2(n_1497),
.B1(n_1542),
.B2(n_1541),
.Y(n_1821)
);

OAI32xp33_ASAP7_75t_L g1822 ( 
.A1(n_1783),
.A2(n_1787),
.A3(n_1789),
.B1(n_1790),
.B2(n_1786),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1785),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1777),
.B(n_1497),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1778),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1754),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1770),
.A2(n_1547),
.B1(n_1541),
.B2(n_1552),
.C(n_1524),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1781),
.A2(n_1618),
.B1(n_1611),
.B2(n_1608),
.C(n_1524),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1757),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1797),
.B(n_1780),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1816),
.A2(n_1788),
.B1(n_1779),
.B2(n_1786),
.C(n_1766),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1794),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1820),
.Y(n_1833)
);

NAND2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1791),
.B(n_1774),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_L g1835 ( 
.A1(n_1791),
.A2(n_1784),
.B(n_1524),
.C(n_1552),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1799),
.B(n_1552),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_L g1837 ( 
.A(n_1792),
.B(n_1520),
.C(n_1518),
.Y(n_1837)
);

OAI211xp5_ASAP7_75t_L g1838 ( 
.A1(n_1822),
.A2(n_1518),
.B(n_1504),
.C(n_1520),
.Y(n_1838)
);

NAND4xp25_ASAP7_75t_L g1839 ( 
.A(n_1818),
.B(n_1520),
.C(n_1504),
.D(n_1518),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1800),
.B(n_1440),
.Y(n_1840)
);

AOI322xp5_ASAP7_75t_L g1841 ( 
.A1(n_1812),
.A2(n_1521),
.A3(n_1504),
.B1(n_1488),
.B2(n_1562),
.C1(n_1540),
.C2(n_1483),
.Y(n_1841)
);

OAI21xp33_ASAP7_75t_L g1842 ( 
.A1(n_1796),
.A2(n_1521),
.B(n_1562),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1806),
.A2(n_1497),
.B(n_1540),
.Y(n_1843)
);

OAI211xp5_ASAP7_75t_SL g1844 ( 
.A1(n_1817),
.A2(n_1521),
.B(n_1527),
.C(n_1445),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1803),
.A2(n_1804),
.B(n_1809),
.Y(n_1845)
);

NOR3xp33_ASAP7_75t_L g1846 ( 
.A(n_1793),
.B(n_1527),
.C(n_1453),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1808),
.A2(n_1433),
.B1(n_1458),
.B2(n_1482),
.C(n_1434),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1793),
.A2(n_1437),
.B(n_1458),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1814),
.B(n_1318),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1814),
.Y(n_1850)
);

AOI221x1_ASAP7_75t_L g1851 ( 
.A1(n_1795),
.A2(n_1434),
.B1(n_1453),
.B2(n_1451),
.C(n_1482),
.Y(n_1851)
);

OAI321xp33_ASAP7_75t_L g1852 ( 
.A1(n_1815),
.A2(n_1488),
.A3(n_1433),
.B1(n_1437),
.B2(n_1479),
.C(n_1435),
.Y(n_1852)
);

NOR3x1_ASAP7_75t_L g1853 ( 
.A(n_1798),
.B(n_1451),
.C(n_1435),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1811),
.A2(n_1479),
.B(n_1467),
.C(n_1472),
.Y(n_1854)
);

NAND4xp25_ASAP7_75t_L g1855 ( 
.A(n_1807),
.B(n_1801),
.C(n_1805),
.D(n_1825),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1828),
.A2(n_1483),
.B(n_1429),
.Y(n_1856)
);

OAI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1811),
.A2(n_1471),
.B(n_1485),
.C(n_1470),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1802),
.A2(n_1470),
.B(n_1465),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1802),
.A2(n_1480),
.B(n_1477),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1824),
.A2(n_1466),
.B(n_1483),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1819),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1833),
.A2(n_1823),
.B(n_1827),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1830),
.A2(n_1826),
.B1(n_1813),
.B2(n_1829),
.C(n_1810),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1832),
.Y(n_1864)
);

AOI322xp5_ASAP7_75t_L g1865 ( 
.A1(n_1834),
.A2(n_1831),
.A3(n_1850),
.B1(n_1861),
.B2(n_1842),
.C1(n_1846),
.C2(n_1840),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1849),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.B(n_1821),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1856),
.A2(n_1326),
.B1(n_1366),
.B2(n_1364),
.C(n_1343),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1839),
.A2(n_1429),
.B(n_1392),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1855),
.B(n_1315),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1845),
.A2(n_1429),
.B(n_1307),
.Y(n_1871)
);

AOI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1852),
.A2(n_1342),
.B1(n_1366),
.B2(n_1364),
.C(n_1325),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1837),
.A2(n_1392),
.B1(n_1318),
.B2(n_1326),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1843),
.A2(n_1274),
.B(n_1212),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1836),
.Y(n_1875)
);

AOI32xp33_ASAP7_75t_L g1876 ( 
.A1(n_1844),
.A2(n_1274),
.A3(n_1133),
.B1(n_1134),
.B2(n_1155),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1853),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1838),
.A2(n_1133),
.B1(n_1134),
.B2(n_1235),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1847),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1847),
.Y(n_1880)
);

OAI31xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1854),
.A2(n_1155),
.A3(n_1150),
.B(n_1148),
.Y(n_1881)
);

AOI32xp33_ASAP7_75t_L g1882 ( 
.A1(n_1841),
.A2(n_1134),
.A3(n_1155),
.B1(n_1130),
.B2(n_1118),
.Y(n_1882)
);

AOI21xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1857),
.A2(n_1081),
.B(n_1125),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1859),
.A2(n_1848),
.B1(n_1858),
.B2(n_1860),
.C(n_1851),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1866),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1864),
.Y(n_1886)
);

XNOR2x1_ASAP7_75t_L g1887 ( 
.A(n_1867),
.B(n_1081),
.Y(n_1887)
);

A2O1A1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1862),
.A2(n_1865),
.B(n_1871),
.C(n_1884),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1870),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1877),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1869),
.A2(n_1081),
.B1(n_1114),
.B2(n_1085),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1879),
.Y(n_1892)
);

AOI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1863),
.A2(n_1255),
.B(n_1130),
.C(n_1126),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1880),
.Y(n_1894)
);

OAI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1873),
.A2(n_1146),
.B1(n_1147),
.B2(n_1150),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1875),
.A2(n_1235),
.B(n_1265),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1874),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1868),
.Y(n_1898)
);

OAI222xp33_ASAP7_75t_L g1899 ( 
.A1(n_1876),
.A2(n_1159),
.B1(n_1126),
.B2(n_1107),
.C1(n_1090),
.C2(n_1091),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1883),
.A2(n_1150),
.B1(n_1148),
.B2(n_1147),
.C(n_1146),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1878),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1881),
.A2(n_1150),
.B(n_1148),
.C(n_1147),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1888),
.A2(n_1872),
.B(n_1881),
.C(n_1882),
.Y(n_1903)
);

A2O1A1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1885),
.A2(n_1263),
.B(n_1118),
.C(n_1114),
.Y(n_1904)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1905 ( 
.A1(n_1890),
.A2(n_1101),
.B(n_1110),
.C(n_1113),
.D(n_1263),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1889),
.A2(n_1113),
.B(n_1110),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1901),
.A2(n_1081),
.B1(n_1146),
.B2(n_1148),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1892),
.A2(n_1265),
.B(n_1233),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1146),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1898),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1886),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1891),
.A2(n_1147),
.B1(n_1233),
.B2(n_1081),
.Y(n_1912)
);

AOI32xp33_ASAP7_75t_L g1913 ( 
.A1(n_1887),
.A2(n_1893),
.A3(n_1895),
.B1(n_1900),
.B2(n_1897),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_SL g1914 ( 
.A1(n_1896),
.A2(n_1083),
.B1(n_1072),
.B2(n_1102),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1899),
.A2(n_1098),
.B1(n_1094),
.B2(n_1102),
.C(n_1080),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1900),
.A2(n_1081),
.B1(n_1098),
.B2(n_1094),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1902),
.A2(n_1073),
.B(n_1080),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1902),
.A2(n_1159),
.B1(n_1073),
.B2(n_1098),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1886),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1911),
.B(n_1083),
.Y(n_1920)
);

INVxp33_ASAP7_75t_SL g1921 ( 
.A(n_1919),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1910),
.B(n_1083),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1910),
.B(n_1083),
.Y(n_1923)
);

NOR2x1_ASAP7_75t_SL g1924 ( 
.A(n_1908),
.B(n_1094),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1903),
.B(n_1098),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1909),
.Y(n_1926)
);

NOR2x1_ASAP7_75t_L g1927 ( 
.A(n_1906),
.B(n_1080),
.Y(n_1927)
);

OAI211xp5_ASAP7_75t_L g1928 ( 
.A1(n_1913),
.A2(n_1080),
.B(n_1076),
.C(n_1094),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1914),
.Y(n_1929)
);

NOR2x1_ASAP7_75t_L g1930 ( 
.A(n_1918),
.B(n_1076),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1907),
.A2(n_1076),
.B(n_1073),
.C(n_1051),
.Y(n_1931)
);

NOR2xp67_ASAP7_75t_L g1932 ( 
.A(n_1912),
.B(n_1076),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1926),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1924),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1921),
.A2(n_1916),
.B1(n_1917),
.B2(n_1904),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1925),
.A2(n_1915),
.B1(n_1905),
.B2(n_1047),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1922),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1929),
.Y(n_1938)
);

OAI211xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1938),
.A2(n_1920),
.B(n_1923),
.C(n_1928),
.Y(n_1939)
);

AOI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1933),
.A2(n_1931),
.B1(n_1932),
.B2(n_1927),
.C(n_1930),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1934),
.Y(n_1941)
);

OAI211xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1935),
.A2(n_1253),
.B(n_1248),
.C(n_1246),
.Y(n_1942)
);

NOR3xp33_ASAP7_75t_L g1943 ( 
.A(n_1937),
.B(n_1240),
.C(n_1089),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1936),
.A2(n_1049),
.B1(n_1051),
.B2(n_1052),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1938),
.B(n_1049),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1941),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1945),
.B(n_1052),
.Y(n_1947)
);

NOR3xp33_ASAP7_75t_SL g1948 ( 
.A(n_1939),
.B(n_1089),
.C(n_1120),
.Y(n_1948)
);

NOR3xp33_ASAP7_75t_L g1949 ( 
.A(n_1940),
.B(n_1089),
.C(n_1120),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1943),
.Y(n_1950)
);

XNOR2xp5_ASAP7_75t_L g1951 ( 
.A(n_1944),
.B(n_1120),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1946),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1950),
.B(n_1947),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1948),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1949),
.B(n_1942),
.Y(n_1955)
);

XNOR2xp5_ASAP7_75t_L g1956 ( 
.A(n_1951),
.B(n_1142),
.Y(n_1956)
);

XNOR2xp5_ASAP7_75t_L g1957 ( 
.A(n_1952),
.B(n_1142),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1954),
.Y(n_1958)
);

AND3x4_ASAP7_75t_L g1959 ( 
.A(n_1955),
.B(n_1052),
.C(n_1049),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1953),
.A2(n_1956),
.B(n_1251),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1952),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1961),
.A2(n_1049),
.B(n_1054),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1958),
.B(n_1960),
.Y(n_1963)
);

AO22x2_ASAP7_75t_L g1964 ( 
.A1(n_1959),
.A2(n_1051),
.B1(n_1052),
.B2(n_1054),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1963),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1965),
.A2(n_1957),
.B1(n_1962),
.B2(n_1964),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1966),
.A2(n_1047),
.B1(n_1064),
.B2(n_1051),
.Y(n_1967)
);

AOI222xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1967),
.A2(n_1047),
.B1(n_1064),
.B2(n_1054),
.C1(n_1059),
.C2(n_1050),
.Y(n_1968)
);

AOI222xp33_ASAP7_75t_L g1969 ( 
.A1(n_1968),
.A2(n_1054),
.B1(n_1064),
.B2(n_1047),
.C1(n_1059),
.C2(n_1050),
.Y(n_1969)
);

AO21x2_ASAP7_75t_L g1970 ( 
.A1(n_1969),
.A2(n_1047),
.B(n_1064),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_SL g1971 ( 
.A1(n_1970),
.A2(n_1064),
.B1(n_1151),
.B2(n_1253),
.Y(n_1971)
);

AOI211xp5_ASAP7_75t_L g1972 ( 
.A1(n_1971),
.A2(n_1151),
.B(n_1248),
.C(n_1246),
.Y(n_1972)
);


endmodule