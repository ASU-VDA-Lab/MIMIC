module real_aes_6263_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g251 ( .A1(n_0), .A2(n_252), .B(n_253), .C(n_256), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_1), .B(n_193), .Y(n_257) );
INVx1_ASAP7_75t_L g432 ( .A(n_2), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_3), .B(n_163), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_4), .A2(n_133), .B(n_136), .C(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_153), .B(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_6), .A2(n_153), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_7), .B(n_193), .Y(n_520) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_8), .A2(n_120), .B(n_173), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_9), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_9), .Y(n_741) );
AND2x6_ASAP7_75t_L g133 ( .A(n_10), .B(n_134), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_11), .A2(n_133), .B(n_136), .C(n_139), .Y(n_135) );
INVx1_ASAP7_75t_L g490 ( .A(n_12), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_13), .B(n_41), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_14), .A2(n_45), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_14), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_15), .B(n_143), .Y(n_476) );
INVx1_ASAP7_75t_L g125 ( .A(n_16), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_17), .B(n_163), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_18), .A2(n_141), .B(n_498), .C(n_500), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_19), .B(n_193), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_20), .B(n_217), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_21), .A2(n_136), .B(n_180), .C(n_213), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_22), .A2(n_145), .B(n_255), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_23), .B(n_143), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_24), .B(n_143), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_25), .Y(n_548) );
INVx1_ASAP7_75t_L g540 ( .A(n_26), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_27), .A2(n_136), .B(n_176), .C(n_180), .Y(n_175) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_28), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_29), .Y(n_472) );
INVx1_ASAP7_75t_L g531 ( .A(n_30), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_31), .A2(n_153), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g131 ( .A(n_32), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_33), .A2(n_155), .B(n_166), .C(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_34), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_35), .A2(n_255), .B(n_517), .C(n_519), .Y(n_516) );
INVxp67_ASAP7_75t_L g532 ( .A(n_36), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_37), .A2(n_78), .B1(n_435), .B2(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_37), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_38), .B(n_178), .Y(n_177) );
CKINVDCx14_ASAP7_75t_R g515 ( .A(n_39), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_40), .A2(n_136), .B(n_180), .C(n_539), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_42), .A2(n_256), .B(n_488), .C(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_43), .B(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_44), .Y(n_148) );
INVx1_ASAP7_75t_L g739 ( .A(n_45), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_46), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_47), .B(n_153), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_48), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_49), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_50), .A2(n_155), .B(n_157), .C(n_166), .Y(n_154) );
INVx1_ASAP7_75t_L g254 ( .A(n_51), .Y(n_254) );
INVx1_ASAP7_75t_L g158 ( .A(n_52), .Y(n_158) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_53), .A2(n_458), .B1(n_732), .B2(n_733), .C1(n_742), .C2(n_745), .Y(n_457) );
INVx1_ASAP7_75t_L g505 ( .A(n_54), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_55), .B(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_56), .A2(n_59), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_56), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_57), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g486 ( .A(n_58), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_59), .Y(n_108) );
INVx1_ASAP7_75t_L g134 ( .A(n_60), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_61), .B(n_153), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_62), .B(n_193), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_63), .A2(n_187), .B(n_189), .C(n_191), .Y(n_186) );
INVx1_ASAP7_75t_L g124 ( .A(n_64), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_65), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g518 ( .A(n_66), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_67), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_68), .B(n_163), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_69), .B(n_193), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_70), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g551 ( .A(n_71), .Y(n_551) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_72), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_73), .B(n_160), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_74), .A2(n_136), .B(n_166), .C(n_227), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_75), .Y(n_185) );
INVx1_ASAP7_75t_L g452 ( .A(n_76), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_77), .A2(n_153), .B(n_485), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_78), .A2(n_104), .B1(n_444), .B2(n_453), .C1(n_456), .C2(n_748), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_78), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_79), .A2(n_153), .B(n_495), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_80), .A2(n_211), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g496 ( .A(n_81), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_82), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_83), .B(n_159), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_84), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_85), .A2(n_153), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g499 ( .A(n_86), .Y(n_499) );
INVx2_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx1_ASAP7_75t_L g475 ( .A(n_88), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_89), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_90), .B(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g429 ( .A(n_91), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g461 ( .A(n_91), .B(n_431), .Y(n_461) );
INVx2_ASAP7_75t_L g731 ( .A(n_91), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_92), .A2(n_136), .B(n_166), .C(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_93), .B(n_153), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_94), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_94), .Y(n_734) );
INVx1_ASAP7_75t_L g202 ( .A(n_95), .Y(n_202) );
INVxp67_ASAP7_75t_L g190 ( .A(n_96), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_97), .B(n_120), .Y(n_491) );
INVx1_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
INVx1_ASAP7_75t_L g228 ( .A(n_99), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_100), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g508 ( .A(n_101), .Y(n_508) );
AND2x2_ASAP7_75t_L g169 ( .A(n_102), .B(n_168), .Y(n_169) );
OAI321xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_427), .A3(n_434), .B1(n_437), .B2(n_438), .C(n_441), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_105), .B(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_107), .B1(n_110), .B2(n_111), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22x1_ASAP7_75t_SL g458 ( .A1(n_110), .A2(n_459), .B1(n_462), .B2(n_728), .Y(n_458) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_111), .A2(n_463), .B1(n_743), .B2(n_744), .Y(n_742) );
OR3x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_325), .C(n_390), .Y(n_111) );
NAND4xp25_ASAP7_75t_SL g112 ( .A(n_113), .B(n_266), .C(n_292), .D(n_315), .Y(n_112) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_194), .B1(n_235), .B2(n_242), .C(n_258), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_115), .A2(n_259), .B1(n_283), .B2(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_170), .Y(n_115) );
INVx1_ASAP7_75t_SL g319 ( .A(n_116), .Y(n_319) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_150), .Y(n_116) );
OR2x2_ASAP7_75t_L g240 ( .A(n_117), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g261 ( .A(n_117), .B(n_171), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_117), .B(n_181), .Y(n_274) );
AND2x2_ASAP7_75t_L g291 ( .A(n_117), .B(n_150), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_117), .B(n_238), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_117), .B(n_290), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_117), .B(n_170), .Y(n_412) );
AOI211xp5_ASAP7_75t_SL g423 ( .A1(n_117), .A2(n_329), .B(n_424), .C(n_425), .Y(n_423) );
INVx5_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_118), .B(n_171), .Y(n_295) );
AND2x2_ASAP7_75t_L g298 ( .A(n_118), .B(n_172), .Y(n_298) );
OR2x2_ASAP7_75t_L g343 ( .A(n_118), .B(n_171), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_118), .B(n_181), .Y(n_352) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_126), .B(n_147), .Y(n_118) );
INVx3_ASAP7_75t_L g193 ( .A(n_119), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_119), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_119), .A2(n_225), .B(n_233), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_119), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_119), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_119), .B(n_543), .Y(n_542) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_119), .A2(n_547), .B(n_553), .Y(n_546) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_120), .A2(n_174), .B(n_175), .Y(n_173) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_120), .Y(n_182) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g149 ( .A(n_121), .Y(n_149) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_122), .B(n_123), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_135), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_128), .A2(n_472), .B(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_128), .A2(n_168), .B(n_537), .C(n_538), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_128), .A2(n_548), .B(n_549), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
AND2x4_ASAP7_75t_L g153 ( .A(n_129), .B(n_133), .Y(n_153) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g191 ( .A(n_130), .Y(n_191) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_131), .Y(n_146) );
INVx1_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
INVx3_ASAP7_75t_L g141 ( .A(n_132), .Y(n_141) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
INVx1_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx4_ASAP7_75t_SL g167 ( .A(n_133), .Y(n_167) );
BUFx3_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
INVx5_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx3_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_137), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_142), .B(n_144), .Y(n_139) );
INVx5_ASAP7_75t_L g163 ( .A(n_141), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_141), .B(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g255 ( .A(n_143), .Y(n_255) );
INVx2_ASAP7_75t_L g488 ( .A(n_143), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_144), .A2(n_177), .B(n_179), .Y(n_176) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx2_ASAP7_75t_L g525 ( .A(n_149), .Y(n_525) );
INVx5_ASAP7_75t_SL g241 ( .A(n_150), .Y(n_241) );
AND2x2_ASAP7_75t_L g260 ( .A(n_150), .B(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_150), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g346 ( .A(n_150), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g378 ( .A(n_150), .B(n_181), .Y(n_378) );
OR2x2_ASAP7_75t_L g384 ( .A(n_150), .B(n_274), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_150), .B(n_334), .Y(n_393) );
OR2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_169), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B(n_168), .Y(n_151) );
BUFx2_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_156), .A2(n_167), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_156), .A2(n_167), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_156), .A2(n_167), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_156), .A2(n_167), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_156), .A2(n_167), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_156), .A2(n_167), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_156), .A2(n_167), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_162), .C(n_164), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_164), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_159), .A2(n_475), .B(n_476), .C(n_477), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_159), .A2(n_477), .B(n_551), .C(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_163), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g252 ( .A(n_163), .Y(n_252) );
OAI22xp33_ASAP7_75t_L g530 ( .A1(n_163), .A2(n_188), .B1(n_531), .B2(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_163), .A2(n_216), .B(n_540), .C(n_541), .Y(n_539) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g256 ( .A(n_165), .Y(n_256) );
INVx1_ASAP7_75t_L g500 ( .A(n_165), .Y(n_500) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_168), .A2(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_168), .A2(n_484), .B(n_491), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_181), .Y(n_170) );
AND2x2_ASAP7_75t_L g275 ( .A(n_171), .B(n_241), .Y(n_275) );
INVx1_ASAP7_75t_SL g288 ( .A(n_171), .Y(n_288) );
OR2x2_ASAP7_75t_L g323 ( .A(n_171), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g329 ( .A(n_171), .B(n_181), .Y(n_329) );
AND2x2_ASAP7_75t_L g387 ( .A(n_171), .B(n_238), .Y(n_387) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_172), .B(n_241), .Y(n_314) );
INVx3_ASAP7_75t_L g238 ( .A(n_181), .Y(n_238) );
OR2x2_ASAP7_75t_L g280 ( .A(n_181), .B(n_241), .Y(n_280) );
AND2x2_ASAP7_75t_L g290 ( .A(n_181), .B(n_288), .Y(n_290) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_181), .Y(n_338) );
AND2x2_ASAP7_75t_L g347 ( .A(n_181), .B(n_261), .Y(n_347) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_192), .Y(n_181) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_182), .A2(n_494), .B(n_501), .Y(n_493) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_182), .A2(n_503), .B(n_509), .Y(n_502) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_182), .A2(n_513), .B(n_520), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_187), .A2(n_228), .B(n_229), .C(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_188), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_188), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g216 ( .A(n_191), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_191), .B(n_530), .Y(n_529) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_193), .A2(n_248), .B(n_257), .Y(n_247) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_194), .A2(n_364), .B1(n_366), .B2(n_368), .C(n_371), .Y(n_363) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
AND2x2_ASAP7_75t_L g337 ( .A(n_196), .B(n_318), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_196), .B(n_396), .Y(n_400) );
OR2x2_ASAP7_75t_L g421 ( .A(n_196), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_196), .B(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx5_ASAP7_75t_L g268 ( .A(n_197), .Y(n_268) );
AND2x2_ASAP7_75t_L g345 ( .A(n_197), .B(n_208), .Y(n_345) );
AND2x2_ASAP7_75t_L g406 ( .A(n_197), .B(n_285), .Y(n_406) );
AND2x2_ASAP7_75t_L g419 ( .A(n_197), .B(n_238), .Y(n_419) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_204), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_222), .Y(n_206) );
AND2x4_ASAP7_75t_L g245 ( .A(n_207), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g264 ( .A(n_207), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
AND2x2_ASAP7_75t_L g340 ( .A(n_207), .B(n_318), .Y(n_340) );
AND2x2_ASAP7_75t_L g350 ( .A(n_207), .B(n_268), .Y(n_350) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_207), .Y(n_358) );
AND2x2_ASAP7_75t_L g370 ( .A(n_207), .B(n_247), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_207), .B(n_302), .Y(n_374) );
AND2x2_ASAP7_75t_L g411 ( .A(n_207), .B(n_406), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_207), .B(n_285), .Y(n_422) );
OR2x2_ASAP7_75t_L g424 ( .A(n_207), .B(n_360), .Y(n_424) );
INVx5_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g310 ( .A(n_208), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g320 ( .A(n_208), .B(n_265), .Y(n_320) );
AND2x2_ASAP7_75t_L g332 ( .A(n_208), .B(n_247), .Y(n_332) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_208), .Y(n_362) );
AND2x4_ASAP7_75t_L g396 ( .A(n_208), .B(n_246), .Y(n_396) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_212), .B(n_217), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_218), .B(n_436), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_221), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx2_ASAP7_75t_L g244 ( .A(n_222), .Y(n_244) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g285 ( .A(n_223), .Y(n_285) );
AND2x2_ASAP7_75t_L g318 ( .A(n_223), .B(n_247), .Y(n_318) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g265 ( .A(n_224), .B(n_247), .Y(n_265) );
BUFx2_ASAP7_75t_L g311 ( .A(n_224), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g519 ( .A(n_231), .Y(n_519) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_237), .B(n_319), .Y(n_398) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_238), .B(n_261), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_238), .B(n_241), .Y(n_300) );
AND2x2_ASAP7_75t_L g355 ( .A(n_238), .B(n_291), .Y(n_355) );
AOI221xp5_ASAP7_75t_SL g292 ( .A1(n_239), .A2(n_293), .B1(n_301), .B2(n_303), .C(n_307), .Y(n_292) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g287 ( .A(n_240), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g328 ( .A(n_240), .B(n_329), .Y(n_328) );
OAI321xp33_ASAP7_75t_L g335 ( .A1(n_240), .A2(n_294), .A3(n_336), .B1(n_338), .B2(n_339), .C(n_341), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_241), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_244), .B(n_396), .Y(n_414) );
AND2x2_ASAP7_75t_L g301 ( .A(n_245), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_245), .B(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
AND2x2_ASAP7_75t_L g284 ( .A(n_246), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_246), .B(n_359), .Y(n_389) );
INVx1_ASAP7_75t_L g426 ( .A(n_246), .Y(n_426) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_255), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g477 ( .A(n_256), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B(n_263), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_260), .A2(n_370), .B(n_419), .C(n_420), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_261), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_261), .B(n_299), .Y(n_365) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_265), .B(n_268), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_265), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_265), .B(n_350), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_269), .B1(n_281), .B2(n_286), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g282 ( .A(n_268), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g305 ( .A(n_268), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g317 ( .A(n_268), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_268), .B(n_311), .Y(n_353) );
OR2x2_ASAP7_75t_L g360 ( .A(n_268), .B(n_285), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_268), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g410 ( .A(n_268), .B(n_396), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .B1(n_276), .B2(n_278), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g316 ( .A(n_271), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_274), .A2(n_289), .B1(n_357), .B2(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g404 ( .A(n_275), .Y(n_404) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_279), .A2(n_316), .B1(n_319), .B2(n_320), .C(n_321), .Y(n_315) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g294 ( .A(n_280), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_284), .B(n_350), .Y(n_382) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_285), .Y(n_302) );
INVx1_ASAP7_75t_L g306 ( .A(n_285), .Y(n_306) );
NAND2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g324 ( .A(n_291), .Y(n_324) );
AND2x2_ASAP7_75t_L g333 ( .A(n_291), .B(n_334), .Y(n_333) );
NAND2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx2_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g377 ( .A(n_298), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_301), .A2(n_327), .B1(n_330), .B2(n_333), .C(n_335), .Y(n_326) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_305), .B(n_362), .Y(n_361) );
AOI21xp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_309), .B(n_312), .Y(n_307) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_312), .Y(n_409) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
OR2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g372 ( .A(n_317), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_317), .B(n_377), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_320), .B(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NAND4xp25_ASAP7_75t_L g325 ( .A(n_326), .B(n_344), .C(n_363), .D(n_376), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g334 ( .A(n_329), .Y(n_334) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g367 ( .A(n_338), .B(n_343), .Y(n_367) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B(n_348), .C(n_356), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_346), .A2(n_388), .B(n_416), .C(n_423), .Y(n_415) );
INVx1_ASAP7_75t_SL g375 ( .A(n_347), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_353), .B2(n_354), .Y(n_348) );
INVx1_ASAP7_75t_L g379 ( .A(n_353), .Y(n_379) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_359), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_359), .B(n_370), .Y(n_403) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g380 ( .A(n_370), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_375), .Y(n_371) );
INVxp33_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI322xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .A3(n_380), .B1(n_381), .B2(n_383), .C1(n_385), .C2(n_388), .Y(n_376) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g390 ( .A(n_391), .B(n_408), .C(n_415), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B1(n_397), .B2(n_399), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g407 ( .A(n_396), .Y(n_407) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_413), .Y(n_408) );
NAND2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g440 ( .A(n_429), .Y(n_440) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_429), .Y(n_443) );
BUFx2_ASAP7_75t_L g455 ( .A(n_429), .Y(n_455) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_430), .B(n_731), .Y(n_747) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g730 ( .A(n_431), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g437 ( .A(n_434), .Y(n_437) );
NAND2xp33_ASAP7_75t_L g749 ( .A(n_439), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
CKINVDCx6p67_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_449), .A2(n_450), .B(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_SL g750 ( .A(n_449), .B(n_451), .Y(n_750) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g743 ( .A(n_460), .Y(n_743) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_683), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_595), .C(n_633), .D(n_654), .E(n_671), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_567), .C(n_588), .Y(n_465) );
OAI221xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_510), .B1(n_534), .B2(n_554), .C(n_558), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_480), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_469), .B(n_556), .Y(n_575) );
OR2x2_ASAP7_75t_L g602 ( .A(n_469), .B(n_493), .Y(n_602) );
AND2x2_ASAP7_75t_L g616 ( .A(n_469), .B(n_493), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_469), .B(n_483), .Y(n_630) );
AND2x2_ASAP7_75t_L g668 ( .A(n_469), .B(n_632), .Y(n_668) );
AND2x2_ASAP7_75t_L g697 ( .A(n_469), .B(n_607), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_469), .B(n_579), .Y(n_714) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g594 ( .A(n_470), .B(n_492), .Y(n_594) );
BUFx3_ASAP7_75t_L g619 ( .A(n_470), .Y(n_619) );
AND2x2_ASAP7_75t_L g648 ( .A(n_470), .B(n_493), .Y(n_648) );
AND3x2_ASAP7_75t_L g661 ( .A(n_470), .B(n_662), .C(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g584 ( .A(n_480), .Y(n_584) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
AOI32xp33_ASAP7_75t_L g639 ( .A1(n_481), .A2(n_591), .A3(n_640), .B1(n_643), .B2(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g566 ( .A(n_482), .B(n_492), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_482), .B(n_594), .Y(n_637) );
AND2x2_ASAP7_75t_L g644 ( .A(n_482), .B(n_616), .Y(n_644) );
OR2x2_ASAP7_75t_L g650 ( .A(n_482), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_482), .B(n_605), .Y(n_675) );
OR2x2_ASAP7_75t_L g693 ( .A(n_482), .B(n_522), .Y(n_693) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g557 ( .A(n_483), .B(n_502), .Y(n_557) );
INVx2_ASAP7_75t_L g579 ( .A(n_483), .Y(n_579) );
OR2x2_ASAP7_75t_L g601 ( .A(n_483), .B(n_502), .Y(n_601) );
AND2x2_ASAP7_75t_L g606 ( .A(n_483), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_483), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g662 ( .A(n_483), .B(n_556), .Y(n_662) );
INVx1_ASAP7_75t_SL g713 ( .A(n_492), .Y(n_713) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
INVx1_ASAP7_75t_SL g556 ( .A(n_493), .Y(n_556) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_493), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_493), .B(n_642), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_493), .B(n_579), .C(n_697), .Y(n_708) );
INVx2_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_502), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
INVx1_ASAP7_75t_L g643 ( .A(n_511), .Y(n_643) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g561 ( .A(n_512), .B(n_545), .Y(n_561) );
INVx2_ASAP7_75t_L g578 ( .A(n_512), .Y(n_578) );
AND2x2_ASAP7_75t_L g583 ( .A(n_512), .B(n_546), .Y(n_583) );
AND2x2_ASAP7_75t_L g598 ( .A(n_512), .B(n_535), .Y(n_598) );
AND2x2_ASAP7_75t_L g610 ( .A(n_512), .B(n_582), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_521), .B(n_626), .Y(n_625) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_521), .B(n_583), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_521), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_521), .B(n_577), .Y(n_705) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g544 ( .A(n_522), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_522), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g587 ( .A(n_522), .B(n_535), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_522), .B(n_545), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_522), .B(n_653), .Y(n_652) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_526), .B(n_533), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_524), .A2(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_533), .Y(n_573) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_535), .B(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g577 ( .A(n_535), .B(n_578), .Y(n_577) );
INVx3_ASAP7_75t_SL g582 ( .A(n_535), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_535), .B(n_569), .Y(n_635) );
OR2x2_ASAP7_75t_L g645 ( .A(n_535), .B(n_571), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_535), .B(n_613), .Y(n_673) );
OR2x2_ASAP7_75t_L g703 ( .A(n_535), .B(n_545), .Y(n_703) );
AND2x2_ASAP7_75t_L g707 ( .A(n_535), .B(n_546), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_535), .B(n_583), .Y(n_720) );
AND2x2_ASAP7_75t_L g727 ( .A(n_535), .B(n_609), .Y(n_727) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .Y(n_535) );
INVx1_ASAP7_75t_SL g670 ( .A(n_544), .Y(n_670) );
AND2x2_ASAP7_75t_L g609 ( .A(n_545), .B(n_571), .Y(n_609) );
AND2x2_ASAP7_75t_L g623 ( .A(n_545), .B(n_578), .Y(n_623) );
AND2x2_ASAP7_75t_L g626 ( .A(n_545), .B(n_582), .Y(n_626) );
INVx1_ASAP7_75t_L g653 ( .A(n_545), .Y(n_653) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g565 ( .A(n_546), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_555), .A2(n_601), .B(n_725), .C(n_726), .Y(n_724) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g631 ( .A(n_556), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_557), .B(n_574), .Y(n_589) );
AND2x2_ASAP7_75t_L g615 ( .A(n_557), .B(n_616), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_562), .B(n_566), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_560), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g586 ( .A(n_561), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_561), .B(n_582), .Y(n_627) );
AND2x2_ASAP7_75t_L g718 ( .A(n_561), .B(n_569), .Y(n_718) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g591 ( .A(n_565), .B(n_578), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_576), .Y(n_592) );
OAI322xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_575), .A3(n_576), .B1(n_579), .B2(n_580), .C1(n_584), .C2(n_585), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_574), .Y(n_568) );
AND2x2_ASAP7_75t_L g679 ( .A(n_569), .B(n_591), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_569), .B(n_643), .Y(n_725) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g622 ( .A(n_571), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g688 ( .A(n_575), .B(n_601), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_576), .B(n_670), .Y(n_669) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_577), .B(n_609), .Y(n_666) );
AND2x2_ASAP7_75t_L g612 ( .A(n_578), .B(n_582), .Y(n_612) );
AND2x2_ASAP7_75t_L g620 ( .A(n_579), .B(n_621), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_579), .A2(n_658), .B(n_718), .C(n_719), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_580), .A2(n_593), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_582), .B(n_609), .Y(n_649) );
AND2x2_ASAP7_75t_L g655 ( .A(n_582), .B(n_623), .Y(n_655) );
AND2x2_ASAP7_75t_L g689 ( .A(n_582), .B(n_591), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_583), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g699 ( .A(n_583), .Y(n_699) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_587), .A2(n_615), .B1(n_617), .B2(n_622), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_590), .B1(n_592), .B2(n_593), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_589), .A2(n_625), .B1(n_627), .B2(n_628), .Y(n_624) );
INVxp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_594), .A2(n_696), .B1(n_698), .B2(n_700), .C(n_704), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_599), .B(n_603), .C(n_624), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x2_ASAP7_75t_L g665 ( .A(n_601), .B(n_618), .Y(n_665) );
INVx1_ASAP7_75t_L g716 ( .A(n_601), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_602), .A2(n_604), .B1(n_608), .B2(n_611), .C(n_614), .Y(n_603) );
INVx2_ASAP7_75t_SL g658 ( .A(n_602), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g723 ( .A(n_605), .Y(n_723) );
AND2x2_ASAP7_75t_L g647 ( .A(n_606), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g632 ( .A(n_607), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g694 ( .A(n_610), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_618), .B(n_720), .Y(n_719) );
CKINVDCx16_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_L g663 ( .A(n_621), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_622), .A2(n_634), .B(n_636), .C(n_638), .Y(n_633) );
INVx1_ASAP7_75t_L g711 ( .A(n_625), .Y(n_711) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_629), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx2_ASAP7_75t_L g642 ( .A(n_632), .Y(n_642) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_645), .B1(n_646), .B2(n_649), .C1(n_650), .C2(n_652), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g678 ( .A(n_642), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_645), .B(n_699), .Y(n_698) );
NAND2xp33_ASAP7_75t_SL g676 ( .A(n_646), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g651 ( .A(n_648), .Y(n_651) );
AND2x2_ASAP7_75t_L g715 ( .A(n_648), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g681 ( .A(n_651), .B(n_678), .Y(n_681) );
INVx1_ASAP7_75t_L g710 ( .A(n_652), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B(n_659), .C(n_664), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_658), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AOI322xp5_ASAP7_75t_L g709 ( .A1(n_661), .A2(n_689), .A3(n_694), .B1(n_710), .B2(n_711), .C1(n_712), .C2(n_715), .Y(n_709) );
AND2x2_ASAP7_75t_L g696 ( .A(n_662), .B(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_669), .Y(n_664) );
INVxp33_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_676), .B2(n_679), .C(n_680), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND5xp2_ASAP7_75t_L g683 ( .A(n_684), .B(n_695), .C(n_709), .D(n_717), .E(n_721), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B(n_690), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp33_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_697), .A2(n_722), .B(n_723), .C(n_724), .Y(n_721) );
AOI31xp33_ASAP7_75t_L g704 ( .A1(n_699), .A2(n_705), .A3(n_706), .B(n_708), .Y(n_704) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g722 ( .A(n_720), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g744 ( .A(n_729), .Y(n_744) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_737), .Y(n_740) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx3_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
endmodule