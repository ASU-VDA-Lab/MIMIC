module real_jpeg_29287_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_293;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx11_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_1),
.A2(n_44),
.B1(n_47),
.B2(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_44),
.B1(n_77),
.B2(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_77),
.B1(n_78),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_2),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_126),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_126),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_2),
.A2(n_47),
.B1(n_51),
.B2(n_126),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_29),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_4),
.A2(n_29),
.B(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_153),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_4),
.A2(n_10),
.B(n_47),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_120),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_4),
.A2(n_89),
.B1(n_142),
.B2(n_244),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_7),
.A2(n_77),
.B1(n_78),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_7),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_155),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_155),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_7),
.A2(n_47),
.B1(n_51),
.B2(n_155),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_8),
.A2(n_47),
.B1(n_51),
.B2(n_58),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_9),
.A2(n_40),
.B1(n_47),
.B2(n_51),
.Y(n_139)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_11),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_11),
.A2(n_77),
.B1(n_78),
.B2(n_149),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_149),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_11),
.A2(n_47),
.B1(n_51),
.B2(n_149),
.Y(n_236)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_38),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_14),
.A2(n_38),
.B1(n_47),
.B2(n_51),
.Y(n_172)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_102),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_86),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_60),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_25),
.B(n_70),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_25),
.A2(n_33),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_25),
.A2(n_33),
.B1(n_148),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_25),
.A2(n_33),
.B1(n_181),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_27),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_27),
.B(n_35),
.Y(n_197)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_29),
.A2(n_30),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_29),
.B(n_74),
.Y(n_169)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_30),
.A2(n_81),
.B1(n_152),
.B2(n_169),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_30),
.A2(n_34),
.A3(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_194)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_33),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_35),
.A2(n_50),
.B(n_153),
.C(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_37),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_42),
.A2(n_55),
.B(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_45),
.B(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_55),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_46),
.A2(n_55),
.B1(n_97),
.B2(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_46),
.A2(n_53),
.B(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_46),
.A2(n_55),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_46),
.A2(n_55),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_46),
.A2(n_55),
.B1(n_203),
.B2(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_46),
.B(n_153),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_90),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_51),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_64),
.B(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_84),
.B2(n_85),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_67),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_67),
.A2(n_69),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_83),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_72),
.A2(n_124),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_72),
.B(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_72),
.A2(n_124),
.B1(n_125),
.B2(n_161),
.Y(n_279)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.C(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_73),
.B(n_100),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_73),
.A2(n_80),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_78),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g152 ( 
.A(n_78),
.B(n_153),
.CON(n_152),
.SN(n_152)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_80),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B(n_99),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_99),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_88),
.A2(n_96),
.B1(n_106),
.B2(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_93),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_89),
.A2(n_90),
.B1(n_139),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_89),
.A2(n_115),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_89),
.A2(n_142),
.B1(n_236),
.B2(n_244),
.Y(n_243)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_92),
.A2(n_113),
.B(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_94),
.A2(n_141),
.B(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_96),
.Y(n_296)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_108),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_103),
.B(n_107),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_108),
.A2(n_109),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_119),
.C(n_122),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_110),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_111),
.B(n_117),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_116),
.A2(n_193),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_119),
.Y(n_293)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_127),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_299),
.B(n_304),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_286),
.B(n_298),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_185),
.B(n_267),
.C(n_285),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_173),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_134),
.B(n_173),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_156),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_136),
.B(n_143),
.C(n_156),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_137),
.B(n_138),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_142),
.B(n_153),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_151),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_167),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_158),
.B(n_163),
.C(n_167),
.Y(n_283)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_166),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_170),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_179),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_174),
.A2(n_175),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_266),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_259),
.B(n_265),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_214),
.B(n_258),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_205),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_189),
.B(n_205),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.C(n_201),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_190),
.A2(n_191),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_194),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_212),
.C(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_252),
.B(n_257),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_232),
.B(n_251),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_240),
.B(n_250),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_283),
.B2(n_284),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.C(n_284),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_278),
.C(n_281),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.C(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);


endmodule