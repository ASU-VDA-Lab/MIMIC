module fake_jpeg_16631_n_50 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_50);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_50;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_11),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_6),
.B(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_0),
.B1(n_12),
.B2(n_17),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2x1_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_29),
.B1(n_36),
.B2(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_37),
.CI(n_38),
.CON(n_46),
.SN(n_46)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_36),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_46),
.C(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_43),
.Y(n_50)
);


endmodule