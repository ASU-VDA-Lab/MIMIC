module fake_ariane_1938_n_1610 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1610);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1610;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_246;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g171 ( 
.A(n_33),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_19),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_72),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_42),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_14),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_75),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_4),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_129),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_28),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_45),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_122),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_68),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_63),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_36),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_66),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_89),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_20),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_133),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_67),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_34),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_41),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_22),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_69),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_103),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_18),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_35),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_116),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_77),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_137),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_119),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_16),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_147),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_80),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_148),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_28),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_30),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_139),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_48),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_79),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_102),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_51),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_92),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_78),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_88),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_114),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_51),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_54),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_112),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_21),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_149),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_157),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_117),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_54),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_155),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_156),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_105),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_22),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_42),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_29),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_108),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_58),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_23),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_144),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_24),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_154),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_128),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

BUFx8_ASAP7_75t_SL g286 ( 
.A(n_106),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_138),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_62),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_76),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_71),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_135),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_95),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_140),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_52),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_91),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_6),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_50),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_168),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_57),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_90),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_146),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_7),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_50),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_94),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_25),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_33),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_169),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_49),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_19),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_30),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_83),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_12),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_27),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_85),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_61),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_64),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_12),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_23),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_158),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_109),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_73),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_121),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_44),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_143),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_130),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_52),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_163),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_49),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_46),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_7),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_44),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_40),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_21),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_93),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_98),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_87),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_127),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_6),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_55),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_151),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_113),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_74),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_165),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_36),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_201),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_201),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_210),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_308),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_259),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_259),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_200),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_210),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_188),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_231),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_231),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_251),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_280),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_327),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_174),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_263),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_251),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_180),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_262),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_181),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_294),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_176),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_171),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_281),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_294),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_178),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_200),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_178),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_219),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_203),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_219),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_303),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_281),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_298),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_183),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_298),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_205),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_223),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_292),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_183),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_228),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_236),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_185),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_241),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_247),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_182),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_248),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_174),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_303),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_185),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_186),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_255),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_195),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_267),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_174),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_186),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_179),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_278),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_282),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_297),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_299),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_310),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_321),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_184),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_179),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_268),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_195),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_316),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_186),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_204),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_266),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_191),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_193),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_194),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_209),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_204),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_213),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_204),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_214),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_279),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_208),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_286),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g442 ( 
.A(n_216),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_365),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_372),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_173),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_351),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_380),
.A2(n_218),
.B(n_217),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_348),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_208),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_348),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_349),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_432),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_351),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_425),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_222),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_349),
.A2(n_224),
.B(n_220),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_368),
.Y(n_475)
);

BUFx8_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_356),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_422),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_229),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_350),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_352),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_433),
.B(n_222),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_438),
.A2(n_249),
.B(n_238),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_350),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_354),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_438),
.B(n_250),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_355),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_386),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_356),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_355),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_357),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_406),
.A2(n_271),
.B(n_265),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_353),
.B(n_276),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_357),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_358),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_378),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_381),
.Y(n_505)
);

BUFx8_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_358),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_359),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_359),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_366),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_366),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_374),
.B(n_277),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_404),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_442),
.B(n_173),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_367),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_391),
.B(n_287),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_367),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_400),
.B(n_288),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_369),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_362),
.B(n_192),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_447),
.A2(n_364),
.B1(n_392),
.B2(n_363),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_SL g523 ( 
.A1(n_472),
.A2(n_439),
.B(n_408),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_452),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_468),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_492),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_472),
.B(n_411),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_472),
.B(n_411),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_468),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_468),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_468),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_468),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_444),
.Y(n_537)
);

AO21x2_ASAP7_75t_L g538 ( 
.A1(n_456),
.A2(n_302),
.B(n_300),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_468),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_487),
.B(n_428),
.Y(n_542)
);

BUFx6f_ASAP7_75t_SL g543 ( 
.A(n_513),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_468),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_467),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_501),
.B(n_360),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_463),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_447),
.A2(n_364),
.B1(n_392),
.B2(n_363),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_489),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_487),
.Y(n_552)
);

AND3x2_ASAP7_75t_L g553 ( 
.A(n_454),
.B(n_441),
.C(n_409),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_487),
.B(n_389),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_501),
.B(n_361),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_500),
.B(n_406),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_467),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_513),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_491),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_488),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_514),
.B(n_428),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_491),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_514),
.B(n_429),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_491),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_471),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_471),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_520),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_412),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_489),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_491),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_489),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_479),
.B(n_429),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_447),
.B(n_435),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_489),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_489),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_513),
.Y(n_584)
);

XNOR2x2_ASAP7_75t_R g585 ( 
.A(n_466),
.B(n_440),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_446),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_501),
.B(n_435),
.Y(n_589)
);

NOR2x1p5_ASAP7_75t_L g590 ( 
.A(n_479),
.B(n_266),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_501),
.B(n_388),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_447),
.B(n_469),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_504),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_474),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_501),
.B(n_393),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_496),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_447),
.B(n_437),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_469),
.B(n_430),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_508),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_473),
.A2(n_373),
.B1(n_407),
.B2(n_426),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_478),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_513),
.B(n_401),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_469),
.B(n_410),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_508),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_478),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_478),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_513),
.B(n_454),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_481),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_511),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_496),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_520),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_473),
.A2(n_396),
.B1(n_403),
.B2(n_254),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_481),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_446),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_481),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_481),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_483),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_483),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_483),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_453),
.B(n_329),
.C(n_319),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_483),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_484),
.B(n_413),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_459),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_453),
.B(n_329),
.C(n_319),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_511),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_511),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_495),
.B(n_516),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_495),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_473),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_470),
.B(n_459),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_460),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_460),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_466),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_495),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_460),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_460),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_511),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_511),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_500),
.B(n_414),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_461),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_511),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_461),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_511),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_486),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_516),
.A2(n_230),
.B1(n_270),
.B2(n_272),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_486),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_461),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_512),
.B(n_390),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_461),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_449),
.B(n_176),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_462),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_470),
.B(n_187),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_511),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_512),
.B(n_394),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_527),
.B(n_476),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_545),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_546),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_552),
.B(n_470),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_552),
.B(n_476),
.Y(n_662)
);

INVx6_ASAP7_75t_L g663 ( 
.A(n_626),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_528),
.B(n_476),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_614),
.B(n_382),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_625),
.B(n_518),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_567),
.B(n_482),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_572),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_554),
.A2(n_476),
.B1(n_493),
.B2(n_486),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_557),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_542),
.B(n_486),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_572),
.B(n_505),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_560),
.B(n_486),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_625),
.B(n_506),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_651),
.B(n_506),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_614),
.B(n_385),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_657),
.B(n_506),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_642),
.B(n_506),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_557),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_584),
.B(n_506),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_402),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_584),
.B(n_493),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_603),
.B(n_189),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_642),
.B(n_630),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_563),
.B(n_505),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_526),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_632),
.A2(n_642),
.B1(n_592),
.B2(n_556),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_565),
.B(n_482),
.Y(n_688)
);

OAI221xp5_ASAP7_75t_L g689 ( 
.A1(n_523),
.A2(n_274),
.B1(n_331),
.B2(n_333),
.C(n_335),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_554),
.B(n_395),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_554),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_556),
.B(n_475),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_556),
.B(n_581),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_579),
.B(n_190),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_640),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_556),
.B(n_475),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_554),
.B(n_397),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_581),
.B(n_477),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_581),
.B(n_477),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_598),
.B(n_196),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_543),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_567),
.B(n_480),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_593),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_606),
.B(n_480),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_551),
.B(n_497),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_640),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_569),
.B(n_449),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_640),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_551),
.B(n_497),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_551),
.B(n_497),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_599),
.B(n_497),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_573),
.B(n_497),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_573),
.B(n_515),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_610),
.B(n_515),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_573),
.B(n_515),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_543),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_591),
.B(n_515),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_522),
.B(n_202),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_537),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_575),
.B(n_580),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_595),
.B(n_515),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_550),
.A2(n_335),
.B1(n_336),
.B2(n_334),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_575),
.B(n_451),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_473),
.B1(n_230),
.B2(n_315),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_576),
.B(n_336),
.C(n_331),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_648),
.A2(n_315),
.B1(n_326),
.B2(n_270),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_597),
.B(n_264),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_526),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_548),
.B(n_455),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_615),
.B(n_455),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_549),
.B(n_457),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_597),
.B(n_264),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_613),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_549),
.B(n_457),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_633),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_589),
.B(n_458),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_558),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_547),
.B(n_555),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_613),
.B(n_605),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_632),
.A2(n_473),
.B1(n_465),
.B2(n_462),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_634),
.A2(n_473),
.B1(n_465),
.B2(n_462),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_562),
.B(n_571),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_562),
.B(n_269),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_634),
.A2(n_462),
.B1(n_465),
.B2(n_464),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_571),
.B(n_464),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_582),
.B(n_269),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_559),
.B(n_494),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_655),
.B(n_502),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_569),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_588),
.B(n_502),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_SL g752 ( 
.A(n_543),
.B(n_175),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_647),
.B(n_324),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_635),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_636),
.B(n_507),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_635),
.B(n_507),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_590),
.B(n_553),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_638),
.B(n_510),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_623),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_638),
.B(n_510),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_639),
.B(n_517),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_641),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_641),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_585),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_588),
.B(n_517),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_647),
.B(n_398),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_604),
.Y(n_767)
);

AND2x2_ASAP7_75t_SL g768 ( 
.A(n_639),
.B(n_317),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_643),
.B(n_519),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_643),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_645),
.B(n_519),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_650),
.B(n_465),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_650),
.B(n_652),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_652),
.B(n_485),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_654),
.B(n_485),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_L g776 ( 
.A(n_627),
.B(n_485),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_654),
.B(n_485),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_649),
.B(n_324),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_631),
.B(n_211),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_SL g780 ( 
.A(n_525),
.B(n_221),
.C(n_212),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_637),
.B(n_498),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_641),
.B(n_330),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_531),
.B(n_237),
.C(n_232),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_604),
.Y(n_784)
);

OAI22xp33_ASAP7_75t_L g785 ( 
.A1(n_649),
.A2(n_509),
.B1(n_503),
.B2(n_498),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_637),
.B(n_239),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_417),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_531),
.B(n_240),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_608),
.B(n_498),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_609),
.B(n_498),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_695),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_690),
.B(n_414),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_666),
.B(n_609),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_660),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_724),
.A2(n_618),
.B1(n_620),
.B2(n_621),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_724),
.A2(n_618),
.B1(n_620),
.B2(n_621),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_701),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_768),
.B(n_641),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_768),
.B(n_641),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_691),
.B(n_503),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_658),
.A2(n_656),
.B1(n_628),
.B2(n_529),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_726),
.A2(n_611),
.B1(n_622),
.B2(n_624),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_687),
.B(n_531),
.Y(n_803)
);

AND2x2_ASAP7_75t_SL g804 ( 
.A(n_687),
.B(n_318),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_701),
.Y(n_805)
);

AND2x2_ASAP7_75t_SL g806 ( 
.A(n_669),
.B(n_323),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_684),
.B(n_720),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_695),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_664),
.A2(n_656),
.B1(n_628),
.B2(n_533),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_663),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_663),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_711),
.B(n_611),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_664),
.B(n_540),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_663),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_671),
.B(n_540),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_766),
.B(n_616),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_685),
.B(n_540),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_675),
.A2(n_677),
.B(n_671),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_686),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_665),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_SL g821 ( 
.A(n_783),
.B(n_256),
.C(n_244),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_750),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_695),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_766),
.B(n_619),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_668),
.B(n_415),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_690),
.B(n_415),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_676),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_691),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_735),
.B(n_525),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_703),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_739),
.A2(n_533),
.B1(n_536),
.B2(n_541),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_749),
.B(n_544),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_SL g833 ( 
.A(n_727),
.B(n_258),
.C(n_257),
.Y(n_833)
);

BUFx6f_ASAP7_75t_SL g834 ( 
.A(n_733),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_695),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_737),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_688),
.B(n_521),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_706),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

AO22x1_ASAP7_75t_L g840 ( 
.A1(n_764),
.A2(n_261),
.B1(n_312),
.B2(n_307),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_SL g841 ( 
.A(n_693),
.B(n_521),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_754),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_697),
.B(n_416),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_770),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_688),
.B(n_524),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_738),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_701),
.B(n_503),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_681),
.Y(n_848)
);

CKINVDCx6p67_ASAP7_75t_R g849 ( 
.A(n_716),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_728),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_706),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_755),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_757),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_723),
.A2(n_564),
.B1(n_646),
.B2(n_644),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_698),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_706),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_697),
.B(n_416),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_708),
.B(n_530),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_699),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_726),
.A2(n_503),
.B1(n_509),
.B2(n_538),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_702),
.B(n_418),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_661),
.B(n_532),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_716),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_674),
.B(n_532),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_759),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_748),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_779),
.B(n_786),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_707),
.B(n_419),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_708),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_767),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_667),
.B(n_420),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_756),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_758),
.Y(n_874)
);

O2A1O1Ixp5_ASAP7_75t_L g875 ( 
.A1(n_682),
.A2(n_534),
.B(n_629),
.C(n_535),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_760),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_761),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_659),
.Y(n_878)
);

BUFx12f_ASAP7_75t_L g879 ( 
.A(n_787),
.Y(n_879)
);

INVx5_ASAP7_75t_L g880 ( 
.A(n_716),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_708),
.B(n_535),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_762),
.B(n_539),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_704),
.B(n_561),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_762),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_717),
.A2(n_490),
.B(n_499),
.C(n_456),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_769),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_771),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_729),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_787),
.B(n_421),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_670),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_751),
.B(n_765),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_692),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_787),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_696),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_763),
.B(n_566),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_719),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_765),
.B(n_568),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_679),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_789),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_790),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_740),
.B(n_423),
.C(n_285),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_731),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_734),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_763),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_746),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_772),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_774),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_775),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_700),
.B(n_574),
.Y(n_909)
);

CKINVDCx8_ASAP7_75t_R g910 ( 
.A(n_717),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_721),
.B(n_577),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_705),
.A2(n_710),
.B(n_709),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_743),
.Y(n_913)
);

NOR2x2_ASAP7_75t_L g914 ( 
.A(n_722),
.B(n_577),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_777),
.Y(n_915)
);

NOR2x2_ASAP7_75t_L g916 ( 
.A(n_718),
.B(n_725),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_678),
.B(n_578),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_SL g918 ( 
.A1(n_736),
.A2(n_586),
.B(n_583),
.C(n_612),
.Y(n_918)
);

OR2x2_ASAP7_75t_SL g919 ( 
.A(n_780),
.B(n_369),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_683),
.A2(n_509),
.B1(n_538),
.B2(n_222),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_781),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_773),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_730),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_SL g924 ( 
.A(n_783),
.B(n_295),
.C(n_275),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_732),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_714),
.B(n_596),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_689),
.B(n_752),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_694),
.A2(n_607),
.B(n_602),
.C(n_601),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_736),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_600),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_929),
.B(n_662),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_896),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_880),
.B(n_797),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_891),
.A2(n_713),
.B(n_712),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_794),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_867),
.A2(n_744),
.B(n_747),
.C(n_788),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_812),
.A2(n_715),
.B(n_785),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_818),
.A2(n_776),
.B(n_788),
.C(n_778),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_817),
.A2(n_753),
.B(n_680),
.C(n_673),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_837),
.A2(n_782),
.B(n_741),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_SL g941 ( 
.A(n_834),
.B(n_745),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_845),
.A2(n_741),
.B(n_742),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_SL g943 ( 
.A(n_819),
.B(n_304),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_804),
.A2(n_745),
.B1(n_742),
.B2(n_607),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_822),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_804),
.A2(n_602),
.B1(n_601),
.B2(n_314),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_857),
.B(n_305),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_922),
.A2(n_347),
.B1(n_337),
.B2(n_340),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_839),
.A2(n_339),
.B(n_325),
.C(n_376),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_L g950 ( 
.A(n_880),
.B(n_850),
.Y(n_950)
);

CKINVDCx6p67_ASAP7_75t_R g951 ( 
.A(n_834),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_910),
.B(n_839),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_912),
.A2(n_538),
.B(n_617),
.Y(n_953)
);

BUFx8_ASAP7_75t_L g954 ( 
.A(n_820),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_829),
.A2(n_448),
.B(n_371),
.C(n_322),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_848),
.B(n_198),
.Y(n_956)
);

AO32x1_ASAP7_75t_L g957 ( 
.A1(n_854),
.A2(n_450),
.A3(n_445),
.B1(n_443),
.B2(n_653),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_880),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_827),
.B(n_309),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_830),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_912),
.A2(n_617),
.B(n_587),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_807),
.A2(n_617),
.B(n_587),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_849),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_866),
.A2(n_338),
.B1(n_343),
.B2(n_344),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_893),
.B(n_797),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_880),
.Y(n_966)
);

NOR2x1_ASAP7_75t_L g967 ( 
.A(n_805),
.B(n_328),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_806),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_872),
.B(n_587),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_813),
.A2(n_448),
.B(n_450),
.C(n_445),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_904),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_792),
.B(n_0),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_826),
.B(n_4),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_829),
.A2(n_448),
.B(n_445),
.C(n_443),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_828),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_897),
.A2(n_587),
.B(n_617),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_828),
.B(n_172),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_874),
.B(n_653),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_826),
.B(n_206),
.Y(n_979)
);

AO21x1_ASAP7_75t_L g980 ( 
.A1(n_841),
.A2(n_450),
.B(n_445),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_843),
.B(n_9),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_852),
.B(n_10),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_883),
.A2(n_253),
.B(n_207),
.Y(n_983)
);

BUFx8_ASAP7_75t_L g984 ( 
.A(n_879),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_843),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_SL g986 ( 
.A1(n_918),
.A2(n_443),
.B(n_11),
.C(n_13),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_853),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_825),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_876),
.B(n_10),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_877),
.B(n_11),
.Y(n_990)
);

NOR2xp67_ASAP7_75t_SL g991 ( 
.A(n_805),
.B(n_225),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_927),
.B(n_226),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_865),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_886),
.A2(n_296),
.B1(n_227),
.B2(n_233),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_853),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_887),
.B(n_653),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_923),
.B(n_653),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_889),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_793),
.A2(n_301),
.B1(n_234),
.B2(n_235),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_806),
.B(n_653),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_846),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_925),
.B(n_242),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_791),
.Y(n_1003)
);

AOI33xp33_ASAP7_75t_L g1004 ( 
.A1(n_868),
.A2(n_443),
.A3(n_15),
.B1(n_18),
.B2(n_24),
.B3(n_26),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_802),
.B(n_13),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_885),
.A2(n_653),
.B(n_346),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_SL g1007 ( 
.A(n_821),
.B(n_293),
.C(n_245),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_802),
.B(n_29),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_SL g1009 ( 
.A(n_924),
.B(n_291),
.C(n_243),
.Y(n_1009)
);

OA22x2_ASAP7_75t_L g1010 ( 
.A1(n_861),
.A2(n_290),
.B1(n_246),
.B2(n_252),
.Y(n_1010)
);

OAI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_800),
.A2(n_283),
.B1(n_289),
.B2(n_284),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_800),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_888),
.B(n_177),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_924),
.B(n_260),
.C(n_306),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_892),
.B(n_31),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_864),
.A2(n_909),
.B(n_902),
.C(n_903),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_800),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_871),
.B(n_31),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_875),
.A2(n_197),
.B(n_177),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_870),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_863),
.Y(n_1021)
);

INVxp33_ASAP7_75t_L g1022 ( 
.A(n_901),
.Y(n_1022)
);

AOI221x1_ASAP7_75t_L g1023 ( 
.A1(n_841),
.A2(n_446),
.B1(n_215),
.B2(n_197),
.C(n_177),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_916),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_873),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_847),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_878),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_836),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_1028)
);

BUFx4f_ASAP7_75t_SL g1029 ( 
.A(n_810),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_SL g1030 ( 
.A1(n_798),
.A2(n_37),
.B(n_38),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_916),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_909),
.A2(n_446),
.B(n_197),
.C(n_177),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_905),
.A2(n_446),
.B(n_197),
.C(n_177),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_842),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_894),
.B(n_39),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_871),
.B(n_39),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_844),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_855),
.B(n_40),
.Y(n_1038)
);

OAI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_859),
.A2(n_43),
.B(n_47),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_833),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_811),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_913),
.B(n_48),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_814),
.B(n_53),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_847),
.B(n_53),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_862),
.A2(n_197),
.B(n_177),
.C(n_55),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_860),
.B(n_197),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_937),
.A2(n_815),
.B(n_918),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_995),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_992),
.A2(n_798),
.B(n_799),
.C(n_901),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_936),
.A2(n_799),
.B(n_862),
.C(n_860),
.Y(n_1050)
);

AOI211x1_ASAP7_75t_L g1051 ( 
.A1(n_1028),
.A2(n_840),
.B(n_803),
.C(n_908),
.Y(n_1051)
);

AO221x2_ASAP7_75t_L g1052 ( 
.A1(n_1028),
.A2(n_914),
.B1(n_919),
.B2(n_906),
.C(n_930),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_963),
.B(n_791),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_934),
.A2(n_926),
.B(n_832),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_1008),
.A2(n_914),
.B1(n_803),
.B2(n_900),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_988),
.B(n_899),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_935),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_980),
.A2(n_885),
.A3(n_917),
.B(n_911),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_1045),
.A2(n_928),
.B(n_907),
.C(n_915),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_968),
.A2(n_816),
.B1(n_824),
.B2(n_831),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_948),
.A2(n_928),
.B(n_882),
.C(n_881),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1016),
.A2(n_847),
.B(n_791),
.Y(n_1062)
);

AO21x2_ASAP7_75t_L g1063 ( 
.A1(n_1006),
.A2(n_895),
.B(n_858),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1006),
.A2(n_801),
.B(n_809),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_985),
.B(n_795),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_952),
.B(n_795),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_945),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_941),
.B(n_791),
.Y(n_1068)
);

AND3x2_ASAP7_75t_L g1069 ( 
.A(n_1024),
.B(n_898),
.C(n_890),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_932),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_960),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_998),
.B(n_796),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1031),
.B(n_796),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_SL g1074 ( 
.A1(n_948),
.A2(n_913),
.B(n_856),
.C(n_884),
.Y(n_1074)
);

AOI221x1_ASAP7_75t_L g1075 ( 
.A1(n_1039),
.A2(n_921),
.B1(n_808),
.B2(n_884),
.C(n_823),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_975),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1044),
.A2(n_920),
.B1(n_851),
.B2(n_869),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_1004),
.A2(n_838),
.B(n_808),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_965),
.B(n_869),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_984),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_939),
.A2(n_931),
.B(n_1022),
.C(n_949),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_SL g1082 ( 
.A(n_1021),
.B(n_835),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_959),
.B(n_835),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_946),
.A2(n_59),
.B(n_60),
.Y(n_1084)
);

AO21x2_ASAP7_75t_L g1085 ( 
.A1(n_1033),
.A2(n_81),
.B(n_84),
.Y(n_1085)
);

AOI211x1_ASAP7_75t_L g1086 ( 
.A1(n_972),
.A2(n_86),
.B(n_99),
.C(n_100),
.Y(n_1086)
);

AND3x4_ASAP7_75t_L g1087 ( 
.A(n_950),
.B(n_107),
.C(n_111),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_938),
.A2(n_118),
.B(n_124),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_979),
.B(n_166),
.Y(n_1089)
);

OAI22x1_ASAP7_75t_L g1090 ( 
.A1(n_1040),
.A2(n_125),
.B1(n_131),
.B2(n_134),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_970),
.A2(n_976),
.B(n_962),
.Y(n_1091)
);

CKINVDCx14_ASAP7_75t_R g1092 ( 
.A(n_993),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1012),
.Y(n_1093)
);

NOR4xp25_ASAP7_75t_L g1094 ( 
.A(n_1030),
.B(n_150),
.C(n_955),
.D(n_986),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_974),
.A2(n_1038),
.B(n_989),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_999),
.A2(n_946),
.B1(n_964),
.B2(n_990),
.Y(n_1096)
);

INVx3_ASAP7_75t_SL g1097 ( 
.A(n_951),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_994),
.A2(n_981),
.B(n_973),
.C(n_999),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_956),
.B(n_947),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1044),
.B(n_1000),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_SL g1101 ( 
.A1(n_1036),
.A2(n_1018),
.B(n_994),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_958),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_969),
.A2(n_944),
.B(n_1000),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_969),
.A2(n_944),
.B(n_957),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_957),
.A2(n_1013),
.B(n_978),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_SL g1106 ( 
.A(n_1007),
.B(n_1014),
.C(n_1009),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1011),
.B(n_966),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1015),
.A2(n_1035),
.B(n_996),
.Y(n_1108)
);

AO21x1_ASAP7_75t_L g1109 ( 
.A1(n_1042),
.A2(n_997),
.B(n_978),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_984),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1034),
.B(n_1037),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1017),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_977),
.B(n_982),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_958),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1002),
.A2(n_983),
.B(n_967),
.C(n_971),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_958),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1003),
.A2(n_1026),
.B(n_933),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1027),
.A2(n_1020),
.A3(n_1025),
.B(n_1001),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1029),
.Y(n_1119)
);

AOI211x1_ASAP7_75t_L g1120 ( 
.A1(n_943),
.A2(n_991),
.B(n_1010),
.C(n_1043),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_966),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_L g1122 ( 
.A(n_1041),
.B(n_954),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_942),
.A2(n_940),
.B(n_937),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_985),
.B(n_857),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_985),
.B(n_839),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_942),
.A2(n_940),
.B(n_937),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_988),
.B(n_668),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_988),
.B(n_668),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1005),
.A2(n_804),
.B1(n_806),
.B2(n_768),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_985),
.B(n_857),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_992),
.A2(n_867),
.B(n_658),
.C(n_664),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_988),
.B(n_668),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_953),
.A2(n_1019),
.B(n_961),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_987),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_952),
.B(n_867),
.Y(n_1135)
);

AOI211x1_ASAP7_75t_L g1136 ( 
.A1(n_1028),
.A2(n_972),
.B(n_981),
.C(n_973),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_988),
.B(n_668),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1008),
.A2(n_929),
.B1(n_867),
.B2(n_724),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_1006),
.A2(n_867),
.B(n_818),
.C(n_980),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_985),
.B(n_839),
.Y(n_1140)
);

AOI221x1_ASAP7_75t_L g1141 ( 
.A1(n_1039),
.A2(n_1045),
.B1(n_867),
.B2(n_1005),
.C(n_1006),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_932),
.Y(n_1142)
);

NAND3x1_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_648),
.C(n_952),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_952),
.B(n_728),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_985),
.B(n_857),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1005),
.A2(n_804),
.B1(n_806),
.B2(n_768),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_948),
.A2(n_726),
.B1(n_722),
.B2(n_685),
.C(n_550),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_953),
.A2(n_1019),
.B(n_961),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_952),
.B(n_867),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_945),
.Y(n_1150)
);

AO22x2_ASAP7_75t_L g1151 ( 
.A1(n_1008),
.A2(n_466),
.B1(n_946),
.B2(n_1046),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_988),
.B(n_668),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_992),
.A2(n_867),
.B(n_658),
.C(n_664),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_980),
.A2(n_1023),
.A3(n_1032),
.B(n_942),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_992),
.A2(n_867),
.B(n_658),
.C(n_664),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_958),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1151),
.A2(n_1052),
.B1(n_1146),
.B2(n_1129),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1135),
.B(n_1149),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1096),
.A2(n_1081),
.B(n_1101),
.C(n_1147),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_1049),
.A2(n_1064),
.B(n_1050),
.C(n_1089),
.Y(n_1160)
);

BUFx8_ASAP7_75t_SL g1161 ( 
.A(n_1080),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1123),
.A2(n_1126),
.B(n_1047),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1102),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1124),
.B(n_1130),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_1100),
.B(n_1062),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1054),
.A2(n_1126),
.B(n_1123),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1111),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1151),
.A2(n_1088),
.B1(n_1138),
.B2(n_1090),
.C(n_1084),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1066),
.B(n_1099),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1082),
.B(n_1068),
.Y(n_1170)
);

INVx6_ASAP7_75t_L g1171 ( 
.A(n_1119),
.Y(n_1171)
);

CKINVDCx14_ASAP7_75t_R g1172 ( 
.A(n_1092),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1057),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1145),
.B(n_1076),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1058),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1070),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1109),
.A2(n_1141),
.A3(n_1075),
.B(n_1077),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_SL g1178 ( 
.A1(n_1098),
.A2(n_1095),
.B(n_1146),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1101),
.B(n_1138),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1139),
.A2(n_1129),
.B(n_1088),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1067),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1071),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_1134),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1136),
.A2(n_1144),
.B1(n_1142),
.B2(n_1143),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1095),
.A2(n_1061),
.B(n_1108),
.Y(n_1185)
);

OAI21xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1107),
.A2(n_1094),
.B(n_1074),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1058),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1125),
.B(n_1140),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1059),
.A2(n_1117),
.B(n_1077),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1112),
.B(n_1093),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1056),
.B(n_1113),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1058),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1094),
.A2(n_1060),
.B(n_1115),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_1097),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_1063),
.A2(n_1085),
.B(n_1078),
.Y(n_1195)
);

BUFx4f_ASAP7_75t_SL g1196 ( 
.A(n_1150),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1156),
.A2(n_1121),
.B(n_1083),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1055),
.A2(n_1120),
.B1(n_1128),
.B2(n_1132),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1078),
.A2(n_1127),
.B(n_1137),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1073),
.B(n_1152),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1053),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1114),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1106),
.A2(n_1065),
.B(n_1122),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1112),
.B(n_1093),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1072),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1154),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1051),
.A2(n_1086),
.B1(n_1087),
.B2(n_1110),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1114),
.B(n_1116),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1069),
.B(n_1114),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1116),
.B(n_1048),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1154),
.A2(n_1091),
.B(n_1133),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_1008),
.B2(n_1147),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1111),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1111),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_L g1215 ( 
.A(n_1131),
.B(n_1153),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1131),
.A2(n_1153),
.B(n_1155),
.C(n_867),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_867),
.B2(n_1147),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1134),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1091),
.A2(n_1148),
.B(n_1133),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1091),
.A2(n_1148),
.B(n_1133),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1076),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1100),
.B(n_1026),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1124),
.B(n_1130),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1091),
.A2(n_1148),
.B(n_1133),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1147),
.B(n_992),
.C(n_1131),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1109),
.A2(n_1104),
.A3(n_1105),
.B(n_1103),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1111),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1123),
.A2(n_1126),
.B(n_1047),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_867),
.B2(n_1147),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1111),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_1008),
.B2(n_1147),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1129),
.A2(n_1146),
.B(n_1153),
.C(n_1131),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_867),
.B2(n_1147),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1111),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1129),
.A2(n_1008),
.B1(n_1146),
.B2(n_1066),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1080),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1129),
.A2(n_1146),
.B(n_1153),
.C(n_1131),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1135),
.B(n_1149),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1079),
.B(n_1012),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_L g1240 ( 
.A(n_1147),
.B(n_1096),
.C(n_1131),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1135),
.B(n_1149),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1111),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1124),
.B(n_1130),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1123),
.A2(n_1126),
.B(n_1047),
.Y(n_1244)
);

AOI221xp5_ASAP7_75t_L g1245 ( 
.A1(n_1147),
.A2(n_726),
.B1(n_1138),
.B2(n_1096),
.C(n_1101),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1151),
.A2(n_1052),
.B1(n_1146),
.B2(n_1129),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1135),
.B(n_1149),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_867),
.B2(n_1147),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1118),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1129),
.A2(n_1146),
.B1(n_1008),
.B2(n_1147),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_SL g1251 ( 
.A(n_1096),
.B(n_867),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1111),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1111),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1147),
.B(n_992),
.C(n_1131),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1070),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1254),
.C(n_1240),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1179),
.A2(n_1218),
.B1(n_1183),
.B2(n_1246),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1179),
.B(n_1169),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1167),
.B(n_1213),
.Y(n_1259)
);

AOI221x1_ASAP7_75t_SL g1260 ( 
.A1(n_1217),
.A2(n_1229),
.B1(n_1233),
.B2(n_1248),
.C(n_1212),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1214),
.B(n_1227),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1230),
.B(n_1234),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1193),
.A2(n_1166),
.B(n_1211),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1196),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1173),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1159),
.A2(n_1245),
.B(n_1251),
.C(n_1240),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1242),
.B(n_1252),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1215),
.A2(n_1160),
.B(n_1216),
.C(n_1237),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1243),
.B(n_1200),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1215),
.A2(n_1160),
.B(n_1216),
.C(n_1237),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1245),
.A2(n_1168),
.B(n_1232),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1253),
.B(n_1205),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1185),
.B(n_1212),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1183),
.B(n_1218),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1188),
.B(n_1174),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1255),
.B(n_1221),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1161),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1232),
.A2(n_1157),
.B(n_1246),
.C(n_1180),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1190),
.B(n_1204),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1157),
.A2(n_1186),
.B(n_1198),
.C(n_1203),
.Y(n_1280)
);

CKINVDCx8_ASAP7_75t_R g1281 ( 
.A(n_1236),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1231),
.B(n_1250),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1161),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1231),
.B(n_1250),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1207),
.A2(n_1199),
.B(n_1184),
.C(n_1189),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1158),
.A2(n_1247),
.B1(n_1241),
.B2(n_1238),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1196),
.Y(n_1287)
);

AOI221x1_ASAP7_75t_SL g1288 ( 
.A1(n_1191),
.A2(n_1210),
.B1(n_1178),
.B2(n_1235),
.C(n_1221),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1201),
.B(n_1181),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1197),
.Y(n_1290)
);

AOI221x1_ASAP7_75t_SL g1291 ( 
.A1(n_1194),
.A2(n_1187),
.B1(n_1172),
.B2(n_1209),
.C(n_1206),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1162),
.A2(n_1228),
.B1(n_1244),
.B2(n_1165),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1219),
.A2(n_1224),
.B(n_1220),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1194),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1244),
.A2(n_1165),
.B1(n_1170),
.B2(n_1172),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1175),
.A2(n_1192),
.B1(n_1171),
.B2(n_1222),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1175),
.A2(n_1192),
.B1(n_1171),
.B2(n_1222),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1208),
.A2(n_1195),
.B(n_1239),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1177),
.B(n_1226),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1163),
.B(n_1202),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1177),
.B(n_1226),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1249),
.B(n_1179),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1161),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1161),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1182),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1193),
.A2(n_1166),
.B(n_1211),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1193),
.A2(n_1166),
.B(n_1211),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1221),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1245),
.A2(n_1179),
.B1(n_1146),
.B2(n_1129),
.Y(n_1309)
);

INVx8_ASAP7_75t_L g1310 ( 
.A(n_1161),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1176),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1164),
.B(n_1223),
.Y(n_1312)
);

INVx3_ASAP7_75t_SL g1313 ( 
.A(n_1236),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1179),
.B(n_1169),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1254),
.C(n_1240),
.Y(n_1315)
);

OAI211xp5_ASAP7_75t_L g1316 ( 
.A1(n_1159),
.A2(n_1179),
.B(n_1251),
.C(n_1245),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1179),
.B(n_1169),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1251),
.A2(n_1153),
.B(n_1131),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1164),
.B(n_1223),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1193),
.A2(n_1166),
.B(n_1211),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1245),
.A2(n_1179),
.B1(n_1146),
.B2(n_1129),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1164),
.B(n_1223),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1193),
.A2(n_1166),
.B(n_1211),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1179),
.B(n_1169),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1254),
.C(n_1240),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1221),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1161),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1159),
.A2(n_1225),
.B(n_1254),
.C(n_1240),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1298),
.B(n_1271),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1308),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1326),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1263),
.B(n_1306),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1263),
.B(n_1306),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1307),
.B(n_1320),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1265),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1290),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1309),
.A2(n_1321),
.B1(n_1284),
.B2(n_1282),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1307),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1299),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1301),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1323),
.B(n_1292),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1323),
.B(n_1292),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1293),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1302),
.B(n_1279),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1302),
.B(n_1275),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1276),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1309),
.A2(n_1273),
.B(n_1278),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1293),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1273),
.A2(n_1280),
.B(n_1318),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1282),
.A2(n_1284),
.B(n_1285),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1311),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1272),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1266),
.A2(n_1295),
.B(n_1267),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1296),
.B(n_1297),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1259),
.A2(n_1267),
.B(n_1262),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1272),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1259),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1316),
.B(n_1324),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1261),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1296),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1261),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1258),
.Y(n_1362)
);

AOI33xp33_ASAP7_75t_L g1363 ( 
.A1(n_1256),
.A2(n_1328),
.A3(n_1315),
.B1(n_1325),
.B2(n_1270),
.B3(n_1268),
.Y(n_1363)
);

NOR4xp25_ASAP7_75t_SL g1364 ( 
.A(n_1360),
.B(n_1327),
.C(n_1277),
.D(n_1283),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1329),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1362),
.B(n_1359),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1362),
.B(n_1314),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1335),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1330),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1358),
.A2(n_1317),
.B1(n_1258),
.B2(n_1324),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_1349),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1344),
.B(n_1314),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1341),
.B(n_1312),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1330),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1359),
.B(n_1317),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1358),
.B(n_1305),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1341),
.B(n_1322),
.Y(n_1377)
);

INVx4_ASAP7_75t_SL g1378 ( 
.A(n_1329),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1341),
.B(n_1300),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1342),
.B(n_1319),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1331),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1342),
.B(n_1269),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1343),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1331),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1332),
.B(n_1333),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1336),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1355),
.B(n_1286),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1348),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1370),
.B(n_1349),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1368),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1371),
.A2(n_1347),
.B1(n_1349),
.B2(n_1350),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1373),
.B(n_1346),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1371),
.A2(n_1347),
.B1(n_1349),
.B2(n_1350),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1378),
.B(n_1360),
.Y(n_1395)
);

OAI33xp33_ASAP7_75t_L g1396 ( 
.A1(n_1370),
.A2(n_1257),
.A3(n_1352),
.B1(n_1356),
.B2(n_1345),
.B3(n_1357),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_R g1397 ( 
.A(n_1364),
.B(n_1303),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1368),
.Y(n_1398)
);

OAI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1371),
.A2(n_1288),
.B1(n_1260),
.B2(n_1291),
.C(n_1388),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1372),
.B(n_1346),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1387),
.Y(n_1401)
);

AOI33xp33_ASAP7_75t_L g1402 ( 
.A1(n_1386),
.A2(n_1337),
.A3(n_1363),
.B1(n_1333),
.B2(n_1332),
.B3(n_1334),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1375),
.B(n_1357),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1371),
.A2(n_1337),
.B1(n_1329),
.B2(n_1354),
.C(n_1356),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1373),
.B(n_1351),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1384),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1375),
.B(n_1361),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1366),
.B(n_1374),
.C(n_1369),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_L g1409 ( 
.A(n_1369),
.B(n_1381),
.C(n_1374),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1364),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1367),
.B(n_1361),
.Y(n_1411)
);

NAND2x1_ASAP7_75t_L g1412 ( 
.A(n_1379),
.B(n_1354),
.Y(n_1412)
);

AOI211xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1376),
.A2(n_1334),
.B(n_1333),
.C(n_1338),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1381),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1385),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1385),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1383),
.B(n_1340),
.C(n_1339),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1414),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1415),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1398),
.Y(n_1420)
);

CKINVDCx14_ASAP7_75t_R g1421 ( 
.A(n_1405),
.Y(n_1421)
);

INVxp33_ASAP7_75t_SL g1422 ( 
.A(n_1410),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1415),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1402),
.B(n_1365),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1413),
.B(n_1386),
.Y(n_1425)
);

INVx4_ASAP7_75t_SL g1426 ( 
.A(n_1395),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1391),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1412),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1390),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1417),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1392),
.A2(n_1389),
.B(n_1383),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1410),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1393),
.B(n_1386),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1416),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1400),
.B(n_1382),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1399),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1402),
.B(n_1382),
.Y(n_1437)
);

AOI21xp33_ASAP7_75t_L g1438 ( 
.A1(n_1394),
.A2(n_1347),
.B(n_1350),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1408),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1401),
.Y(n_1440)
);

NOR2x1p5_ASAP7_75t_L g1441 ( 
.A(n_1412),
.B(n_1294),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1409),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1426),
.B(n_1393),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1427),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1439),
.B(n_1403),
.Y(n_1445)
);

NAND5xp2_ASAP7_75t_L g1446 ( 
.A(n_1436),
.B(n_1274),
.C(n_1397),
.D(n_1404),
.E(n_1405),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1431),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1426),
.B(n_1373),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1432),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1426),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1426),
.B(n_1377),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1426),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1431),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1426),
.B(n_1377),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1425),
.B(n_1421),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1437),
.B(n_1400),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1439),
.B(n_1407),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1437),
.B(n_1411),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1436),
.A2(n_1347),
.B(n_1350),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1431),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1433),
.B(n_1377),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1431),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1433),
.B(n_1380),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1422),
.B(n_1304),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1428),
.B(n_1424),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1431),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1442),
.Y(n_1467)
);

AND2x4_ASAP7_75t_SL g1468 ( 
.A(n_1428),
.B(n_1395),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1442),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1420),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1441),
.B(n_1406),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1430),
.B(n_1428),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1420),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1467),
.A2(n_1396),
.B1(n_1353),
.B2(n_1438),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1467),
.B(n_1430),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1455),
.B(n_1434),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1434),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1450),
.B(n_1418),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1470),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1428),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1470),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1449),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1452),
.B(n_1418),
.Y(n_1483)
);

NAND4xp25_ASAP7_75t_L g1484 ( 
.A(n_1469),
.B(n_1419),
.C(n_1423),
.D(n_1440),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1466),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1469),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1449),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1473),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1464),
.Y(n_1489)
);

AND2x4_ASAP7_75t_SL g1490 ( 
.A(n_1443),
.B(n_1471),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1452),
.B(n_1310),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1468),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1448),
.B(n_1440),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1459),
.A2(n_1353),
.B1(n_1438),
.B2(n_1466),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1466),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1448),
.B(n_1419),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1445),
.B(n_1457),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1473),
.Y(n_1498)
);

NOR2xp67_ASAP7_75t_R g1499 ( 
.A(n_1466),
.B(n_1432),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1451),
.B(n_1423),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_L g1501 ( 
.A(n_1472),
.B(n_1310),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1444),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1472),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1472),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1444),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1447),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1445),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1456),
.B(n_1435),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1456),
.B(n_1429),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1502),
.B(n_1468),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1479),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1476),
.B(n_1451),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1476),
.B(n_1454),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1481),
.Y(n_1517)
);

CKINVDCx16_ASAP7_75t_R g1518 ( 
.A(n_1489),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1481),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1488),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_SL g1521 ( 
.A(n_1475),
.B(n_1310),
.Y(n_1521)
);

NOR2x1_ASAP7_75t_L g1522 ( 
.A(n_1475),
.B(n_1446),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1474),
.A2(n_1446),
.B1(n_1459),
.B2(n_1453),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_SL g1524 ( 
.A(n_1489),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1502),
.B(n_1443),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1489),
.Y(n_1526)
);

AND3x1_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1477),
.C(n_1502),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1477),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1458),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1488),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1454),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1461),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1507),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1474),
.A2(n_1447),
.B1(n_1453),
.B2(n_1460),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1493),
.B(n_1461),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1463),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1522),
.A2(n_1494),
.B1(n_1510),
.B2(n_1462),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_SL g1538 ( 
.A1(n_1522),
.A2(n_1492),
.B(n_1499),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1524),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1511),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1526),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1511),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_L g1543 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1543)
);

OAI211xp5_ASAP7_75t_L g1544 ( 
.A1(n_1526),
.A2(n_1484),
.B(n_1487),
.C(n_1482),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1523),
.A2(n_1494),
.B1(n_1432),
.B2(n_1447),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1513),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1534),
.A2(n_1453),
.B1(n_1462),
.B2(n_1460),
.Y(n_1547)
);

O2A1O1Ixp5_ASAP7_75t_L g1548 ( 
.A1(n_1516),
.A2(n_1495),
.B(n_1485),
.C(n_1507),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1513),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_L g1550 ( 
.A1(n_1514),
.A2(n_1484),
.B(n_1496),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1521),
.A2(n_1510),
.B1(n_1462),
.B2(n_1460),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1518),
.B(n_1504),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1518),
.B(n_1496),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1517),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1514),
.B(n_1500),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1539),
.B(n_1526),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1556),
.B(n_1508),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1552),
.B(n_1529),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1553),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1539),
.B(n_1515),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1541),
.B(n_1515),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1543),
.B(n_1512),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1550),
.B(n_1512),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1544),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1545),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1544),
.B(n_1535),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1561),
.B(n_1535),
.Y(n_1569)
);

NOR3xp33_ASAP7_75t_L g1570 ( 
.A(n_1565),
.B(n_1537),
.C(n_1548),
.Y(n_1570)
);

NAND4xp25_ASAP7_75t_L g1571 ( 
.A(n_1557),
.B(n_1548),
.C(n_1521),
.D(n_1512),
.Y(n_1571)
);

OAI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1565),
.A2(n_1547),
.B1(n_1527),
.B2(n_1533),
.C(n_1505),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1566),
.A2(n_1551),
.B1(n_1527),
.B2(n_1538),
.C(n_1533),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1563),
.A2(n_1512),
.B(n_1525),
.Y(n_1574)
);

OAI21xp33_ASAP7_75t_L g1575 ( 
.A1(n_1564),
.A2(n_1532),
.B(n_1525),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1563),
.B(n_1281),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1568),
.A2(n_1529),
.B1(n_1499),
.B2(n_1554),
.C(n_1555),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1559),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_L g1579 ( 
.A(n_1578),
.B(n_1557),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1570),
.A2(n_1533),
.B1(n_1485),
.B2(n_1495),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1572),
.A2(n_1560),
.B1(n_1562),
.B2(n_1558),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1569),
.Y(n_1582)
);

AOI32xp33_ASAP7_75t_L g1583 ( 
.A1(n_1573),
.A2(n_1560),
.A3(n_1567),
.B1(n_1549),
.B2(n_1546),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1579),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1581),
.B(n_1582),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1580),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1583),
.B(n_1575),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1579),
.Y(n_1588)
);

XNOR2xp5_ASAP7_75t_L g1589 ( 
.A(n_1579),
.B(n_1571),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1584),
.A2(n_1577),
.B1(n_1574),
.B2(n_1525),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1586),
.A2(n_1542),
.B1(n_1519),
.B2(n_1520),
.C(n_1530),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1588),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1589),
.Y(n_1593)
);

AOI321xp33_ASAP7_75t_L g1594 ( 
.A1(n_1585),
.A2(n_1519),
.A3(n_1520),
.B1(n_1530),
.B2(n_1525),
.C(n_1465),
.Y(n_1594)
);

NAND4xp75_ASAP7_75t_L g1595 ( 
.A(n_1592),
.B(n_1587),
.C(n_1531),
.D(n_1483),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1593),
.B(n_1576),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1590),
.B(n_1483),
.C(n_1478),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1595),
.Y(n_1598)
);

OAI322xp33_ASAP7_75t_L g1599 ( 
.A1(n_1598),
.A2(n_1596),
.A3(n_1597),
.B1(n_1594),
.B2(n_1591),
.C1(n_1503),
.C2(n_1506),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1599),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1599),
.A2(n_1503),
.B1(n_1506),
.B2(n_1480),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1600),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1601),
.A2(n_1498),
.B(n_1531),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1602),
.A2(n_1480),
.B(n_1478),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1604),
.Y(n_1605)
);

AOI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1605),
.A2(n_1603),
.B(n_1498),
.Y(n_1606)
);

AOI222xp33_ASAP7_75t_L g1607 ( 
.A1(n_1606),
.A2(n_1532),
.B1(n_1480),
.B2(n_1536),
.C1(n_1313),
.C2(n_1501),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1607),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1608),
.A2(n_1480),
.B1(n_1536),
.B2(n_1509),
.Y(n_1609)
);

AOI211xp5_ASAP7_75t_L g1610 ( 
.A1(n_1609),
.A2(n_1264),
.B(n_1287),
.C(n_1289),
.Y(n_1610)
);


endmodule