module fake_jpeg_10778_n_470 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_470);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_470;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_48),
.B(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

CKINVDCx11_ASAP7_75t_R g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_72),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_14),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_78),
.B(n_80),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_11),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_11),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_1),
.Y(n_112)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_86),
.B(n_87),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_22),
.B(n_1),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_90),
.Y(n_116)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_92),
.Y(n_123)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_22),
.B1(n_43),
.B2(n_38),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_99),
.A2(n_27),
.B1(n_3),
.B2(n_5),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_114),
.Y(n_167)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_31),
.B(n_38),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_111),
.A2(n_8),
.B(n_10),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_112),
.B(n_133),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_47),
.A2(n_20),
.B1(n_17),
.B2(n_42),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_128),
.B1(n_37),
.B2(n_30),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_54),
.B1(n_88),
.B2(n_85),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_118),
.A2(n_27),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_64),
.A2(n_20),
.B1(n_43),
.B2(n_38),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_37),
.B1(n_30),
.B2(n_45),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_31),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_130),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_72),
.B1(n_20),
.B2(n_42),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g129 ( 
.A(n_57),
.B(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_31),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_55),
.B(n_43),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_17),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_104),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_56),
.B(n_42),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_140),
.B(n_3),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_52),
.A2(n_45),
.B(n_44),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_35),
.Y(n_166)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_150),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_29),
.B1(n_45),
.B2(n_44),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_151),
.A2(n_155),
.B1(n_161),
.B2(n_165),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_74),
.B1(n_71),
.B2(n_91),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_152),
.A2(n_154),
.B1(n_158),
.B2(n_183),
.Y(n_230)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_164),
.Y(n_214)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_157),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_51),
.B1(n_49),
.B2(n_44),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_162),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_129),
.B(n_109),
.C(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_163),
.B(n_173),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_166),
.A2(n_202),
.B(n_10),
.Y(n_218)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_34),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_93),
.B(n_29),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_174),
.B(n_175),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_29),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_121),
.C(n_124),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_180),
.C(n_181),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_111),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_177),
.A2(n_190),
.B1(n_155),
.B2(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_1),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_104),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_116),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_126),
.A2(n_135),
.B1(n_136),
.B2(n_103),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_192),
.B1(n_201),
.B2(n_146),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_125),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_2),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_141),
.B1(n_101),
.B2(n_144),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_2),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_8),
.Y(n_215)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_27),
.B1(n_5),
.B2(n_6),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_27),
.B(n_7),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_96),
.B(n_95),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_123),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_203),
.Y(n_228)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_97),
.Y(n_198)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_101),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_136),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_98),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_143),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_206),
.A2(n_210),
.B(n_225),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_167),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_213),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_95),
.B(n_96),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_211),
.B(n_215),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_150),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_217),
.A2(n_219),
.B1(n_235),
.B2(n_252),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_171),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_172),
.A2(n_106),
.B1(n_139),
.B2(n_144),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_106),
.B(n_102),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_221),
.A2(n_232),
.B(n_222),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_182),
.A2(n_102),
.B(n_143),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_240),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_230),
.B1(n_213),
.B2(n_239),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_146),
.B1(n_160),
.B2(n_156),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_169),
.B1(n_152),
.B2(n_160),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_236),
.A2(n_239),
.B1(n_237),
.B2(n_249),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_169),
.A2(n_188),
.B1(n_186),
.B2(n_185),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_161),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_248),
.C(n_211),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_202),
.A2(n_195),
.B(n_165),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_243),
.A2(n_247),
.B(n_250),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_229),
.B1(n_240),
.B2(n_221),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_177),
.A2(n_163),
.B(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_176),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_159),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_164),
.A2(n_170),
.B(n_189),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_253),
.B(n_295),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_260),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_212),
.A2(n_193),
.B1(n_197),
.B2(n_168),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_205),
.B(n_203),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_259),
.B(n_265),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_209),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_278),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_190),
.B1(n_157),
.B2(n_153),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_263),
.A2(n_271),
.B1(n_273),
.B2(n_292),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_264),
.B(n_266),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g265 ( 
.A(n_205),
.B(n_198),
.C(n_204),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_194),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_267),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_191),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_285),
.B1(n_290),
.B2(n_245),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_230),
.A2(n_233),
.B1(n_207),
.B2(n_206),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_215),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_277),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_228),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_280),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_228),
.B(n_227),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_218),
.B(n_225),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_284),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_289),
.Y(n_300)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_229),
.B(n_220),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_210),
.B(n_224),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_288),
.B(n_294),
.C(n_251),
.D(n_223),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_238),
.B(n_249),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_244),
.A2(n_237),
.B1(n_224),
.B2(n_226),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_216),
.B(n_231),
.C(n_246),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_298),
.A2(n_310),
.B1(n_288),
.B2(n_271),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_301),
.B(n_305),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_245),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_307),
.A2(n_266),
.B(n_257),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_223),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_312),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_241),
.B1(n_284),
.B2(n_255),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_256),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_323),
.Y(n_337)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_256),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_241),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_295),
.C(n_266),
.Y(n_358)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_327),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_241),
.B1(n_292),
.B2(n_263),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_290),
.B1(n_255),
.B2(n_258),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_254),
.B(n_260),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_331),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_275),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_332),
.B(n_276),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_268),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_333),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_310),
.B1(n_314),
.B2(n_318),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_287),
.B(n_279),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_343),
.B(n_344),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_323),
.Y(n_338)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_281),
.B(n_258),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_271),
.Y(n_346)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_264),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_357),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_348),
.B(n_363),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_296),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_359),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_298),
.A2(n_271),
.B1(n_287),
.B2(n_286),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_362),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_352),
.A2(n_317),
.B(n_304),
.Y(n_374)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_271),
.Y(n_355)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_303),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_361),
.Y(n_368)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_318),
.A2(n_267),
.B(n_276),
.Y(n_360)
);

XOR2x2_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_325),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_270),
.C(n_274),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_300),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_303),
.C(n_314),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_365),
.A2(n_385),
.B1(n_389),
.B2(n_364),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_381),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_297),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_372),
.B(n_377),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_386),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_313),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_336),
.A2(n_307),
.B(n_317),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_380),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_351),
.A2(n_328),
.B(n_329),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_352),
.A2(n_328),
.B(n_308),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_364),
.B(n_306),
.Y(n_383)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_319),
.Y(n_384)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_343),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_343),
.A2(n_311),
.B(n_321),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_311),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_387),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_337),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_360),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_373),
.A2(n_334),
.B1(n_346),
.B2(n_355),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_393),
.A2(n_387),
.B1(n_384),
.B2(n_375),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_361),
.C(n_357),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_397),
.C(n_400),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_383),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_398),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_358),
.C(n_363),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_348),
.C(n_337),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_340),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_402),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_344),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_390),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_367),
.A2(n_342),
.B1(n_362),
.B2(n_345),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_405),
.A2(n_411),
.B1(n_379),
.B2(n_370),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_339),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_407),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_365),
.B(n_341),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_369),
.B1(n_380),
.B2(n_389),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_390),
.B1(n_371),
.B2(n_373),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_371),
.A2(n_341),
.B1(n_354),
.B2(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_409),
.B(n_370),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_414),
.B(n_415),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_385),
.C(n_374),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_422),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_417),
.A2(n_410),
.B1(n_399),
.B2(n_382),
.Y(n_438)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_366),
.C(n_381),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_420),
.B(n_421),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_366),
.C(n_378),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_405),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_424),
.B(n_426),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_386),
.C(n_379),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_335),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_382),
.C(n_375),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_407),
.C(n_398),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_404),
.B(n_391),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_430),
.A2(n_431),
.B(n_425),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_SL g431 ( 
.A(n_415),
.B(n_406),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_437),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_391),
.C(n_393),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_423),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_335),
.C(n_349),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_425),
.C(n_423),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_441),
.A2(n_418),
.B1(n_428),
.B2(n_359),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_426),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_446),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_435),
.B(n_420),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_439),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_444),
.A2(n_450),
.B1(n_438),
.B2(n_448),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_430),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_421),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_448),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_345),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_356),
.B(n_316),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_451),
.B(n_429),
.Y(n_458)
);

NOR2x1p5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_456),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_455),
.B(n_446),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_433),
.C(n_432),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_433),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_458),
.A2(n_315),
.B1(n_326),
.B2(n_443),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_460),
.B(n_457),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_461),
.B(n_462),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_459),
.A2(n_453),
.B(n_454),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_315),
.Y(n_467)
);

NOR3xp33_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_455),
.C(n_456),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_L g468 ( 
.A1(n_466),
.A2(n_467),
.B(n_463),
.Y(n_468)
);

AOI21xp33_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_316),
.B(n_299),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_299),
.Y(n_470)
);


endmodule