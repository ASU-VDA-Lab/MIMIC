module fake_jpeg_7041_n_291 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_291);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_20),
.Y(n_49)
);

NAND2xp67_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_29),
.B(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_17),
.B1(n_13),
.B2(n_35),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_73),
.B1(n_53),
.B2(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_47),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_69),
.B1(n_15),
.B2(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22x1_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_35),
.B1(n_34),
.B2(n_31),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_73),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_45),
.B1(n_42),
.B2(n_53),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_45),
.B1(n_53),
.B2(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_39),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_28),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_97),
.C(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_43),
.B1(n_15),
.B2(n_55),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_43),
.B1(n_23),
.B2(n_21),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_76),
.B1(n_24),
.B2(n_22),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_28),
.C(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_101),
.B(n_104),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_90),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_108),
.B1(n_101),
.B2(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_75),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_70),
.C(n_74),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_91),
.C(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_76),
.B1(n_75),
.B2(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_76),
.B1(n_62),
.B2(n_61),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_112),
.B1(n_121),
.B2(n_95),
.Y(n_143)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_114),
.B(n_22),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_67),
.B1(n_66),
.B2(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_23),
.B(n_21),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_119),
.Y(n_123)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_91),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_57),
.B1(n_34),
.B2(n_31),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_21),
.B(n_89),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_131),
.B(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_83),
.B1(n_51),
.B2(n_41),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_107),
.C(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_28),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_18),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_142),
.B(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_90),
.B(n_60),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_85),
.B1(n_83),
.B2(n_51),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_108),
.B1(n_103),
.B2(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_164),
.C(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_121),
.B1(n_119),
.B2(n_116),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_110),
.B1(n_85),
.B2(n_100),
.Y(n_153)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_26),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_144),
.B(n_123),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_141),
.B1(n_130),
.B2(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_100),
.B1(n_41),
.B2(n_26),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_26),
.B1(n_18),
.B2(n_16),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_41),
.B1(n_26),
.B2(n_18),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_18),
.B1(n_16),
.B2(n_2),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_170),
.B1(n_140),
.B2(n_124),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_132),
.B1(n_135),
.B2(n_125),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_168),
.B(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_177),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_137),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_180),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_135),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_183),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_135),
.C(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_126),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_138),
.C(n_124),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_194),
.B(n_165),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_147),
.B1(n_146),
.B2(n_167),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_200),
.B1(n_184),
.B2(n_188),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_152),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_168),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_147),
.B1(n_166),
.B2(n_148),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_192),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_211),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_158),
.B1(n_150),
.B2(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_176),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_163),
.B1(n_136),
.B2(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_136),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_225),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_0),
.B(n_3),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_183),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_176),
.B(n_186),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_227),
.B(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_189),
.C(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_175),
.C(n_172),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_231),
.C(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_175),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_SL g232 ( 
.A(n_198),
.B(n_0),
.C(n_1),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_3),
.B(n_4),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_211),
.B1(n_199),
.B2(n_209),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_213),
.B1(n_195),
.B2(n_16),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_238),
.A2(n_242),
.B1(n_244),
.B2(n_232),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_195),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_229),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_227),
.B1(n_231),
.B2(n_224),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_5),
.B(n_6),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_3),
.C(n_4),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_221),
.C(n_6),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_224),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.C(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_6),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_258),
.B(n_259),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_8),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_268),
.B(n_271),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_262),
.B(n_267),
.Y(n_279)
);

FAx1_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_236),
.CI(n_239),
.CON(n_264),
.SN(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_234),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_9),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_244),
.C(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_8),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_274),
.B(n_278),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_249),
.B(n_257),
.C(n_12),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_275),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_11),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_11),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_281),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_264),
.C(n_11),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_280),
.C(n_284),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_283),
.C(n_279),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_288),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_286),
.B(n_274),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_12),
.B(n_277),
.Y(n_291)
);


endmodule