module fake_jpeg_728_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_42),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_62),
.Y(n_79)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_2),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_12),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_17),
.B(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_64),
.B1(n_36),
.B2(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_82),
.B1(n_26),
.B2(n_22),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_92),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_36),
.B1(n_24),
.B2(n_30),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_73),
.B1(n_89),
.B2(n_60),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_31),
.C(n_38),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_99),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_39),
.B1(n_27),
.B2(n_30),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_32),
.B1(n_33),
.B2(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_33),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_38),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_37),
.B1(n_31),
.B2(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_50),
.B(n_17),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_32),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_57),
.B1(n_86),
.B2(n_99),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_17),
.C(n_26),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_35),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_26),
.B1(n_22),
.B2(n_7),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_29),
.B(n_26),
.C(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_26),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_48),
.B1(n_49),
.B2(n_47),
.Y(n_116)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_35),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_87),
.B(n_77),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_68),
.C(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_2),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_80),
.B1(n_102),
.B2(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_78),
.B1(n_75),
.B2(n_88),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_153),
.B1(n_159),
.B2(n_161),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_128),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_124),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_78),
.B1(n_75),
.B2(n_88),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_127),
.B1(n_129),
.B2(n_118),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_102),
.B1(n_98),
.B2(n_83),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_80),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_130),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_110),
.Y(n_165)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_128),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_157),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_172),
.Y(n_199)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NOR4xp25_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_128),
.C(n_119),
.D(n_129),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_184),
.A3(n_148),
.B1(n_153),
.B2(n_150),
.C1(n_116),
.C2(n_22),
.Y(n_200)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_115),
.B1(n_114),
.B2(n_111),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_178),
.B1(n_158),
.B2(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_106),
.B1(n_120),
.B2(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_182),
.B(n_139),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_123),
.C(n_132),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_186),
.C(n_126),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_159),
.B(n_135),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_131),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_139),
.B1(n_147),
.B2(n_151),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_192),
.B1(n_203),
.B2(n_204),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_198),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_170),
.B1(n_164),
.B2(n_151),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_138),
.B(n_162),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_197),
.B(n_188),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_140),
.B(n_163),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_171),
.C(n_8),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_150),
.B1(n_116),
.B2(n_121),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_155),
.B1(n_4),
.B2(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_208),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_198),
.C(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_213),
.C(n_3),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_181),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_190),
.A3(n_197),
.B1(n_199),
.B2(n_174),
.C1(n_172),
.C2(n_201),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_179),
.C(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_155),
.Y(n_215)
);

NAND4xp25_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_195),
.C(n_199),
.D(n_204),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_187),
.B(n_178),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_199),
.B1(n_203),
.B2(n_191),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_221),
.B1(n_210),
.B2(n_214),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_202),
.B1(n_201),
.B2(n_185),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_214),
.C(n_8),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_217),
.B1(n_212),
.B2(n_216),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_212),
.B(n_207),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_233),
.B(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_225),
.B1(n_222),
.B2(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_235),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_227),
.B(n_226),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_10),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_3),
.B(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_230),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_241),
.B(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_232),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_226),
.B(n_10),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_244),
.B1(n_235),
.B2(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_234),
.C(n_228),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_239),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_248),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_249),
.Y(n_252)
);


endmodule