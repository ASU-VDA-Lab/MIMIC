module fake_netlist_6_1074_n_84 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_84);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_84;

wire n_52;
wire n_46;
wire n_21;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_78;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

AND2x4_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_9),
.B(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_6),
.A2(n_7),
.B1(n_13),
.B2(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_1),
.B(n_4),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_25),
.Y(n_42)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_34),
.B(n_33),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_23),
.B(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_22),
.B(n_24),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_54),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_59),
.Y(n_69)
);

OAI31xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_32),
.A3(n_59),
.B(n_27),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_65),
.B(n_68),
.Y(n_71)
);

AOI321xp33_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_8),
.A3(n_35),
.B1(n_31),
.B2(n_20),
.C(n_21),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_21),
.B(n_29),
.Y(n_73)
);

AOI211xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_31),
.B(n_29),
.C(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_21),
.C(n_29),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_21),
.C(n_29),
.Y(n_77)
);

AOI211xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_29),
.B(n_37),
.C(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_75),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_71),
.B1(n_80),
.B2(n_77),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_75),
.B(n_74),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_37),
.B(n_82),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_37),
.B(n_39),
.Y(n_84)
);


endmodule