module real_aes_10662_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_1584;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_0), .A2(n_34), .B1(n_636), .B2(n_688), .C(n_689), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_0), .A2(n_275), .B1(n_361), .B2(n_642), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_1), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_2), .A2(n_69), .B1(n_482), .B2(n_894), .Y(n_1075) );
INVx1_ASAP7_75t_L g1104 ( .A(n_2), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_3), .A2(n_270), .B1(n_939), .B2(n_1158), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_3), .A2(n_270), .B1(n_950), .B2(n_1165), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_4), .A2(n_6), .B1(n_1249), .B2(n_1262), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_5), .B(n_698), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_7), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_8), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_8), .B(n_213), .Y(n_380) );
AND2x2_ASAP7_75t_L g388 ( .A(n_8), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g432 ( .A(n_8), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g1129 ( .A(n_9), .Y(n_1129) );
AOI22xp5_ASAP7_75t_L g1255 ( .A1(n_10), .A2(n_246), .B1(n_1256), .B2(n_1259), .Y(n_1255) );
INVx1_ASAP7_75t_L g596 ( .A(n_11), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_11), .A2(n_386), .B1(n_413), .B2(n_614), .C(n_620), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g1495 ( .A(n_12), .Y(n_1495) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_13), .A2(n_93), .B1(n_573), .B2(n_575), .Y(n_718) );
INVx1_ASAP7_75t_L g736 ( .A(n_13), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_14), .Y(n_1205) );
CKINVDCx14_ASAP7_75t_R g1265 ( .A(n_15), .Y(n_1265) );
INVx1_ASAP7_75t_L g1573 ( .A(n_16), .Y(n_1573) );
OAI22xp5_ASAP7_75t_L g1578 ( .A1(n_16), .A2(n_77), .B1(n_534), .B2(n_535), .Y(n_1578) );
INVx1_ASAP7_75t_L g707 ( .A(n_17), .Y(n_707) );
INVx1_ASAP7_75t_L g630 ( .A(n_18), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_18), .A2(n_25), .B1(n_573), .B2(n_575), .Y(n_643) );
INVx1_ASAP7_75t_L g856 ( .A(n_19), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_19), .A2(n_210), .B1(n_898), .B2(n_899), .Y(n_897) );
XNOR2xp5_ASAP7_75t_L g902 ( .A(n_20), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g1498 ( .A(n_21), .Y(n_1498) );
INVx2_ASAP7_75t_L g323 ( .A(n_22), .Y(n_323) );
OR2x2_ASAP7_75t_L g349 ( .A(n_22), .B(n_321), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_23), .A2(n_140), .B1(n_357), .B2(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g441 ( .A(n_23), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_24), .A2(n_230), .B1(n_898), .B2(n_899), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_24), .A2(n_230), .B1(n_450), .B2(n_535), .Y(n_1109) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_25), .A2(n_132), .B1(n_634), .B2(n_635), .C(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g325 ( .A(n_26), .Y(n_325) );
BUFx2_ASAP7_75t_L g370 ( .A(n_26), .Y(n_370) );
BUFx2_ASAP7_75t_L g375 ( .A(n_26), .Y(n_375) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_26), .B(n_380), .Y(n_1502) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_27), .A2(n_205), .B1(n_875), .B2(n_933), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_27), .A2(n_205), .B1(n_999), .B2(n_1000), .Y(n_998) );
INVx1_ASAP7_75t_L g916 ( .A(n_28), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_28), .A2(n_203), .B1(n_931), .B2(n_933), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_29), .A2(n_38), .B1(n_1473), .B2(n_1474), .C(n_1475), .Y(n_1472) );
INVx1_ASAP7_75t_L g1514 ( .A(n_29), .Y(n_1514) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_30), .A2(n_107), .B1(n_472), .B2(n_920), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_30), .A2(n_107), .B1(n_625), .B2(n_688), .C(n_689), .Y(n_1200) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_31), .A2(n_60), .B1(n_295), .B2(n_864), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_31), .A2(n_177), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_32), .A2(n_54), .B1(n_311), .B2(n_328), .Y(n_608) );
INVx1_ASAP7_75t_L g639 ( .A(n_32), .Y(n_639) );
INVx1_ASAP7_75t_L g1041 ( .A(n_33), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_33), .A2(n_58), .B1(n_573), .B2(n_575), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_34), .A2(n_56), .B1(n_573), .B2(n_575), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_35), .A2(n_238), .B1(n_920), .B2(n_922), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g942 ( .A1(n_35), .A2(n_238), .B1(n_935), .B2(n_943), .Y(n_942) );
XNOR2xp5_ASAP7_75t_L g1066 ( .A(n_36), .B(n_1067), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_37), .Y(n_1191) );
INVx1_ASAP7_75t_L g1511 ( .A(n_38), .Y(n_1511) );
CKINVDCx5p33_ASAP7_75t_R g1557 ( .A(n_39), .Y(n_1557) );
AOI22xp33_ASAP7_75t_SL g1187 ( .A1(n_40), .A2(n_44), .B1(n_343), .B2(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1196 ( .A(n_40), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_41), .A2(n_276), .B1(n_875), .B2(n_876), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_41), .A2(n_276), .B1(n_891), .B2(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g1567 ( .A(n_42), .Y(n_1567) );
OAI211xp5_ASAP7_75t_SL g1585 ( .A1(n_42), .A2(n_417), .B(n_1586), .C(n_1592), .Y(n_1585) );
INVx1_ASAP7_75t_L g557 ( .A(n_43), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_43), .A2(n_78), .B1(n_573), .B2(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g1195 ( .A(n_44), .Y(n_1195) );
INVx1_ASAP7_75t_L g812 ( .A(n_45), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_45), .A2(n_153), .B1(n_878), .B2(n_881), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_46), .A2(n_239), .B1(n_827), .B2(n_910), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_46), .A2(n_239), .B1(n_851), .B2(n_955), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_47), .A2(n_73), .B1(n_625), .B2(n_635), .C(n_688), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_47), .A2(n_73), .B1(n_781), .B2(n_782), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_48), .A2(n_169), .B1(n_450), .B2(n_455), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_48), .A2(n_169), .B1(n_485), .B2(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g326 ( .A(n_49), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g1562 ( .A(n_50), .Y(n_1562) );
AOI221xp5_ASAP7_75t_L g1591 ( .A1(n_51), .A2(n_278), .B1(n_428), .B2(n_635), .C(n_688), .Y(n_1591) );
OAI22xp33_ASAP7_75t_L g1597 ( .A1(n_51), .A2(n_55), .B1(n_573), .B2(n_575), .Y(n_1597) );
INVx1_ASAP7_75t_L g600 ( .A(n_52), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g627 ( .A1(n_52), .A2(n_417), .B(n_628), .C(n_637), .Y(n_627) );
INVx1_ASAP7_75t_L g524 ( .A(n_53), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_53), .A2(n_64), .B1(n_534), .B2(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g638 ( .A(n_54), .Y(n_638) );
INVx1_ASAP7_75t_L g1587 ( .A(n_55), .Y(n_1587) );
INVx1_ASAP7_75t_L g684 ( .A(n_56), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_57), .A2(n_269), .B1(n_522), .B2(n_668), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_57), .A2(n_269), .B1(n_450), .B2(n_455), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g1044 ( .A1(n_58), .A2(n_67), .B1(n_935), .B2(n_1045), .C(n_1046), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_59), .A2(n_147), .B1(n_898), .B2(n_899), .Y(n_1026) );
INVx1_ASAP7_75t_L g1058 ( .A(n_59), .Y(n_1058) );
OAI22xp33_ASAP7_75t_L g976 ( .A1(n_60), .A2(n_237), .B1(n_977), .B2(n_979), .Y(n_976) );
INVx1_ASAP7_75t_L g824 ( .A(n_61), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_61), .A2(n_124), .B1(n_883), .B2(n_885), .Y(n_882) );
INVx1_ASAP7_75t_L g1590 ( .A(n_62), .Y(n_1590) );
OAI22xp33_ASAP7_75t_L g1596 ( .A1(n_62), .A2(n_278), .B1(n_357), .B2(n_361), .Y(n_1596) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_63), .A2(n_95), .B1(n_1249), .B2(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g523 ( .A(n_64), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_65), .A2(n_386), .B1(n_391), .B2(n_403), .C(n_413), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_65), .A2(n_277), .B1(n_482), .B2(n_483), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_66), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_67), .A2(n_211), .B1(n_361), .B2(n_642), .Y(n_1064) );
INVx1_ASAP7_75t_L g1136 ( .A(n_68), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_68), .A2(n_136), .B1(n_950), .B2(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1102 ( .A(n_69), .Y(n_1102) );
AO221x1_ASAP7_75t_L g1203 ( .A1(n_70), .A2(n_86), .B1(n_634), .B2(n_636), .C(n_843), .Y(n_1203) );
INVx1_ASAP7_75t_L g1214 ( .A(n_70), .Y(n_1214) );
AOI22xp5_ASAP7_75t_SL g1270 ( .A1(n_71), .A2(n_83), .B1(n_1243), .B2(n_1249), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_72), .A2(n_249), .B1(n_352), .B2(n_483), .Y(n_1076) );
OAI211xp5_ASAP7_75t_SL g1089 ( .A1(n_72), .A2(n_417), .B(n_1090), .C(n_1098), .Y(n_1089) );
CKINVDCx16_ASAP7_75t_R g1247 ( .A(n_74), .Y(n_1247) );
INVx1_ASAP7_75t_L g402 ( .A(n_75), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_75), .A2(n_219), .B1(n_475), .B2(n_478), .Y(n_474) );
INVx1_ASAP7_75t_L g1138 ( .A(n_76), .Y(n_1138) );
AOI22xp33_ASAP7_75t_SL g1167 ( .A1(n_76), .A2(n_216), .B1(n_922), .B2(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1570 ( .A(n_77), .Y(n_1570) );
INVx1_ASAP7_75t_L g555 ( .A(n_78), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_79), .A2(n_128), .B1(n_974), .B2(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_SL g995 ( .A1(n_79), .A2(n_128), .B1(n_933), .B2(n_939), .Y(n_995) );
INVx1_ASAP7_75t_L g1132 ( .A(n_80), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_80), .A2(n_130), .B1(n_931), .B2(n_1154), .Y(n_1153) );
XNOR2x2_ASAP7_75t_L g803 ( .A(n_81), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g971 ( .A(n_82), .Y(n_971) );
OAI222xp33_ASAP7_75t_L g983 ( .A1(n_82), .A2(n_177), .B1(n_195), .B2(n_984), .C1(n_985), .C2(n_986), .Y(n_983) );
INVx1_ASAP7_75t_L g1082 ( .A(n_84), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_84), .A2(n_189), .B1(n_843), .B2(n_1046), .C(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g605 ( .A(n_85), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_85), .A2(n_148), .B1(n_534), .B2(n_535), .Y(n_612) );
INVx1_ASAP7_75t_L g1216 ( .A(n_86), .Y(n_1216) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_87), .A2(n_103), .B1(n_428), .B2(n_753), .C(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g790 ( .A(n_87), .Y(n_790) );
OAI222xp33_ASAP7_75t_L g1120 ( .A1(n_88), .A2(n_191), .B1(n_234), .B2(n_910), .C1(n_1121), .C2(n_1124), .Y(n_1120) );
INVx1_ASAP7_75t_L g1139 ( .A(n_88), .Y(n_1139) );
AO22x2_ASAP7_75t_L g1115 ( .A1(n_89), .A2(n_1116), .B1(n_1117), .B2(n_1173), .Y(n_1115) );
INVxp67_ASAP7_75t_SL g1116 ( .A(n_89), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_90), .A2(n_113), .B1(n_1152), .B2(n_1161), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_90), .A2(n_113), .B1(n_920), .B2(n_922), .Y(n_1163) );
INVx1_ASAP7_75t_L g321 ( .A(n_91), .Y(n_321) );
INVx1_ASAP7_75t_L g467 ( .A(n_91), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_92), .A2(n_167), .B1(n_922), .B2(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g961 ( .A(n_92), .Y(n_961) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_93), .A2(n_222), .B1(n_636), .B2(n_680), .C(n_689), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_94), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_96), .A2(n_98), .B1(n_328), .B2(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1048 ( .A(n_96), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_97), .A2(n_137), .B1(n_924), .B2(n_925), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_97), .A2(n_137), .B1(n_939), .B2(n_940), .Y(n_938) );
INVx1_ASAP7_75t_L g1049 ( .A(n_98), .Y(n_1049) );
XNOR2xp5_ASAP7_75t_L g1551 ( .A(n_99), .B(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g709 ( .A(n_100), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_100), .A2(n_386), .B1(n_724), .B2(n_728), .C(n_732), .Y(n_723) );
AOI22x1_ASAP7_75t_L g1175 ( .A1(n_101), .A2(n_1176), .B1(n_1177), .B2(n_1217), .Y(n_1175) );
INVxp67_ASAP7_75t_SL g1217 ( .A(n_101), .Y(n_1217) );
INVx1_ASAP7_75t_L g1128 ( .A(n_102), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1151 ( .A1(n_102), .A2(n_234), .B1(n_943), .B2(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g793 ( .A(n_103), .Y(n_793) );
XNOR2xp5_ASAP7_75t_L g580 ( .A(n_104), .B(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_105), .A2(n_250), .B1(n_1256), .B2(n_1314), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_106), .Y(n_1072) );
CKINVDCx20_ASAP7_75t_R g1354 ( .A(n_108), .Y(n_1354) );
AOI221xp5_ASAP7_75t_L g1486 ( .A1(n_109), .A2(n_164), .B1(n_949), .B2(n_1004), .C(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1531 ( .A(n_109), .Y(n_1531) );
CKINVDCx5p33_ASAP7_75t_R g1071 ( .A(n_110), .Y(n_1071) );
INVx1_ASAP7_75t_L g763 ( .A(n_111), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_111), .A2(n_248), .B1(n_477), .B2(n_480), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_112), .A2(n_186), .B1(n_892), .B2(n_999), .Y(n_1074) );
INVx1_ASAP7_75t_L g1106 ( .A(n_112), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_114), .A2(n_231), .B1(n_750), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_114), .A2(n_231), .B1(n_477), .B2(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g906 ( .A(n_115), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_115), .A2(n_200), .B1(n_635), .B2(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1028 ( .A(n_116), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_116), .A2(n_386), .B1(n_732), .B2(n_1051), .C(n_1055), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1564 ( .A(n_117), .Y(n_1564) );
INVx1_ASAP7_75t_L g514 ( .A(n_118), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_119), .A2(n_192), .B1(n_922), .B2(n_1184), .Y(n_1183) );
OAI221xp5_ASAP7_75t_L g1202 ( .A1(n_119), .A2(n_417), .B1(n_1203), .B2(n_1204), .C(n_1208), .Y(n_1202) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_120), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_121), .A2(n_225), .B1(n_949), .B2(n_950), .Y(n_1181) );
AOI22xp33_ASAP7_75t_SL g1198 ( .A1(n_121), .A2(n_225), .B1(n_399), .B2(n_1199), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g1471 ( .A(n_122), .Y(n_1471) );
INVx1_ASAP7_75t_L g1566 ( .A(n_123), .Y(n_1566) );
OAI221xp5_ASAP7_75t_L g1579 ( .A1(n_123), .A2(n_386), .B1(n_413), .B2(n_1580), .C(n_1584), .Y(n_1579) );
INVx1_ASAP7_75t_L g807 ( .A(n_124), .Y(n_807) );
INVx1_ASAP7_75t_L g286 ( .A(n_125), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g1479 ( .A1(n_126), .A2(n_252), .B1(n_1480), .B2(n_1483), .Y(n_1479) );
OAI221xp5_ASAP7_75t_L g1518 ( .A1(n_126), .A2(n_252), .B1(n_1519), .B2(n_1522), .C(n_1525), .Y(n_1518) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_127), .Y(n_913) );
INVx1_ASAP7_75t_L g710 ( .A(n_129), .Y(n_710) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_129), .A2(n_417), .B(n_734), .C(n_739), .Y(n_733) );
INVx1_ASAP7_75t_L g1131 ( .A(n_130), .Y(n_1131) );
INVx1_ASAP7_75t_L g766 ( .A(n_131), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_131), .A2(n_266), .B1(n_352), .B2(n_785), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_132), .A2(n_161), .B1(n_361), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_133), .A2(n_236), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g794 ( .A(n_133), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_134), .A2(n_235), .B1(n_1256), .B2(n_1259), .Y(n_1269) );
INVx1_ASAP7_75t_L g844 ( .A(n_135), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_135), .A2(n_215), .B1(n_482), .B2(n_894), .Y(n_896) );
INVx1_ASAP7_75t_L g1135 ( .A(n_136), .Y(n_1135) );
XOR2xp5_ASAP7_75t_L g306 ( .A(n_138), .B(n_307), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_138), .A2(n_141), .B1(n_1243), .B2(n_1316), .Y(n_1315) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_139), .Y(n_586) );
INVx1_ASAP7_75t_L g426 ( .A(n_140), .Y(n_426) );
CKINVDCx14_ASAP7_75t_R g1266 ( .A(n_142), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1273 ( .A1(n_143), .A2(n_173), .B1(n_1256), .B2(n_1259), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_144), .A2(n_227), .B1(n_447), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g797 ( .A(n_144), .Y(n_797) );
INVx1_ASAP7_75t_L g531 ( .A(n_145), .Y(n_531) );
INVx1_ASAP7_75t_L g355 ( .A(n_146), .Y(n_355) );
INVx1_ASAP7_75t_L g1061 ( .A(n_147), .Y(n_1061) );
INVx1_ASAP7_75t_L g603 ( .A(n_148), .Y(n_603) );
INVx1_ASAP7_75t_L g350 ( .A(n_149), .Y(n_350) );
INVx1_ASAP7_75t_L g798 ( .A(n_150), .Y(n_798) );
INVx1_ASAP7_75t_L g334 ( .A(n_151), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_152), .Y(n_817) );
INVx1_ASAP7_75t_L g821 ( .A(n_153), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_154), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_155), .A2(n_243), .B1(n_949), .B2(n_950), .Y(n_948) );
INVx1_ASAP7_75t_L g957 ( .A(n_155), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_156), .A2(n_233), .B1(n_527), .B2(n_529), .Y(n_715) );
INVx1_ASAP7_75t_L g741 ( .A(n_156), .Y(n_741) );
INVx1_ASAP7_75t_L g989 ( .A(n_157), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_157), .A2(n_162), .B1(n_898), .B2(n_899), .Y(n_1006) );
INVx1_ASAP7_75t_L g712 ( .A(n_158), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_158), .A2(n_265), .B1(n_534), .B2(n_535), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_159), .A2(n_190), .B1(n_871), .B2(n_872), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_159), .A2(n_190), .B1(n_469), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_160), .A2(n_247), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
INVx1_ASAP7_75t_L g1535 ( .A(n_160), .Y(n_1535) );
INVx1_ASAP7_75t_L g632 ( .A(n_161), .Y(n_632) );
INVx1_ASAP7_75t_L g990 ( .A(n_162), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_163), .A2(n_193), .B1(n_1477), .B2(n_1478), .Y(n_1476) );
INVx1_ASAP7_75t_L g1507 ( .A(n_163), .Y(n_1507) );
INVx1_ASAP7_75t_L g1533 ( .A(n_164), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_165), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_166), .Y(n_1462) );
INVx1_ASAP7_75t_L g953 ( .A(n_167), .Y(n_953) );
INVx1_ASAP7_75t_L g408 ( .A(n_168), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_168), .A2(n_197), .B1(n_469), .B2(n_472), .Y(n_468) );
AOI22x1_ASAP7_75t_SL g963 ( .A1(n_170), .A2(n_964), .B1(n_1007), .B2(n_1008), .Y(n_963) );
INVx1_ASAP7_75t_L g1007 ( .A(n_170), .Y(n_1007) );
AO221x2_ASAP7_75t_L g1263 ( .A1(n_170), .A2(n_261), .B1(n_1249), .B2(n_1262), .C(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1087 ( .A(n_171), .Y(n_1087) );
CKINVDCx16_ASAP7_75t_R g1250 ( .A(n_172), .Y(n_1250) );
INVx1_ASAP7_75t_L g968 ( .A(n_174), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_174), .A2(n_237), .B1(n_841), .B2(n_871), .Y(n_996) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_175), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_175), .B(n_286), .Y(n_1230) );
AND3x2_ASAP7_75t_L g1246 ( .A(n_175), .B(n_286), .C(n_1233), .Y(n_1246) );
INVx1_ASAP7_75t_L g664 ( .A(n_176), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_176), .A2(n_386), .B1(n_413), .B2(n_673), .C(n_678), .Y(n_672) );
AOI22xp5_ASAP7_75t_SL g1282 ( .A1(n_178), .A2(n_194), .B1(n_1243), .B2(n_1249), .Y(n_1282) );
CKINVDCx5p33_ASAP7_75t_R g1576 ( .A(n_179), .Y(n_1576) );
INVx1_ASAP7_75t_L g519 ( .A(n_180), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_180), .A2(n_417), .B1(n_549), .B2(n_556), .C(n_563), .Y(n_548) );
INVx2_ASAP7_75t_L g299 ( .A(n_181), .Y(n_299) );
AOI22xp5_ASAP7_75t_SL g1281 ( .A1(n_182), .A2(n_257), .B1(n_1256), .B2(n_1259), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_183), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g526 ( .A1(n_184), .A2(n_185), .B1(n_527), .B2(n_529), .Y(n_526) );
INVx1_ASAP7_75t_L g564 ( .A(n_184), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_185), .Y(n_566) );
INVx1_ASAP7_75t_L g1107 ( .A(n_186), .Y(n_1107) );
INVx1_ASAP7_75t_L g590 ( .A(n_187), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_187), .A2(n_623), .B(n_625), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_188), .A2(n_222), .B1(n_357), .B2(n_361), .Y(n_717) );
INVx1_ASAP7_75t_L g737 ( .A(n_188), .Y(n_737) );
INVx1_ASAP7_75t_L g1084 ( .A(n_189), .Y(n_1084) );
INVx1_ASAP7_75t_L g1141 ( .A(n_191), .Y(n_1141) );
INVx1_ASAP7_75t_L g1201 ( .A(n_192), .Y(n_1201) );
INVx1_ASAP7_75t_L g1516 ( .A(n_193), .Y(n_1516) );
XNOR2xp5_ASAP7_75t_L g1456 ( .A(n_194), .B(n_1457), .Y(n_1456) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_194), .A2(n_1546), .B1(n_1550), .B2(n_1598), .Y(n_1545) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_195), .Y(n_970) );
XNOR2xp5_ASAP7_75t_L g498 ( .A(n_196), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g410 ( .A(n_197), .Y(n_410) );
INVx1_ASAP7_75t_L g825 ( .A(n_198), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_198), .A2(n_228), .B1(n_849), .B2(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g610 ( .A(n_199), .Y(n_610) );
INVx1_ASAP7_75t_L g912 ( .A(n_200), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_201), .A2(n_204), .B1(n_527), .B2(n_529), .Y(n_669) );
INVx1_ASAP7_75t_L g692 ( .A(n_201), .Y(n_692) );
INVx1_ASAP7_75t_L g1233 ( .A(n_202), .Y(n_1233) );
INVx1_ASAP7_75t_L g915 ( .A(n_203), .Y(n_915) );
INVx1_ASAP7_75t_L g691 ( .A(n_204), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g1013 ( .A(n_206), .B(n_1014), .Y(n_1013) );
AO221x2_ASAP7_75t_L g1351 ( .A1(n_206), .A2(n_207), .B1(n_1316), .B2(n_1352), .C(n_1353), .Y(n_1351) );
INVx1_ASAP7_75t_L g1034 ( .A(n_208), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_209), .A2(n_253), .B1(n_688), .B2(n_841), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_209), .A2(n_253), .B1(n_482), .B2(n_483), .Y(n_1001) );
INVx1_ASAP7_75t_L g859 ( .A(n_210), .Y(n_859) );
INVx1_ASAP7_75t_L g1043 ( .A(n_211), .Y(n_1043) );
INVx1_ASAP7_75t_L g652 ( .A(n_212), .Y(n_652) );
INVx1_ASAP7_75t_L g301 ( .A(n_213), .Y(n_301) );
INVx2_ASAP7_75t_L g389 ( .A(n_213), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_214), .A2(n_241), .B1(n_488), .B2(n_891), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_214), .A2(n_241), .B1(n_450), .B2(n_455), .Y(n_1062) );
INVx1_ASAP7_75t_L g862 ( .A(n_215), .Y(n_862) );
INVx1_ASAP7_75t_L g1146 ( .A(n_216), .Y(n_1146) );
INVx1_ASAP7_75t_L g518 ( .A(n_217), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g536 ( .A1(n_217), .A2(n_386), .B1(n_413), .B2(n_537), .C(n_543), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_218), .Y(n_1024) );
INVx1_ASAP7_75t_L g397 ( .A(n_219), .Y(n_397) );
CKINVDCx14_ASAP7_75t_R g1356 ( .A(n_220), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_221), .A2(n_274), .B1(n_506), .B2(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g674 ( .A(n_221), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_223), .B(n_746), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g1560 ( .A(n_224), .Y(n_1560) );
INVx1_ASAP7_75t_L g702 ( .A(n_226), .Y(n_702) );
INVx1_ASAP7_75t_L g796 ( .A(n_227), .Y(n_796) );
INVx1_ASAP7_75t_L g831 ( .A(n_228), .Y(n_831) );
CKINVDCx16_ASAP7_75t_R g1240 ( .A(n_229), .Y(n_1240) );
INVx1_ASAP7_75t_L g1031 ( .A(n_232), .Y(n_1031) );
OAI211xp5_ASAP7_75t_SL g1036 ( .A1(n_232), .A2(n_417), .B(n_1037), .C(n_1047), .Y(n_1036) );
INVx1_ASAP7_75t_L g740 ( .A(n_233), .Y(n_740) );
INVx1_ASAP7_75t_L g788 ( .A(n_236), .Y(n_788) );
INVx1_ASAP7_75t_L g656 ( .A(n_240), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_240), .A2(n_625), .B(n_680), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_242), .Y(n_508) );
INVx1_ASAP7_75t_L g959 ( .A(n_243), .Y(n_959) );
INVx1_ASAP7_75t_L g704 ( .A(n_244), .Y(n_704) );
INVx1_ASAP7_75t_L g1234 ( .A(n_245), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_245), .B(n_1232), .Y(n_1239) );
INVx1_ASAP7_75t_L g1530 ( .A(n_247), .Y(n_1530) );
INVx1_ASAP7_75t_L g764 ( .A(n_248), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g1099 ( .A1(n_249), .A2(n_386), .B1(n_732), .B2(n_1100), .C(n_1105), .Y(n_1099) );
INVx1_ASAP7_75t_L g367 ( .A(n_251), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g1574 ( .A1(n_254), .A2(n_256), .B1(n_527), .B2(n_529), .Y(n_1574) );
INVx1_ASAP7_75t_L g1593 ( .A(n_254), .Y(n_1593) );
INVx1_ASAP7_75t_L g666 ( .A(n_255), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_255), .A2(n_417), .B(n_682), .C(n_690), .Y(n_681) );
INVx1_ASAP7_75t_L g1594 ( .A(n_256), .Y(n_1594) );
CKINVDCx5p33_ASAP7_75t_R g1465 ( .A(n_258), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_259), .Y(n_1025) );
INVx2_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
INVx1_ASAP7_75t_L g552 ( .A(n_262), .Y(n_552) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_262), .A2(n_268), .B1(n_357), .B2(n_361), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_263), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_264), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g714 ( .A(n_265), .Y(n_714) );
INVx1_ASAP7_75t_L g756 ( .A(n_266), .Y(n_756) );
INVx1_ASAP7_75t_L g507 ( .A(n_267), .Y(n_507) );
INVx1_ASAP7_75t_L g558 ( .A(n_268), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g1235 ( .A(n_271), .Y(n_1235) );
BUFx3_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
INVx1_ASAP7_75t_L g360 ( .A(n_272), .Y(n_360) );
BUFx3_ASAP7_75t_L g316 ( .A(n_273), .Y(n_316) );
INVx1_ASAP7_75t_L g346 ( .A(n_273), .Y(n_346) );
INVx1_ASAP7_75t_L g677 ( .A(n_274), .Y(n_677) );
INVx1_ASAP7_75t_L g686 ( .A(n_275), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_277), .A2(n_417), .B1(n_424), .B2(n_433), .C(n_442), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_279), .Y(n_1081) );
INVx1_ASAP7_75t_L g720 ( .A(n_280), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_302), .B(n_1218), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
AND2x4_ASAP7_75t_L g1544 ( .A(n_284), .B(n_290), .Y(n_1544) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g1549 ( .A(n_285), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_285), .B(n_287), .Y(n_1605) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_287), .B(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x6_ASAP7_75t_L g865 ( .A(n_292), .B(n_370), .Y(n_865) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g412 ( .A(n_293), .B(n_301), .Y(n_412) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g625 ( .A(n_294), .B(n_626), .Y(n_625) );
INVx8_ASAP7_75t_L g861 ( .A(n_295), .Y(n_861) );
OR2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_296), .Y(n_409) );
INVx2_ASAP7_75t_SL g545 ( .A(n_296), .Y(n_545) );
INVx1_ASAP7_75t_L g554 ( .A(n_296), .Y(n_554) );
BUFx2_ASAP7_75t_L g731 ( .A(n_296), .Y(n_731) );
OR2x6_ASAP7_75t_L g864 ( .A(n_296), .B(n_855), .Y(n_864) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_296), .B(n_1502), .Y(n_1501) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g383 ( .A(n_298), .B(n_299), .Y(n_383) );
INVx2_ASAP7_75t_L g396 ( .A(n_298), .Y(n_396) );
AND2x4_ASAP7_75t_L g400 ( .A(n_298), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
INVx1_ASAP7_75t_L g423 ( .A(n_298), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_299), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g401 ( .A(n_299), .Y(n_401) );
INVx1_ASAP7_75t_L g406 ( .A(n_299), .Y(n_406) );
INVx1_ASAP7_75t_L g445 ( .A(n_299), .Y(n_445) );
INVx1_ASAP7_75t_L g454 ( .A(n_299), .Y(n_454) );
AND2x4_ASAP7_75t_L g850 ( .A(n_300), .B(n_445), .Y(n_850) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g851 ( .A(n_301), .B(n_852), .Y(n_851) );
OR2x2_ASAP7_75t_L g986 ( .A(n_301), .B(n_852), .Y(n_986) );
XOR2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_644), .Y(n_302) );
XOR2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_579), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_494), .B1(n_495), .B2(n_578), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_306), .Y(n_578) );
NAND4xp75_ASAP7_75t_SL g307 ( .A(n_308), .B(n_366), .C(n_384), .D(n_462), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_341), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_326), .B1(n_327), .B2(n_334), .C(n_335), .Y(n_309) );
INVx1_ASAP7_75t_L g1018 ( .A(n_310), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_310), .A2(n_327), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g528 ( .A(n_311), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_312), .B(n_317), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g1482 ( .A(n_313), .Y(n_1482) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g830 ( .A(n_314), .Y(n_830) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g354 ( .A(n_315), .B(n_332), .Y(n_354) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g339 ( .A(n_316), .B(n_333), .Y(n_339) );
AND2x4_ASAP7_75t_L g359 ( .A(n_316), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x6_ASAP7_75t_L g328 ( .A(n_318), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g340 ( .A(n_318), .Y(n_340) );
OR2x2_ASAP7_75t_L g529 ( .A(n_318), .B(n_329), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_319), .B(n_324), .Y(n_318) );
AND2x2_ASAP7_75t_L g371 ( .A(n_319), .B(n_354), .Y(n_371) );
AND2x4_ASAP7_75t_L g1481 ( .A(n_319), .B(n_1482), .Y(n_1481) );
AND2x4_ASAP7_75t_L g1484 ( .A(n_319), .B(n_330), .Y(n_1484) );
BUFx2_ASAP7_75t_L g1497 ( .A(n_319), .Y(n_1497) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g493 ( .A(n_322), .B(n_467), .Y(n_493) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g466 ( .A(n_323), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g810 ( .A(n_323), .Y(n_810) );
INVx1_ASAP7_75t_L g815 ( .A(n_323), .Y(n_815) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_323), .Y(n_820) );
OR2x6_ASAP7_75t_L g887 ( .A(n_324), .B(n_430), .Y(n_887) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g348 ( .A(n_325), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g1510 ( .A(n_325), .B(n_388), .Y(n_1510) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_326), .A2(n_334), .B1(n_443), .B2(n_446), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_327), .A2(n_335), .B1(n_528), .B2(n_796), .C(n_797), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_327), .A2(n_335), .B1(n_528), .B2(n_1190), .C(n_1191), .Y(n_1189) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x6_ASAP7_75t_L g832 ( .A(n_331), .B(n_815), .Y(n_832) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g345 ( .A(n_333), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_335), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_335), .B(n_583), .C(n_608), .Y(n_582) );
NOR3xp33_ASAP7_75t_SL g653 ( .A(n_335), .B(n_654), .C(n_669), .Y(n_653) );
NOR3xp33_ASAP7_75t_SL g699 ( .A(n_335), .B(n_700), .C(n_715), .Y(n_699) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_335), .Y(n_1016) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_340), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g783 ( .A(n_338), .Y(n_783) );
AND2x4_ASAP7_75t_L g834 ( .A(n_338), .B(n_835), .Y(n_834) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_338), .Y(n_908) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_338), .Y(n_1005) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_339), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_340), .B(n_785), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_350), .B1(n_351), .B2(n_355), .C(n_356), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_342), .A2(n_351), .B1(n_793), .B2(n_794), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_342), .A2(n_351), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1215 ( .A1(n_342), .A2(n_791), .B1(n_1206), .B2(n_1216), .Y(n_1215) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_347), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g949 ( .A(n_344), .Y(n_949) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_345), .Y(n_477) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_345), .Y(n_487) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_345), .Y(n_506) );
BUFx3_ASAP7_75t_L g522 ( .A(n_345), .Y(n_522) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_345), .Y(n_577) );
AND2x6_ASAP7_75t_L g813 ( .A(n_345), .B(n_814), .Y(n_813) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_345), .Y(n_1165) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_345), .Y(n_1170) );
INVx1_ASAP7_75t_L g365 ( .A(n_346), .Y(n_365) );
AND2x2_ASAP7_75t_L g351 ( .A(n_347), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x6_ASAP7_75t_L g357 ( .A(n_348), .B(n_358), .Y(n_357) );
OR2x6_ASAP7_75t_L g361 ( .A(n_348), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g573 ( .A(n_348), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g575 ( .A(n_348), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g642 ( .A(n_348), .B(n_358), .Y(n_642) );
OR2x2_ASAP7_75t_L g1464 ( .A(n_349), .B(n_511), .Y(n_1464) );
INVx2_ASAP7_75t_L g1467 ( .A(n_349), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_349), .B(n_928), .Y(n_1470) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_350), .A2(n_434), .B1(n_437), .B2(n_441), .Y(n_433) );
AOI222xp33_ASAP7_75t_L g1213 ( .A1(n_351), .A2(n_369), .B1(n_789), .B2(n_1205), .C1(n_1209), .C2(n_1214), .Y(n_1213) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g482 ( .A(n_353), .Y(n_482) );
INVx1_ASAP7_75t_L g1473 ( .A(n_353), .Y(n_1473) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx6_ASAP7_75t_L g471 ( .A(n_354), .Y(n_471) );
BUFx2_ASAP7_75t_L g781 ( .A(n_354), .Y(n_781) );
AND2x4_ASAP7_75t_L g818 ( .A(n_354), .B(n_819), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_355), .A2(n_409), .B1(n_425), .B2(n_426), .C(n_427), .Y(n_424) );
CKINVDCx6p67_ASAP7_75t_R g789 ( .A(n_357), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_358), .A2(n_521), .B1(n_523), .B2(n_524), .Y(n_520) );
INVx2_ASAP7_75t_L g779 ( .A(n_358), .Y(n_779) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_359), .Y(n_480) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_359), .Y(n_490) );
INVx1_ASAP7_75t_L g587 ( .A(n_359), .Y(n_587) );
INVx2_ASAP7_75t_L g928 ( .A(n_359), .Y(n_928) );
INVx1_ASAP7_75t_L g364 ( .A(n_360), .Y(n_364) );
CKINVDCx6p67_ASAP7_75t_R g791 ( .A(n_361), .Y(n_791) );
BUFx3_ASAP7_75t_L g513 ( .A(n_362), .Y(n_513) );
OAI221xp5_ASAP7_75t_L g1020 ( .A1(n_362), .A2(n_1021), .B1(n_1024), .B2(n_1025), .C(n_1026), .Y(n_1020) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_362), .A2(n_1022), .B1(n_1566), .B2(n_1567), .Y(n_1565) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g592 ( .A(n_363), .Y(n_592) );
INVx1_ASAP7_75t_L g599 ( .A(n_363), .Y(n_599) );
BUFx4f_ASAP7_75t_L g658 ( .A(n_363), .Y(n_658) );
INVx1_ASAP7_75t_L g1126 ( .A(n_363), .Y(n_1126) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OR2x2_ASAP7_75t_L g511 ( .A(n_364), .B(n_365), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_368), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_368), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_368), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_368), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g746 ( .A(n_368), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_368), .B(n_1034), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_368), .B(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_368), .B(n_1576), .Y(n_1575) );
OR2x6_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
INVx2_ASAP7_75t_L g1503 ( .A(n_369), .Y(n_1503) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x4_ASAP7_75t_L g492 ( .A(n_370), .B(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g607 ( .A(n_370), .B(n_493), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx2_ASAP7_75t_L g772 ( .A(n_373), .Y(n_772) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x6_ASAP7_75t_L g464 ( .A(n_374), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g503 ( .A(n_374), .B(n_465), .Y(n_503) );
BUFx2_ASAP7_75t_L g569 ( .A(n_374), .Y(n_569) );
OR2x2_ASAP7_75t_L g776 ( .A(n_374), .B(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g869 ( .A(n_374), .B(n_412), .Y(n_869) );
AND2x4_ASAP7_75t_L g992 ( .A(n_374), .B(n_412), .Y(n_992) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g461 ( .A(n_375), .Y(n_461) );
OR2x6_ASAP7_75t_L g1528 ( .A(n_375), .B(n_625), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
AND2x2_ASAP7_75t_L g443 ( .A(n_377), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g565 ( .A(n_377), .B(n_444), .Y(n_565) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x6_ASAP7_75t_L g413 ( .A(n_378), .B(n_414), .Y(n_413) );
OR2x6_ASAP7_75t_L g447 ( .A(n_378), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g732 ( .A(n_378), .B(n_414), .Y(n_732) );
INVx1_ASAP7_75t_L g761 ( .A(n_378), .Y(n_761) );
INVx1_ASAP7_75t_L g1212 ( .A(n_378), .Y(n_1212) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g935 ( .A(n_381), .Y(n_935) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g634 ( .A(n_382), .Y(n_634) );
INVx2_ASAP7_75t_SL g680 ( .A(n_382), .Y(n_680) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_383), .Y(n_390) );
OAI31xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_416), .A3(n_449), .B(n_459), .Y(n_384) );
CKINVDCx6p67_ASAP7_75t_R g386 ( .A(n_387), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_387), .A2(n_766), .B1(n_767), .B2(n_768), .C(n_770), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g1197 ( .A1(n_387), .A2(n_1198), .B1(n_1200), .B2(n_1201), .Y(n_1197) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx2_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
AND2x2_ASAP7_75t_L g451 ( .A(n_388), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g431 ( .A(n_389), .Y(n_431) );
INVx1_ASAP7_75t_L g626 ( .A(n_389), .Y(n_626) );
INVx3_ASAP7_75t_L g624 ( .A(n_390), .Y(n_624) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_390), .Y(n_688) );
BUFx2_ASAP7_75t_L g753 ( .A(n_390), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_397), .B1(n_398), .B2(n_402), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g538 ( .A(n_393), .Y(n_538) );
INVx2_ASAP7_75t_L g683 ( .A(n_393), .Y(n_683) );
INVx2_ASAP7_75t_L g735 ( .A(n_393), .Y(n_735) );
BUFx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g1040 ( .A(n_394), .Y(n_1040) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
BUFx2_ASAP7_75t_L g617 ( .A(n_395), .Y(n_617) );
INVx1_ASAP7_75t_L g448 ( .A(n_396), .Y(n_448) );
AND2x4_ASAP7_75t_L g452 ( .A(n_396), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_SL g631 ( .A(n_399), .Y(n_631) );
INVx4_ASAP7_75t_L g685 ( .A(n_399), .Y(n_685) );
BUFx3_ASAP7_75t_L g881 ( .A(n_399), .Y(n_881) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g440 ( .A(n_400), .Y(n_440) );
INVx1_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
INVx1_ASAP7_75t_L g542 ( .A(n_400), .Y(n_542) );
AND2x4_ASAP7_75t_L g422 ( .A(n_401), .B(n_423), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_408), .B1(n_409), .B2(n_410), .C(n_411), .Y(n_403) );
INVx2_ASAP7_75t_L g551 ( .A(n_404), .Y(n_551) );
BUFx3_ASAP7_75t_L g621 ( .A(n_404), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_404), .B(n_1211), .Y(n_1210) );
OAI221xp5_ASAP7_75t_L g1584 ( .A1(n_404), .A2(n_409), .B1(n_546), .B2(n_1562), .C(n_1564), .Y(n_1584) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AND2x2_ASAP7_75t_L g415 ( .A(n_406), .B(n_407), .Y(n_415) );
INVx1_ASAP7_75t_L g852 ( .A(n_407), .Y(n_852) );
BUFx2_ASAP7_75t_L g1054 ( .A(n_409), .Y(n_1054) );
OAI221xp5_ASAP7_75t_L g1051 ( .A1(n_411), .A2(n_1024), .B1(n_1025), .B2(n_1052), .C(n_1054), .Y(n_1051) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_411), .A2(n_1101), .B1(n_1102), .B2(n_1103), .C(n_1104), .Y(n_1100) );
BUFx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g547 ( .A(n_412), .Y(n_547) );
INVx2_ASAP7_75t_L g770 ( .A(n_413), .Y(n_770) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g425 ( .A(n_415), .Y(n_425) );
INVx2_ASAP7_75t_L g985 ( .A(n_415), .Y(n_985) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_415), .Y(n_1053) );
INVx8_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI221xp5_ASAP7_75t_SL g748 ( .A1(n_418), .A2(n_749), .B1(n_752), .B2(n_756), .C(n_757), .Y(n_748) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
AND2x4_ASAP7_75t_L g456 ( .A(n_419), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g755 ( .A(n_421), .Y(n_755) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_422), .Y(n_635) );
BUFx3_ASAP7_75t_L g689 ( .A(n_422), .Y(n_689) );
BUFx6f_ASAP7_75t_L g843 ( .A(n_422), .Y(n_843) );
AND2x4_ASAP7_75t_L g845 ( .A(n_422), .B(n_846), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_425), .A2(n_512), .B1(n_514), .B2(n_544), .C(n_546), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_425), .A2(n_546), .B1(n_706), .B2(n_707), .C(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_425), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_427), .A2(n_550), .B1(n_552), .B2(n_553), .C(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g1046 ( .A(n_429), .Y(n_1046) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g636 ( .A(n_430), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g847 ( .A(n_431), .Y(n_847) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g629 ( .A(n_436), .Y(n_629) );
INVx2_ASAP7_75t_L g1207 ( .A(n_436), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g1582 ( .A(n_436), .Y(n_1582) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g676 ( .A(n_439), .Y(n_676) );
INVx2_ASAP7_75t_L g1589 ( .A(n_439), .Y(n_1589) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g562 ( .A(n_440), .Y(n_562) );
INVx3_ASAP7_75t_L g619 ( .A(n_440), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_443), .A2(n_446), .B1(n_691), .B2(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1592 ( .A1(n_443), .A2(n_446), .B1(n_1593), .B2(n_1594), .Y(n_1592) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g760 ( .A(n_445), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_446), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_446), .A2(n_565), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_446), .A2(n_565), .B1(n_740), .B2(n_741), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_446), .A2(n_565), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_446), .A2(n_565), .B1(n_1071), .B2(n_1072), .Y(n_1098) );
CKINVDCx11_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g1524 ( .A(n_448), .Y(n_1524) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g534 ( .A(n_451), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_451), .A2(n_456), .B1(n_763), .B2(n_764), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_451), .A2(n_456), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_452), .Y(n_750) );
AND2x4_ASAP7_75t_L g854 ( .A(n_452), .B(n_855), .Y(n_854) );
BUFx2_ASAP7_75t_L g875 ( .A(n_452), .Y(n_875) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_452), .Y(n_880) );
INVx1_ASAP7_75t_L g932 ( .A(n_452), .Y(n_932) );
BUFx2_ASAP7_75t_L g939 ( .A(n_452), .Y(n_939) );
BUFx6f_ASAP7_75t_L g1199 ( .A(n_452), .Y(n_1199) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g535 ( .A(n_456), .Y(n_535) );
INVx1_ASAP7_75t_L g941 ( .A(n_457), .Y(n_941) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g769 ( .A(n_458), .Y(n_769) );
OAI31xp33_ASAP7_75t_L g611 ( .A1(n_459), .A2(n_612), .A3(n_613), .B(n_627), .Y(n_611) );
OAI31xp33_ASAP7_75t_L g670 ( .A1(n_459), .A2(n_671), .A3(n_672), .B(n_681), .Y(n_670) );
OAI31xp33_ASAP7_75t_L g1088 ( .A1(n_459), .A2(n_1089), .A3(n_1099), .B(n_1109), .Y(n_1088) );
OAI21xp5_ASAP7_75t_L g1192 ( .A1(n_459), .A2(n_1193), .B(n_1202), .Y(n_1192) );
BUFx8_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g1459 ( .A(n_460), .Y(n_1459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g837 ( .A(n_461), .B(n_838), .Y(n_837) );
AND2x4_ASAP7_75t_L g980 ( .A(n_461), .B(n_838), .Y(n_980) );
AOI33xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_468), .A3(n_474), .B1(n_481), .B2(n_484), .B3(n_491), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_464), .Y(n_889) );
OAI22xp5_ASAP7_75t_SL g1019 ( .A1(n_464), .A2(n_662), .B1(n_1020), .B2(n_1027), .Y(n_1019) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g777 ( .A(n_466), .Y(n_777) );
BUFx3_ASAP7_75t_L g1488 ( .A(n_466), .Y(n_1488) );
INVx1_ASAP7_75t_L g838 ( .A(n_467), .Y(n_838) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_470), .Y(n_1003) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g811 ( .A(n_471), .Y(n_811) );
INVx2_ASAP7_75t_L g921 ( .A(n_471), .Y(n_921) );
BUFx6f_ASAP7_75t_L g947 ( .A(n_471), .Y(n_947) );
INVx1_ASAP7_75t_L g1168 ( .A(n_471), .Y(n_1168) );
INVx2_ASAP7_75t_SL g1186 ( .A(n_471), .Y(n_1186) );
AOI222xp33_ASAP7_75t_L g823 ( .A1(n_472), .A2(n_824), .B1(n_825), .B2(n_826), .C1(n_831), .C2(n_832), .Y(n_823) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g483 ( .A(n_473), .Y(n_483) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_473), .Y(n_785) );
INVx2_ASAP7_75t_SL g895 ( .A(n_473), .Y(n_895) );
AND2x4_ASAP7_75t_L g1494 ( .A(n_473), .B(n_1467), .Y(n_1494) );
AND2x4_ASAP7_75t_L g1496 ( .A(n_473), .B(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_476), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g999 ( .A(n_476), .Y(n_999) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_479), .A2(n_505), .B1(n_507), .B2(n_508), .Y(n_504) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g604 ( .A(n_480), .Y(n_604) );
INVx1_ASAP7_75t_L g703 ( .A(n_480), .Y(n_703) );
BUFx3_ASAP7_75t_L g1478 ( .A(n_480), .Y(n_1478) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g585 ( .A(n_487), .Y(n_585) );
INVx1_ASAP7_75t_L g602 ( .A(n_487), .Y(n_602) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g892 ( .A(n_489), .Y(n_892) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_490), .Y(n_661) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_490), .Y(n_668) );
AND2x6_ASAP7_75t_L g822 ( .A(n_490), .B(n_809), .Y(n_822) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_490), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_491), .Y(n_662) );
BUFx4f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx4_ASAP7_75t_L g525 ( .A(n_492), .Y(n_525) );
BUFx4f_ASAP7_75t_L g900 ( .A(n_492), .Y(n_900) );
AOI33xp33_ASAP7_75t_L g997 ( .A1(n_492), .A2(n_889), .A3(n_998), .B1(n_1001), .B2(n_1002), .B3(n_1006), .Y(n_997) );
INVx1_ASAP7_75t_L g1475 ( .A(n_493), .Y(n_1475) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND4x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_530), .C(n_532), .D(n_570), .Y(n_499) );
NOR3xp33_ASAP7_75t_SL g500 ( .A(n_501), .B(n_502), .C(n_526), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g1554 ( .A(n_501), .B(n_1555), .C(n_1574), .Y(n_1554) );
OAI33xp33_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .A3(n_509), .B1(n_515), .B2(n_520), .B3(n_525), .Y(n_502) );
OAI33xp33_ASAP7_75t_L g583 ( .A1(n_503), .A2(n_584), .A3(n_589), .B1(n_594), .B2(n_601), .B3(n_606), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_503), .A2(n_655), .B1(n_662), .B2(n_663), .Y(n_654) );
OAI33xp33_ASAP7_75t_L g700 ( .A1(n_503), .A2(n_525), .A3(n_701), .B1(n_705), .B2(n_708), .B3(n_711), .Y(n_700) );
INVx1_ASAP7_75t_SL g1180 ( .A(n_503), .Y(n_1180) );
OAI33xp33_ASAP7_75t_L g1555 ( .A1(n_503), .A2(n_525), .A3(n_1556), .B1(n_1561), .B2(n_1565), .B3(n_1568), .Y(n_1555) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_505), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx3_ASAP7_75t_L g891 ( .A(n_506), .Y(n_891) );
INVx1_ASAP7_75t_L g1569 ( .A(n_506), .Y(n_1569) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_507), .A2(n_508), .B1(n_538), .B2(n_539), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_510), .A2(n_656), .B1(n_657), .B2(n_659), .C(n_660), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_510), .A2(n_664), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g1561 ( .A1(n_510), .A2(n_1562), .B1(n_1563), .B2(n_1564), .Y(n_1561) );
BUFx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g517 ( .A(n_511), .Y(n_517) );
OR2x2_ASAP7_75t_L g977 ( .A(n_511), .B(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g1023 ( .A(n_511), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g515 ( .A1(n_513), .A2(n_516), .B1(n_518), .B2(n_519), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_516), .A2(n_590), .B1(n_591), .B2(n_593), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_516), .A2(n_597), .B1(n_706), .B2(n_707), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_516), .A2(n_657), .B1(n_709), .B2(n_710), .Y(n_708) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g574 ( .A(n_517), .Y(n_574) );
INVx2_ASAP7_75t_L g595 ( .A(n_517), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g1556 ( .A1(n_521), .A2(n_1557), .B1(n_1558), .B2(n_1560), .Y(n_1556) );
INVx2_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI31xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_536), .A3(n_548), .B(n_567), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_538), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_538), .A2(n_674), .B1(n_675), .B2(n_677), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_538), .A2(n_702), .B1(n_704), .B2(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g858 ( .A(n_542), .Y(n_858) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g1539 ( .A(n_551), .Y(n_1539) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1103 ( .A(n_554), .Y(n_1103) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_561), .A2(n_1465), .B1(n_1471), .B2(n_1534), .Y(n_1537) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g727 ( .A(n_562), .Y(n_727) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_562), .Y(n_751) );
INVx2_ASAP7_75t_L g1155 ( .A(n_562), .Y(n_1155) );
OAI31xp33_ASAP7_75t_L g721 ( .A1(n_567), .A2(n_722), .A3(n_723), .B(n_733), .Y(n_721) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
CKINVDCx8_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
OAI31xp33_ASAP7_75t_L g1035 ( .A1(n_569), .A2(n_1036), .A3(n_1050), .B(n_1062), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g898 ( .A(n_577), .Y(n_898) );
BUFx4f_ASAP7_75t_L g924 ( .A(n_577), .Y(n_924) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_577), .B(n_1467), .Y(n_1466) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND4x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_609), .C(n_611), .D(n_640), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g1477 ( .A(n_585), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_586), .A2(n_588), .B1(n_615), .B2(n_618), .Y(n_614) );
INVx1_ASAP7_75t_L g899 ( .A(n_587), .Y(n_899) );
INVx1_ASAP7_75t_L g1000 ( .A(n_587), .Y(n_1000) );
INVx1_ASAP7_75t_L g1572 ( .A(n_587), .Y(n_1572) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
OAI21xp33_ASAP7_75t_SL g620 ( .A1(n_593), .A2(n_621), .B(n_622), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_600), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_595), .A2(n_1028), .B1(n_1029), .B2(n_1031), .C(n_1032), .Y(n_1027) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx2_ASAP7_75t_L g665 ( .A(n_599), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI33xp33_ASAP7_75t_L g774 ( .A1(n_607), .A2(n_775), .A3(n_778), .B1(n_780), .B2(n_784), .B3(n_786), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g944 ( .A(n_607), .B(n_945), .C(n_948), .Y(n_944) );
INVx1_ASAP7_75t_L g1172 ( .A(n_607), .Y(n_1172) );
AOI33xp33_ASAP7_75t_L g1179 ( .A1(n_607), .A2(n_1180), .A3(n_1181), .B1(n_1182), .B2(n_1183), .B3(n_1187), .Y(n_1179) );
OAI221xp5_ASAP7_75t_L g1586 ( .A1(n_615), .A2(n_1587), .B1(n_1588), .B2(n_1590), .C(n_1591), .Y(n_1586) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_619), .Y(n_1060) );
INVx2_ASAP7_75t_L g1159 ( .A(n_619), .Y(n_1159) );
AND2x4_ASAP7_75t_L g1509 ( .A(n_619), .B(n_1510), .Y(n_1509) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_621), .A2(n_659), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g1152 ( .A(n_624), .Y(n_1152) );
INVx1_ASAP7_75t_L g855 ( .A(n_626), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .C(n_633), .Y(n_628) );
INVx1_ASAP7_75t_L g1057 ( .A(n_629), .Y(n_1057) );
BUFx3_ASAP7_75t_L g871 ( .A(n_634), .Y(n_871) );
INVx2_ASAP7_75t_SL g873 ( .A(n_635), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_1009), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_800), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_743), .B2(n_799), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AO22x2_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_696), .B1(n_697), .B2(n_742), .Y(n_648) );
INVx1_ASAP7_75t_L g742 ( .A(n_649), .Y(n_742) );
AND4x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .C(n_670), .D(n_693), .Y(n_650) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g1030 ( .A(n_658), .Y(n_1030) );
INVx2_ASAP7_75t_SL g713 ( .A(n_661), .Y(n_713) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1097 ( .A(n_680), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1515 ( .A(n_680), .B(n_1510), .Y(n_1515) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_685), .A2(n_735), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_734) );
INVx2_ASAP7_75t_SL g876 ( .A(n_685), .Y(n_876) );
INVx1_ASAP7_75t_L g884 ( .A(n_688), .Y(n_884) );
AND2x6_ASAP7_75t_L g1512 ( .A(n_689), .B(n_1510), .Y(n_1512) );
NAND2x1p5_ASAP7_75t_L g1526 ( .A(n_689), .B(n_1521), .Y(n_1526) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND4x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_716), .C(n_719), .D(n_721), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g933 ( .A(n_727), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_727), .A2(n_1205), .B1(n_1206), .B2(n_1207), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g1529 ( .A1(n_729), .A2(n_1052), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
OAI22xp33_ASAP7_75t_L g1538 ( .A1(n_729), .A2(n_1462), .B1(n_1495), .B2(n_1539), .Y(n_1538) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_735), .A2(n_1106), .B1(n_1107), .B2(n_1108), .Y(n_1105) );
INVx2_ASAP7_75t_L g799 ( .A(n_743), .Y(n_799) );
XOR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_798), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .C(n_773), .Y(n_744) );
AOI31xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_762), .A3(n_765), .B(n_771), .Y(n_747) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g1161 ( .A(n_755), .Y(n_1161) );
NAND2x1p5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_759), .A2(n_1143), .B1(n_1190), .B2(n_1191), .Y(n_1211) );
NAND2x1_ASAP7_75t_SL g1520 ( .A(n_759), .B(n_1521), .Y(n_1520) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g1094 ( .A(n_769), .Y(n_1094) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OAI31xp33_ASAP7_75t_L g1577 ( .A1(n_772), .A2(n_1578), .A3(n_1579), .B(n_1585), .Y(n_1577) );
NAND4xp25_ASAP7_75t_L g773 ( .A(n_774), .B(n_787), .C(n_792), .D(n_795), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_775), .B(n_919), .C(n_923), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_775), .B(n_1163), .C(n_1164), .Y(n_1162) );
INVx3_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx3_ASAP7_75t_L g922 ( .A(n_783), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_789), .A2(n_791), .B1(n_1081), .B2(n_1082), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
XNOR2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_901), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI211x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_836), .B(n_839), .C(n_866), .Y(n_804) );
NAND4xp25_ASAP7_75t_SL g805 ( .A(n_806), .B(n_816), .C(n_823), .D(n_833), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_812), .B2(n_813), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_808), .A2(n_818), .B1(n_912), .B2(n_913), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_808), .A2(n_818), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AND2x4_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
INVx1_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_810), .B(n_1123), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_813), .A2(n_822), .B1(n_915), .B2(n_916), .Y(n_914) );
CKINVDCx6p67_ASAP7_75t_R g974 ( .A(n_813), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_813), .A2(n_822), .B1(n_1131), .B2(n_1132), .Y(n_1130) );
INVx1_ASAP7_75t_L g835 ( .A(n_814), .Y(n_835) );
INVx1_ASAP7_75t_L g978 ( .A(n_814), .Y(n_978) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_821), .B2(n_822), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_817), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_860) );
INVx4_ASAP7_75t_L g979 ( .A(n_818), .Y(n_979) );
AND2x4_ASAP7_75t_L g828 ( .A(n_819), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx4_ASAP7_75t_L g975 ( .A(n_822), .Y(n_975) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_828), .A2(n_832), .B1(n_970), .B2(n_971), .Y(n_969) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g1123 ( .A(n_830), .Y(n_1123) );
INVx3_ASAP7_75t_L g910 ( .A(n_832), .Y(n_910) );
INVx5_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
AOI211xp5_ASAP7_75t_L g905 ( .A1(n_834), .A2(n_906), .B(n_907), .C(n_909), .Y(n_905) );
CKINVDCx8_ASAP7_75t_R g972 ( .A(n_834), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g1119 ( .A(n_834), .B(n_1120), .Y(n_1119) );
AOI221x1_ASAP7_75t_L g1117 ( .A1(n_836), .A2(n_1118), .B1(n_1133), .B2(n_1148), .C(n_1149), .Y(n_1117) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
AO211x2_ASAP7_75t_L g903 ( .A1(n_837), .A2(n_904), .B(n_917), .C(n_951), .Y(n_903) );
AOI31xp33_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_853), .A3(n_860), .B(n_865), .Y(n_839) );
AOI211xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_844), .B(n_845), .C(n_848), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_843), .Y(n_943) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_843), .Y(n_1045) );
AOI211xp5_ASAP7_75t_L g952 ( .A1(n_845), .A2(n_872), .B(n_953), .C(n_954), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g982 ( .A(n_845), .B(n_983), .C(n_987), .Y(n_982) );
CKINVDCx11_ASAP7_75t_R g1147 ( .A(n_845), .Y(n_1147) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVxp67_ASAP7_75t_L g1144 ( .A(n_847), .Y(n_1144) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g955 ( .A(n_850), .Y(n_955) );
INVx2_ASAP7_75t_L g984 ( .A(n_850), .Y(n_984) );
INVx1_ASAP7_75t_L g1143 ( .A(n_852), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_856), .B1(n_857), .B2(n_859), .Y(n_853) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_854), .A2(n_957), .B1(n_958), .B2(n_959), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g988 ( .A1(n_854), .A2(n_958), .B1(n_989), .B2(n_990), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_854), .A2(n_857), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
AND2x4_ASAP7_75t_L g857 ( .A(n_855), .B(n_858), .Y(n_857) );
AND2x4_ASAP7_75t_L g958 ( .A(n_855), .B(n_858), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_861), .A2(n_913), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_861), .A2(n_962), .B1(n_1129), .B2(n_1146), .Y(n_1145) );
INVx4_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx5_ASAP7_75t_L g962 ( .A(n_864), .Y(n_962) );
AOI31xp33_ASAP7_75t_L g951 ( .A1(n_865), .A2(n_952), .A3(n_956), .B(n_960), .Y(n_951) );
AO21x1_ASAP7_75t_SL g981 ( .A1(n_865), .A2(n_982), .B(n_988), .Y(n_981) );
CKINVDCx16_ASAP7_75t_R g1148 ( .A(n_865), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_888), .Y(n_866) );
AOI33xp33_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_870), .A3(n_874), .B1(n_877), .B2(n_882), .B3(n_886), .Y(n_867) );
BUFx3_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NAND3xp33_ASAP7_75t_L g937 ( .A(n_869), .B(n_938), .C(n_942), .Y(n_937) );
INVx2_ASAP7_75t_SL g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g885 ( .A(n_873), .Y(n_885) );
INVx3_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_880), .B(n_1510), .Y(n_1517) );
INVx1_ASAP7_75t_L g1108 ( .A(n_881), .Y(n_1108) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AOI222xp33_ASAP7_75t_L g1137 ( .A1(n_885), .A2(n_1138), .B1(n_1139), .B2(n_1140), .C1(n_1141), .C2(n_1142), .Y(n_1137) );
AOI33xp33_ASAP7_75t_L g991 ( .A1(n_886), .A2(n_992), .A3(n_993), .B1(n_994), .B2(n_995), .B3(n_996), .Y(n_991) );
INVx6_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx5_ASAP7_75t_L g936 ( .A(n_887), .Y(n_936) );
AOI33xp33_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .A3(n_893), .B1(n_896), .B2(n_897), .B3(n_900), .Y(n_888) );
AOI33xp33_ASAP7_75t_L g1073 ( .A1(n_889), .A2(n_900), .A3(n_1074), .B1(n_1075), .B2(n_1076), .B3(n_1077), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_894), .B(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g1474 ( .A(n_895), .Y(n_1474) );
XNOR2x1_ASAP7_75t_L g901 ( .A(n_902), .B(n_963), .Y(n_901) );
NAND3xp33_ASAP7_75t_L g904 ( .A(n_905), .B(n_911), .C(n_914), .Y(n_904) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
NAND4xp25_ASAP7_75t_L g917 ( .A(n_918), .B(n_929), .C(n_937), .D(n_944), .Y(n_917) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g950 ( .A(n_926), .Y(n_950) );
INVx2_ASAP7_75t_SL g1559 ( .A(n_926), .Y(n_1559) );
INVx2_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g1491 ( .A(n_928), .Y(n_1491) );
NAND3xp33_ASAP7_75t_L g929 ( .A(n_930), .B(n_934), .C(n_936), .Y(n_929) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g1536 ( .A(n_933), .Y(n_1536) );
NAND3xp33_ASAP7_75t_L g1150 ( .A(n_936), .B(n_1151), .C(n_1153), .Y(n_1150) );
CKINVDCx8_ASAP7_75t_R g1540 ( .A(n_936), .Y(n_1540) );
INVx1_ASAP7_75t_L g1042 ( .A(n_940), .Y(n_1042) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx4_ASAP7_75t_L g1490 ( .A(n_947), .Y(n_1490) );
INVx1_ASAP7_75t_L g1140 ( .A(n_955), .Y(n_1140) );
AND4x1_ASAP7_75t_L g964 ( .A(n_965), .B(n_981), .C(n_991), .D(n_997), .Y(n_964) );
NAND4xp25_ASAP7_75t_L g1008 ( .A(n_965), .B(n_981), .C(n_991), .D(n_997), .Y(n_1008) );
OAI31xp33_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_973), .A3(n_976), .B(n_980), .Y(n_965) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_969), .C(n_972), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g1156 ( .A(n_992), .B(n_1157), .C(n_1160), .Y(n_1156) );
BUFx6f_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
AO22x2_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1012), .B1(n_1112), .B2(n_1113), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
AO22x1_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1066), .B1(n_1110), .B2(n_1111), .Y(n_1012) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1013), .Y(n_1111) );
AND4x1_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1033), .C(n_1035), .D(n_1063), .Y(n_1014) );
NOR3xp33_ASAP7_75t_SL g1015 ( .A(n_1016), .B(n_1017), .C(n_1019), .Y(n_1015) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1041), .B1(n_1042), .B2(n_1043), .C(n_1044), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx2_ASAP7_75t_L g1534 ( .A(n_1039), .Y(n_1534) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_1040), .Y(n_1091) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1058), .B1(n_1059), .B2(n_1061), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_1060), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1066), .Y(n_1110) );
AND3x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1086), .C(n_1088), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1079), .Y(n_1068) );
NAND3xp33_ASAP7_75t_SL g1069 ( .A(n_1070), .B(n_1073), .C(n_1078), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1083), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1090 ( .A1(n_1081), .A2(n_1085), .B1(n_1091), .B2(n_1092), .C(n_1095), .Y(n_1090) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
OAI22x1_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1115), .B1(n_1174), .B2(n_1175), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1117), .Y(n_1173) );
NAND3xp33_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1127), .C(n_1130), .Y(n_1118) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1563 ( .A(n_1126), .Y(n_1563) );
NAND4xp25_ASAP7_75t_SL g1133 ( .A(n_1134), .B(n_1137), .C(n_1145), .D(n_1147), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
NAND4xp25_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1156), .C(n_1162), .D(n_1166), .Y(n_1149) );
A2O1A1Ixp33_ASAP7_75t_L g1208 ( .A1(n_1152), .A2(n_1209), .B(n_1210), .C(n_1212), .Y(n_1208) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1154), .Y(n_1583) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1169), .C(n_1171), .Y(n_1166) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1174 ( .A(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
NAND4xp75_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1192), .C(n_1213), .D(n_1215), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1189), .Y(n_1178) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1197), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1452), .B1(n_1454), .B2(n_1541), .C(n_1545), .Y(n_1218) );
AND3x1_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1410), .C(n_1440), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1309), .B1(n_1317), .B2(n_1361), .C(n_1388), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1294), .Y(n_1221) );
O2A1O1Ixp33_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1275), .B(n_1278), .C(n_1283), .Y(n_1222) );
AOI21xp5_ASAP7_75t_L g1422 ( .A1(n_1223), .A2(n_1423), .B(n_1425), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1251), .Y(n_1223) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1224), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1224), .B(n_1307), .Y(n_1409) );
INVx2_ASAP7_75t_L g1425 ( .A(n_1224), .Y(n_1425) );
INVx2_ASAP7_75t_SL g1224 ( .A(n_1225), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1225), .B(n_1297), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_1225), .B(n_1279), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1225), .B(n_1280), .Y(n_1322) );
HB1xp67_ASAP7_75t_L g1338 ( .A(n_1225), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1225), .B(n_1310), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_1226), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1226), .B(n_1279), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1226), .B(n_1280), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1241), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1235), .B1(n_1236), .B2(n_1240), .Y(n_1227) );
BUFx3_ASAP7_75t_L g1355 ( .A(n_1228), .Y(n_1355) );
BUFx6f_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_1229), .A2(n_1238), .B1(n_1265), .B2(n_1266), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1231), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1230), .B(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1230), .Y(n_1258) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1231), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1234), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1604 ( .A(n_1232), .Y(n_1604) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1234), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1236), .Y(n_1357) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1239), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1247), .B1(n_1248), .B2(n_1250), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
BUFx3_ASAP7_75t_L g1352 ( .A(n_1243), .Y(n_1352) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1246), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1244), .B(n_1246), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1602 ( .A(n_1244), .Y(n_1602) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
AND2x4_ASAP7_75t_L g1249 ( .A(n_1245), .B(n_1246), .Y(n_1249) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1248), .Y(n_1316) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1248), .Y(n_1453) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1267), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1252), .B(n_1307), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1252), .B(n_1272), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1252), .B(n_1286), .Y(n_1406) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1253), .B(n_1307), .Y(n_1374) );
NOR2xp33_ASAP7_75t_L g1411 ( .A(n_1253), .B(n_1412), .Y(n_1411) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1253), .B(n_1350), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1263), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1254), .B(n_1263), .Y(n_1277) );
INVx2_ASAP7_75t_L g1291 ( .A(n_1254), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1254), .B(n_1305), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1254), .B(n_1304), .Y(n_1371) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1254), .B(n_1305), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1261), .Y(n_1254) );
AND2x4_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1258), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1259 ( .A(n_1258), .B(n_1260), .Y(n_1259) );
BUFx2_ASAP7_75t_L g1314 ( .A(n_1259), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1263), .B(n_1291), .Y(n_1290) );
INVx2_ASAP7_75t_SL g1304 ( .A(n_1263), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1263), .B(n_1272), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1263), .B(n_1305), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1267), .B(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1267), .B(n_1290), .Y(n_1321) );
INVxp67_ASAP7_75t_SL g1372 ( .A(n_1267), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1271), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1268), .B(n_1277), .Y(n_1287) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1268), .Y(n_1297) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1268), .Y(n_1307) );
BUFx2_ASAP7_75t_L g1326 ( .A(n_1268), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1268), .B(n_1305), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1268), .B(n_1332), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1271), .B(n_1290), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1271), .B(n_1277), .Y(n_1334) );
NOR2x1_ASAP7_75t_L g1382 ( .A(n_1271), .B(n_1304), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g1435 ( .A(n_1271), .B(n_1291), .Y(n_1435) );
BUFx2_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVxp67_ASAP7_75t_L g1286 ( .A(n_1272), .Y(n_1286) );
BUFx3_ASAP7_75t_L g1305 ( .A(n_1272), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1274), .Y(n_1272) );
AOI21xp5_ASAP7_75t_L g1445 ( .A1(n_1275), .A2(n_1425), .B(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1277), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1277), .B(n_1349), .Y(n_1348) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_1277), .A2(n_1369), .B1(n_1370), .B2(n_1372), .C(n_1373), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1277), .B(n_1307), .Y(n_1431) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1278), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1278), .B(n_1326), .Y(n_1443) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1279), .B(n_1312), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_1279), .B(n_1395), .Y(n_1394) );
A2O1A1Ixp33_ASAP7_75t_SL g1440 ( .A1(n_1279), .A2(n_1358), .B(n_1441), .C(n_1442), .Y(n_1440) );
INVx3_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1280), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_1280), .B(n_1312), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1280), .B(n_1311), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
AOI21xp5_ASAP7_75t_L g1283 ( .A1(n_1284), .A2(n_1288), .B(n_1292), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_1285), .A2(n_1341), .B1(n_1428), .B2(n_1430), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1286), .B(n_1290), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1286), .B(n_1371), .Y(n_1421) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1290), .B(n_1307), .Y(n_1417) );
A2O1A1Ixp33_ASAP7_75t_L g1376 ( .A1(n_1291), .A2(n_1377), .B(n_1380), .C(n_1383), .Y(n_1376) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
O2A1O1Ixp33_ASAP7_75t_L g1347 ( .A1(n_1293), .A2(n_1348), .B(n_1351), .C(n_1358), .Y(n_1347) );
OAI21xp5_ASAP7_75t_L g1389 ( .A1(n_1293), .A2(n_1296), .B(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1293), .B(n_1297), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1293), .B(n_1448), .Y(n_1447) );
AOI211xp5_ASAP7_75t_SL g1294 ( .A1(n_1295), .A2(n_1296), .B(n_1299), .C(n_1301), .Y(n_1294) );
A2O1A1Ixp33_ASAP7_75t_SL g1419 ( .A1(n_1295), .A2(n_1418), .B(n_1420), .C(n_1422), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1297), .B(n_1435), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1298), .B(n_1300), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g1444 ( .A(n_1298), .B(n_1336), .Y(n_1444) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1300), .Y(n_1369) );
NOR2xp33_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1306), .Y(n_1301) );
OAI221xp5_ASAP7_75t_L g1317 ( .A1(n_1302), .A2(n_1318), .B1(n_1339), .B2(n_1340), .C(n_1342), .Y(n_1317) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1305), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1305), .B(n_1320), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1305), .B(n_1431), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1307), .B(n_1332), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1307), .B(n_1336), .Y(n_1335) );
OAI21xp33_ASAP7_75t_L g1404 ( .A1(n_1307), .A2(n_1330), .B(n_1405), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1308), .B(n_1310), .Y(n_1341) );
AOI221xp5_ASAP7_75t_L g1400 ( .A1(n_1308), .A2(n_1343), .B1(n_1401), .B2(n_1404), .C(n_1407), .Y(n_1400) );
AOI21xp5_ASAP7_75t_L g1416 ( .A1(n_1308), .A2(n_1417), .B(n_1418), .Y(n_1416) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1310), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1311), .Y(n_1360) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1312), .Y(n_1339) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1312), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1315), .Y(n_1312) );
AOI22xp5_ASAP7_75t_L g1361 ( .A1(n_1318), .A2(n_1362), .B1(n_1365), .B2(n_1376), .Y(n_1361) );
AND3x1_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1323), .C(n_1333), .Y(n_1318) );
OAI21xp5_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1321), .B(n_1322), .Y(n_1319) );
AOI221xp5_ASAP7_75t_L g1342 ( .A1(n_1321), .A2(n_1343), .B1(n_1345), .B2(n_1346), .C(n_1347), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1322), .B(n_1379), .Y(n_1378) );
A2O1A1Ixp33_ASAP7_75t_L g1432 ( .A1(n_1322), .A2(n_1351), .B(n_1433), .C(n_1436), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1327), .B1(n_1328), .B2(n_1331), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AOI21xp5_ASAP7_75t_L g1436 ( .A1(n_1325), .A2(n_1329), .B(n_1405), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1327), .Y(n_1325) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1326), .Y(n_1379) );
NAND2xp5_ASAP7_75t_SL g1402 ( .A(n_1326), .B(n_1403), .Y(n_1402) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_1327), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1330), .Y(n_1328) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1331), .Y(n_1415) );
OAI21xp33_ASAP7_75t_L g1333 ( .A1(n_1334), .A2(n_1335), .B(n_1337), .Y(n_1333) );
AOI221xp5_ASAP7_75t_L g1392 ( .A1(n_1334), .A2(n_1335), .B1(n_1346), .B2(n_1393), .C(n_1396), .Y(n_1392) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1335), .Y(n_1414) );
INVxp67_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
NOR2xp33_ASAP7_75t_L g1450 ( .A(n_1338), .B(n_1451), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1339), .B(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1341), .B(n_1345), .Y(n_1439) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1346), .Y(n_1429) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1351), .B(n_1359), .Y(n_1358) );
INVx3_ASAP7_75t_L g1364 ( .A(n_1351), .Y(n_1364) );
AOI31xp33_ASAP7_75t_L g1388 ( .A1(n_1351), .A2(n_1389), .A3(n_1392), .B(n_1400), .Y(n_1388) );
INVx3_ASAP7_75t_L g1418 ( .A(n_1351), .Y(n_1418) );
OAI22xp33_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1355), .B1(n_1356), .B2(n_1357), .Y(n_1353) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
AOI211xp5_ASAP7_75t_L g1365 ( .A1(n_1360), .A2(n_1366), .B(n_1368), .C(n_1375), .Y(n_1365) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1360), .Y(n_1398) );
NAND3xp33_ASAP7_75t_SL g1408 ( .A(n_1360), .B(n_1371), .C(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g1396 ( .A(n_1370), .B(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
AOI21xp33_ASAP7_75t_L g1437 ( .A1(n_1375), .A2(n_1438), .B(n_1439), .Y(n_1437) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1379), .B(n_1382), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1379), .B(n_1421), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1379), .B(n_1403), .Y(n_1424) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1386), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1387), .B(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
OR2x2_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1399), .Y(n_1397) );
A2O1A1Ixp33_ASAP7_75t_L g1413 ( .A1(n_1399), .A2(n_1414), .B(n_1415), .C(n_1416), .Y(n_1413) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
O2A1O1Ixp33_ASAP7_75t_L g1410 ( .A1(n_1411), .A2(n_1413), .B(n_1419), .C(n_1426), .Y(n_1410) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1420), .Y(n_1441) );
INVx2_ASAP7_75t_L g1448 ( .A(n_1421), .Y(n_1448) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
NAND3xp33_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1432), .C(n_1437), .Y(n_1426) );
INVxp67_ASAP7_75t_SL g1433 ( .A(n_1434), .Y(n_1433) );
OAI211xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1444), .B(n_1445), .C(n_1449), .Y(n_1442) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
HB1xp67_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1504), .Y(n_1457) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_1459), .A2(n_1460), .B1(n_1498), .B2(n_1499), .Y(n_1458) );
NAND3xp33_ASAP7_75t_SL g1460 ( .A(n_1461), .B(n_1468), .C(n_1485), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_1462), .A2(n_1463), .B1(n_1465), .B2(n_1466), .Y(n_1461) );
INVx6_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
AOI221xp5_ASAP7_75t_L g1468 ( .A1(n_1469), .A2(n_1471), .B1(n_1472), .B2(n_1476), .C(n_1479), .Y(n_1468) );
INVx4_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx4_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx2_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g1485 ( .A1(n_1486), .A2(n_1489), .B1(n_1492), .B2(n_1495), .C(n_1496), .Y(n_1485) );
INVx3_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
INVx2_ASAP7_75t_SL g1493 ( .A(n_1494), .Y(n_1493) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
AND2x4_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1503), .Y(n_1500) );
INVx3_ASAP7_75t_L g1521 ( .A(n_1502), .Y(n_1521) );
NOR3xp33_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1518), .C(n_1527), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1513), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_1507), .A2(n_1508), .B1(n_1511), .B2(n_1512), .Y(n_1506) );
BUFx2_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_1514), .A2(n_1515), .B1(n_1516), .B2(n_1517), .Y(n_1513) );
HB1xp67_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
NAND2x1p5_ASAP7_75t_L g1523 ( .A(n_1521), .B(n_1524), .Y(n_1523) );
BUFx4f_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
BUFx2_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
OAI33xp33_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1529), .A3(n_1532), .B1(n_1537), .B2(n_1538), .B3(n_1540), .Y(n_1527) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_1533), .A2(n_1534), .B1(n_1535), .B2(n_1536), .Y(n_1532) );
INVx2_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
CKINVDCx5p33_ASAP7_75t_R g1547 ( .A(n_1548), .Y(n_1547) );
A2O1A1Ixp33_ASAP7_75t_L g1600 ( .A1(n_1549), .A2(n_1601), .B(n_1603), .C(n_1605), .Y(n_1600) );
INVxp33_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
HB1xp67_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
AND4x1_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1575), .C(n_1577), .D(n_1595), .Y(n_1553) );
OAI22xp5_ASAP7_75t_L g1580 ( .A1(n_1557), .A2(n_1560), .B1(n_1581), .B2(n_1583), .Y(n_1580) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
OAI22xp5_ASAP7_75t_L g1568 ( .A1(n_1569), .A2(n_1570), .B1(n_1571), .B2(n_1573), .Y(n_1568) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
NOR2xp33_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1597), .Y(n_1595) );
BUFx2_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
HB1xp67_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
endmodule