module fake_jpeg_4768_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_9),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_39),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_53),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_58),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_17),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_56),
.Y(n_102)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_25),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_69),
.Y(n_138)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_26),
.B1(n_16),
.B2(n_25),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_15),
.B1(n_31),
.B2(n_18),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_91),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_16),
.B1(n_26),
.B2(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_97),
.B1(n_104),
.B2(n_12),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_96),
.B1(n_106),
.B2(n_108),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_41),
.A2(n_34),
.B1(n_25),
.B2(n_35),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_93),
.B(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_41),
.A2(n_34),
.B1(n_35),
.B2(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_128)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_56),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_30),
.B1(n_31),
.B2(n_29),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_15),
.B1(n_29),
.B2(n_30),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_43),
.B(n_29),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_133),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_47),
.B1(n_31),
.B2(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_125),
.B1(n_132),
.B2(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_42),
.B1(n_29),
.B2(n_15),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_77),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_43),
.B(n_45),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_124),
.CI(n_64),
.CON(n_148),
.SN(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_45),
.B(n_43),
.C(n_18),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_31),
.B1(n_18),
.B2(n_2),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_92),
.B(n_75),
.C(n_63),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_137),
.B(n_77),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_79),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_0),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_61),
.B(n_1),
.C(n_4),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_69),
.C(n_62),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_68),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_5),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_157),
.B1(n_163),
.B2(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_143),
.B(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_150),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_126),
.B1(n_138),
.B2(n_123),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

XOR2x1_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_156),
.Y(n_212)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_103),
.B(n_93),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_131),
.B1(n_126),
.B2(n_113),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_158),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_82),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_99),
.B1(n_70),
.B2(n_106),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_5),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_111),
.B(n_107),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_86),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_171),
.B(n_162),
.Y(n_183)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_74),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_86),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_95),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_107),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_83),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_68),
.C(n_108),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_10),
.C(n_144),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_118),
.A2(n_99),
.B1(n_70),
.B2(n_63),
.Y(n_176)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_88),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_88),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_184),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_148),
.B(n_145),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_161),
.B(n_149),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_130),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_120),
.B1(n_127),
.B2(n_123),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_189),
.A2(n_210),
.B1(n_214),
.B2(n_10),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_119),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_211),
.C(n_191),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_153),
.A2(n_115),
.B1(n_116),
.B2(n_125),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_119),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_200),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_158),
.A2(n_115),
.B1(n_138),
.B2(n_141),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_141),
.B1(n_129),
.B2(n_67),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_199),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_141),
.B1(n_129),
.B2(n_67),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_110),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_215),
.C(n_216),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_10),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_154),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_210)
);

OR2x6_ASAP7_75t_L g211 ( 
.A(n_142),
.B(n_110),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_177),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_166),
.A2(n_8),
.B1(n_10),
.B2(n_145),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_173),
.B(n_8),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_148),
.B(n_156),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_226),
.B(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_224),
.B(n_235),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_161),
.B1(n_157),
.B2(n_168),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_143),
.Y(n_229)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_238),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_174),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_168),
.C(n_171),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_237),
.C(n_216),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_171),
.B(n_149),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_185),
.B(n_150),
.C(n_169),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_243),
.B1(n_201),
.B2(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_184),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_197),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_190),
.Y(n_262)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_244),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_181),
.A2(n_189),
.B1(n_188),
.B2(n_200),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_246),
.B(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_181),
.B1(n_210),
.B2(n_211),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_255),
.B1(n_226),
.B2(n_236),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_195),
.Y(n_251)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_266),
.C(n_222),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_245),
.A2(n_186),
.B1(n_211),
.B2(n_199),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_262),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_269),
.B1(n_217),
.B2(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_265),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_215),
.C(n_208),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_182),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_268),
.CI(n_239),
.CON(n_279),
.SN(n_279)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_233),
.B(n_196),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_193),
.B1(n_180),
.B2(n_187),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_271),
.C(n_273),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_222),
.C(n_234),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_225),
.C(n_241),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_255),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_225),
.C(n_243),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_287),
.C(n_237),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_268),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_281),
.B1(n_226),
.B2(n_249),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_242),
.B1(n_232),
.B2(n_217),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_282),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_250),
.A2(n_219),
.B1(n_226),
.B2(n_235),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_220),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_263),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_219),
.C(n_221),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_256),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_295),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_284),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_294),
.B(n_301),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_271),
.C(n_278),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_249),
.B(n_247),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_299),
.B1(n_261),
.B2(n_292),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_237),
.B(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_299),
.B1(n_276),
.B2(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

AOI221xp5_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_244),
.B1(n_279),
.B2(n_296),
.C(n_246),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_310),
.C(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_264),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_273),
.C(n_284),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_297),
.C(n_295),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_283),
.B1(n_252),
.B2(n_274),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_290),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_319),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_294),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_318),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_251),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_260),
.C(n_248),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_257),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_322),
.B1(n_313),
.B2(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_325),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_309),
.B1(n_304),
.B2(n_230),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_315),
.A2(n_296),
.B1(n_311),
.B2(n_279),
.Y(n_328)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_322),
.B(n_316),
.C(n_306),
.D(n_307),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_331),
.B(n_259),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_307),
.C(n_259),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_334),
.B(n_332),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_326),
.A3(n_258),
.B1(n_267),
.B2(n_253),
.C1(n_257),
.C2(n_240),
.Y(n_334)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_253),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_224),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_213),
.Y(n_338)
);


endmodule