module fake_netlist_5_1625_n_581 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_65, n_78, n_74, n_57, n_96, n_37, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_94, n_38, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_85, n_95, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_81, n_28, n_89, n_70, n_68, n_93, n_72, n_32, n_41, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_581);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_96;
input n_37;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_94;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_85;
input n_95;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_89;
input n_70;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;

output n_581;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_136;
wire n_124;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_493;
wire n_111;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_116;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_105;
wire n_280;
wire n_378;
wire n_551;
wire n_382;
wire n_554;
wire n_254;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_119;
wire n_497;
wire n_559;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_106;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_546;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_104;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_145;
wire n_521;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_114;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_107;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_112;
wire n_542;
wire n_463;
wire n_488;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_511;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_102;
wire n_273;
wire n_161;
wire n_349;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_487;
wire n_495;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_103;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_29),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_26),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g105 ( 
.A(n_6),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_5),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_1),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_79),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_32),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_44),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_51),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_46),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_58),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_37),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_72),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_23),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_L g146 ( 
.A(n_69),
.B(n_33),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_35),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_34),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_36),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_40),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_24),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_19),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_2),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_48),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_20),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_21),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_57),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_31),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_17),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_84),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_61),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_63),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_13),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_73),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_14),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_L g180 ( 
.A(n_55),
.B(n_39),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_38),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_30),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_13),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_22),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

BUFx8_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_27),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_103),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_112),
.B(n_43),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_106),
.B(n_114),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_114),
.A2(n_0),
.B(n_4),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_8),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_131),
.B(n_52),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_157),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_131),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_108),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

XNOR2x2_ASAP7_75t_R g233 ( 
.A(n_111),
.B(n_10),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_188),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_178),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_15),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_143),
.B(n_16),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_154),
.A2(n_18),
.B(n_25),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_102),
.B(n_80),
.Y(n_248)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_109),
.A2(n_18),
.B(n_49),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_110),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_159),
.A2(n_59),
.B1(n_60),
.B2(n_87),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_159),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_118),
.B(n_193),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_108),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_124),
.B(n_172),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_127),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_132),
.B(n_171),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_134),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_140),
.B(n_187),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_192),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_137),
.B(n_138),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_145),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_183),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_209),
.B(n_135),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_137),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_214),
.A2(n_169),
.B1(n_147),
.B2(n_135),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_152),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_177),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_214),
.B(n_177),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_149),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_138),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_194),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_249),
.B(n_160),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_201),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_235),
.B(n_174),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_194),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_239),
.B(n_192),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_231),
.B(n_164),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_235),
.B(n_147),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_194),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_158),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_205),
.B(n_153),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g299 ( 
.A1(n_252),
.A2(n_174),
.B1(n_170),
.B2(n_169),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_254),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_203),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_101),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_220),
.B(n_170),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_217),
.A2(n_125),
.B1(n_128),
.B2(n_120),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_220),
.B(n_128),
.Y(n_309)
);

OR2x6_ASAP7_75t_L g310 ( 
.A(n_215),
.B(n_247),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_199),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_256),
.B(n_258),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_250),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_217),
.B1(n_206),
.B2(n_196),
.Y(n_316)
);

BUFx4f_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_206),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_260),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_281),
.B(n_199),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_267),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_268),
.B(n_240),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_207),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_251),
.Y(n_336)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_253),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_267),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_262),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_299),
.B1(n_287),
.B2(n_305),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_281),
.B(n_180),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_295),
.A2(n_264),
.B(n_259),
.C(n_216),
.Y(n_342)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_271),
.B(n_146),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_305),
.A2(n_196),
.B1(n_237),
.B2(n_119),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_294),
.A2(n_104),
.B1(n_121),
.B2(n_123),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_274),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_282),
.B(n_257),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_259),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_317),
.B(n_290),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_296),
.B(n_311),
.C(n_283),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_283),
.Y(n_358)
);

AO32x1_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_312),
.A3(n_307),
.B1(n_296),
.B2(n_298),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_318),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_340),
.A2(n_328),
.B1(n_327),
.B2(n_347),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_341),
.A2(n_310),
.B1(n_249),
.B2(n_130),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_354),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_298),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_341),
.A2(n_307),
.B(n_312),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_227),
.Y(n_366)
);

BUFx8_ASAP7_75t_SL g367 ( 
.A(n_315),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_306),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_310),
.B1(n_249),
.B2(n_133),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_317),
.A2(n_310),
.B1(n_129),
.B2(n_142),
.Y(n_370)
);

BUFx8_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

O2A1O1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_347),
.A2(n_264),
.B(n_225),
.C(n_242),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_211),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_196),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_227),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_308),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_244),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_325),
.B(n_232),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_246),
.Y(n_380)
);

OR2x6_ASAP7_75t_SL g381 ( 
.A(n_350),
.B(n_233),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_286),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_325),
.B(n_244),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

CKINVDCx11_ASAP7_75t_R g386 ( 
.A(n_320),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_286),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_316),
.B(n_126),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_337),
.A2(n_223),
.B1(n_213),
.B2(n_264),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_226),
.C(n_241),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_344),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_343),
.A2(n_291),
.B(n_288),
.C(n_284),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_345),
.A2(n_291),
.B(n_288),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_320),
.B(n_144),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_320),
.B(n_150),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_335),
.B(n_161),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_353),
.B(n_163),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_210),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_342),
.A2(n_302),
.B(n_292),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_324),
.B(n_261),
.Y(n_405)
);

O2A1O1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_355),
.A2(n_218),
.B(n_243),
.C(n_238),
.Y(n_406)
);

NOR2x1_ASAP7_75t_SL g407 ( 
.A(n_331),
.B(n_203),
.Y(n_407)
);

OR2x6_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_233),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_351),
.A2(n_165),
.B1(n_168),
.B2(n_181),
.Y(n_409)
);

INVx3_ASAP7_75t_SL g410 ( 
.A(n_352),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_236),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

AOI221xp5_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_261),
.B1(n_245),
.B2(n_236),
.C(n_212),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_365),
.A2(n_331),
.B(n_216),
.Y(n_414)
);

AO31x2_ASAP7_75t_L g415 ( 
.A1(n_362),
.A2(n_221),
.A3(n_230),
.B(n_222),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_356),
.B(n_378),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_364),
.A2(n_216),
.B(n_185),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_367),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_361),
.A2(n_223),
.B1(n_213),
.B2(n_257),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_386),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_358),
.A2(n_257),
.B(n_224),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

AOI32xp33_ASAP7_75t_L g424 ( 
.A1(n_379),
.A2(n_245),
.A3(n_228),
.B1(n_212),
.B2(n_230),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_228),
.C(n_223),
.Y(n_425)
);

BUFx12f_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_380),
.A2(n_387),
.B(n_383),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_366),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_404),
.A2(n_377),
.B(n_393),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_376),
.B(n_368),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_375),
.Y(n_432)
);

OAI22x1_ASAP7_75t_L g433 ( 
.A1(n_381),
.A2(n_389),
.B1(n_408),
.B2(n_392),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_370),
.A2(n_382),
.B(n_390),
.Y(n_436)
);

A2O1A1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_373),
.A2(n_406),
.B(n_391),
.C(n_411),
.Y(n_437)
);

BUFx10_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

AO21x2_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_398),
.B(n_359),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_408),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_410),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_L g442 ( 
.A1(n_360),
.A2(n_385),
.B1(n_388),
.B2(n_396),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_388),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_407),
.A2(n_397),
.B(n_360),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_360),
.A2(n_395),
.B(n_359),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_359),
.A2(n_409),
.B(n_388),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_402),
.A2(n_361),
.B1(n_313),
.B2(n_328),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_361),
.A2(n_313),
.B(n_328),
.C(n_340),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_366),
.B(n_322),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g452 ( 
.A1(n_357),
.A2(n_341),
.B(n_362),
.Y(n_452)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

AO31x2_ASAP7_75t_L g456 ( 
.A1(n_362),
.A2(n_369),
.A3(n_403),
.B(n_394),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_399),
.Y(n_457)
);

CKINVDCx11_ASAP7_75t_R g458 ( 
.A(n_381),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_361),
.A2(n_313),
.B(n_328),
.C(n_340),
.Y(n_459)
);

AO31x2_ASAP7_75t_L g460 ( 
.A1(n_362),
.A2(n_369),
.A3(n_403),
.B(n_394),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_386),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_320),
.Y(n_462)
);

AOI221xp5_ASAP7_75t_L g463 ( 
.A1(n_384),
.A2(n_299),
.B1(n_268),
.B2(n_309),
.C(n_304),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_459),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_416),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_463),
.B(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_429),
.Y(n_469)
);

AO31x2_ASAP7_75t_L g470 ( 
.A1(n_445),
.A2(n_447),
.A3(n_427),
.B(n_437),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_461),
.Y(n_471)
);

AOI221xp5_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_430),
.B1(n_423),
.B2(n_457),
.C(n_464),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_432),
.B(n_412),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_421),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_448),
.A2(n_424),
.B(n_420),
.C(n_425),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_424),
.B(n_455),
.Y(n_476)
);

AO31x2_ASAP7_75t_L g477 ( 
.A1(n_414),
.A2(n_418),
.A3(n_422),
.B(n_444),
.Y(n_477)
);

AO31x2_ASAP7_75t_L g478 ( 
.A1(n_415),
.A2(n_452),
.A3(n_460),
.B(n_456),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_443),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_428),
.B(n_440),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_454),
.B(n_442),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_419),
.Y(n_482)
);

INVx3_ASAP7_75t_SL g483 ( 
.A(n_453),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_452),
.A2(n_460),
.B(n_456),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_446),
.A2(n_413),
.B(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_456),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_439),
.B(n_438),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_462),
.A2(n_433),
.B(n_438),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

CKINVDCx9p33_ASAP7_75t_R g490 ( 
.A(n_453),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_417),
.A2(n_426),
.B(n_458),
.Y(n_491)
);

AO31x2_ASAP7_75t_L g492 ( 
.A1(n_445),
.A2(n_369),
.A3(n_362),
.B(n_447),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_428),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_493),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_494),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_466),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_466),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_471),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_476),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_468),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_484),
.Y(n_504)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_494),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_475),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_473),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_469),
.B(n_472),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_470),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_470),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_487),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_470),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_481),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_477),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_479),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_502),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_R g517 ( 
.A(n_505),
.B(n_489),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_496),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_488),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_477),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_480),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_483),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_491),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_482),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_506),
.B(n_474),
.Y(n_527)
);

NOR2x1_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_490),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_497),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_498),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_509),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_512),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_503),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_512),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_516),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_507),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_510),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_532),
.B(n_512),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_514),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_516),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_514),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_523),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_513),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_504),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_537),
.B(n_533),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_539),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_531),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_522),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_542),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_540),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_529),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_544),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_552),
.B(n_536),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_537),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_529),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_541),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_541),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_529),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_547),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_560),
.Y(n_561)
);

AOI21xp33_ASAP7_75t_L g562 ( 
.A1(n_556),
.A2(n_524),
.B(n_520),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_555),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_553),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_557),
.B(n_548),
.Y(n_565)
);

AOI211xp5_ASAP7_75t_L g566 ( 
.A1(n_562),
.A2(n_554),
.B(n_527),
.C(n_524),
.Y(n_566)
);

AOI211xp5_ASAP7_75t_SL g567 ( 
.A1(n_562),
.A2(n_522),
.B(n_527),
.C(n_520),
.Y(n_567)
);

AOI222xp33_ASAP7_75t_L g568 ( 
.A1(n_566),
.A2(n_525),
.B1(n_563),
.B2(n_559),
.C1(n_549),
.C2(n_564),
.Y(n_568)
);

OAI211xp5_ASAP7_75t_SL g569 ( 
.A1(n_568),
.A2(n_567),
.B(n_528),
.C(n_561),
.Y(n_569)
);

NOR2x1_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_528),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_570),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_570),
.B(n_525),
.C(n_499),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_519),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_571),
.B(n_565),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_558),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_573),
.B1(n_526),
.B2(n_561),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_575),
.B(n_548),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_553),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_578),
.A2(n_577),
.B(n_517),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_495),
.B(n_547),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_580),
.A2(n_526),
.B1(n_505),
.B2(n_518),
.Y(n_581)
);


endmodule