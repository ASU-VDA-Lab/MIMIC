module fake_jpeg_19294_n_29 (n_3, n_2, n_1, n_0, n_4, n_5, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx3_ASAP7_75t_SL g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_7),
.B(n_10),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_15),
.B1(n_9),
.B2(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_15),
.B(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_17),
.Y(n_19)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_13),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_12),
.B1(n_14),
.B2(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_14),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_21),
.C(n_12),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_24),
.B(n_22),
.Y(n_25)
);

AOI322xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_8),
.A3(n_12),
.B1(n_7),
.B2(n_10),
.C1(n_3),
.C2(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_5),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_3),
.B(n_4),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_4),
.B(n_27),
.Y(n_29)
);


endmodule