module real_aes_6987_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_1), .A2(n_143), .B(n_155), .C(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g262 ( .A(n_2), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_3), .A2(n_170), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_4), .B(n_166), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g169 ( .A1(n_5), .A2(n_170), .B(n_171), .Y(n_169) );
AND2x6_ASAP7_75t_L g143 ( .A(n_6), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_7), .A2(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_8), .B(n_39), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g470 ( .A(n_9), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_10), .B(n_176), .Y(n_458) );
INVx1_ASAP7_75t_L g178 ( .A(n_11), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_12), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
INVx1_ASAP7_75t_L g244 ( .A(n_14), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_15), .A2(n_179), .B(n_245), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_16), .B(n_166), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_17), .B(n_189), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_18), .B(n_170), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_19), .B(n_512), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_20), .A2(n_146), .B(n_230), .C(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_21), .B(n_166), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_22), .B(n_176), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_23), .A2(n_242), .B(n_243), .C(n_245), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_24), .B(n_176), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_25), .Y(n_529) );
INVx1_ASAP7_75t_L g519 ( .A(n_26), .Y(n_519) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_28), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_29), .B(n_176), .Y(n_263) );
INVx1_ASAP7_75t_L g508 ( .A(n_30), .Y(n_508) );
INVx1_ASAP7_75t_L g154 ( .A(n_31), .Y(n_154) );
INVx2_ASAP7_75t_L g148 ( .A(n_32), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_33), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_34), .A2(n_180), .B(n_230), .C(n_497), .Y(n_496) );
INVxp67_ASAP7_75t_L g509 ( .A(n_35), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_36), .A2(n_143), .B(n_155), .C(n_200), .Y(n_199) );
CKINVDCx14_ASAP7_75t_R g495 ( .A(n_37), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_38), .A2(n_155), .B(n_518), .C(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g152 ( .A(n_40), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_41), .A2(n_175), .B(n_205), .C(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_42), .B(n_176), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_43), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_44), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_45), .Y(n_124) );
INVx1_ASAP7_75t_L g485 ( .A(n_46), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g158 ( .A(n_47), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_48), .B(n_170), .Y(n_232) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_49), .A2(n_58), .B1(n_126), .B2(n_712), .C1(n_713), .C2(n_717), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_50), .A2(n_146), .B1(n_149), .B2(n_155), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_51), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_52), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_53), .A2(n_175), .B(n_177), .C(n_180), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g467 ( .A(n_54), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_55), .Y(n_219) );
INVx1_ASAP7_75t_L g172 ( .A(n_56), .Y(n_172) );
INVx1_ASAP7_75t_L g144 ( .A(n_57), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_58), .Y(n_712) );
INVx1_ASAP7_75t_L g139 ( .A(n_59), .Y(n_139) );
INVx1_ASAP7_75t_SL g498 ( .A(n_60), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_62), .B(n_166), .Y(n_489) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_63), .A2(n_444), .B1(n_714), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_63), .Y(n_723) );
INVx1_ASAP7_75t_L g532 ( .A(n_64), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_SL g188 ( .A1(n_65), .A2(n_180), .B(n_189), .C(n_190), .Y(n_188) );
INVxp67_ASAP7_75t_L g191 ( .A(n_66), .Y(n_191) );
INVx1_ASAP7_75t_L g109 ( .A(n_67), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_68), .A2(n_170), .B(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_69), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_70), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_71), .A2(n_170), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g212 ( .A(n_72), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_73), .A2(n_238), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g477 ( .A(n_74), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_75), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_76), .A2(n_143), .B(n_155), .C(n_214), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_77), .A2(n_100), .B1(n_110), .B2(n_726), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_78), .A2(n_170), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g480 ( .A(n_79), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_80), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g456 ( .A(n_82), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_83), .B(n_189), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_84), .A2(n_143), .B(n_155), .C(n_261), .Y(n_260) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_85), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g120 ( .A(n_85), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g443 ( .A(n_85), .Y(n_443) );
OR2x2_ASAP7_75t_L g711 ( .A(n_85), .B(n_122), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_86), .A2(n_155), .B(n_531), .C(n_534), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_87), .B(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_88), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_89), .A2(n_143), .B(n_155), .C(n_227), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_90), .Y(n_234) );
INVx1_ASAP7_75t_L g187 ( .A(n_91), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_92), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_93), .B(n_202), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_94), .B(n_168), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_95), .B(n_168), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_96), .B(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_97), .A2(n_170), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g488 ( .A(n_98), .Y(n_488) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
CKINVDCx12_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g727 ( .A(n_103), .Y(n_727) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g122 ( .A(n_106), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_125), .B1(n_720), .B2(n_721), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_117), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g720 ( .A(n_114), .Y(n_720) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_117), .A2(n_722), .B(n_724), .Y(n_721) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_124), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g725 ( .A(n_120), .Y(n_725) );
NOR2x2_ASAP7_75t_L g719 ( .A(n_121), .B(n_443), .Y(n_719) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g442 ( .A(n_122), .B(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_440), .B1(n_444), .B2(n_711), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_128), .A2(n_440), .B1(n_714), .B2(n_715), .Y(n_713) );
AND3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_365), .C(n_414), .Y(n_128) );
NOR3xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_272), .C(n_310), .Y(n_129) );
OAI222xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_193), .B1(n_247), .B2(n_253), .C1(n_267), .C2(n_270), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_164), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_132), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_132), .B(n_315), .Y(n_406) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g283 ( .A(n_133), .B(n_184), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_133), .B(n_165), .Y(n_291) );
AND2x2_ASAP7_75t_L g326 ( .A(n_133), .B(n_303), .Y(n_326) );
OR2x2_ASAP7_75t_L g350 ( .A(n_133), .B(n_165), .Y(n_350) );
OR2x2_ASAP7_75t_L g358 ( .A(n_133), .B(n_257), .Y(n_358) );
AND2x2_ASAP7_75t_L g361 ( .A(n_133), .B(n_184), .Y(n_361) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g255 ( .A(n_134), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g269 ( .A(n_134), .B(n_184), .Y(n_269) );
AND2x2_ASAP7_75t_L g319 ( .A(n_134), .B(n_257), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_134), .B(n_165), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_134), .B(n_418), .Y(n_439) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_141), .B(n_162), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_135), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g207 ( .A(n_135), .Y(n_207) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_135), .A2(n_258), .B(n_265), .Y(n_257) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_137), .B(n_138), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI22xp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B1(n_158), .B2(n_159), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_172), .B(n_173), .C(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_142), .A2(n_173), .B(n_187), .C(n_188), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_142), .A2(n_173), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_142), .A2(n_173), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_142), .A2(n_173), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_142), .A2(n_173), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_142), .A2(n_173), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_142), .A2(n_173), .B(n_505), .C(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g534 ( .A(n_142), .Y(n_534) );
INVx4_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
NAND2x1p5_ASAP7_75t_L g159 ( .A(n_143), .B(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g170 ( .A(n_143), .B(n_160), .Y(n_170) );
BUFx3_ASAP7_75t_L g522 ( .A(n_143), .Y(n_522) );
INVx2_ASAP7_75t_L g264 ( .A(n_146), .Y(n_264) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
INVx1_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g149 ( .A1(n_150), .A2(n_152), .B1(n_153), .B2(n_154), .Y(n_149) );
INVx2_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
INVx4_ASAP7_75t_L g242 ( .A(n_150), .Y(n_242) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
AND2x2_ASAP7_75t_L g160 ( .A(n_151), .B(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
INVx3_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx1_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx2_ASAP7_75t_L g457 ( .A(n_153), .Y(n_457) );
INVx5_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
BUFx3_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_159), .A2(n_212), .B(n_213), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_159), .A2(n_259), .B(n_260), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_159), .A2(n_453), .B(n_454), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_159), .A2(n_183), .B(n_516), .C(n_517), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_159), .A2(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g510 ( .A(n_161), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_164), .A2(n_358), .B(n_359), .C(n_362), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_164), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_164), .B(n_302), .Y(n_424) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_184), .Y(n_164) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_165), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g282 ( .A(n_165), .Y(n_282) );
AND2x2_ASAP7_75t_L g309 ( .A(n_165), .B(n_303), .Y(n_309) );
INVx1_ASAP7_75t_SL g317 ( .A(n_165), .Y(n_317) );
AND2x2_ASAP7_75t_L g340 ( .A(n_165), .B(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g418 ( .A(n_165), .Y(n_418) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_182), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_SL g208 ( .A(n_167), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_167), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_167), .B(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_167), .A2(n_528), .B(n_535), .Y(n_527) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_168), .A2(n_185), .B(n_192), .Y(n_184) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_168), .Y(n_474) );
BUFx2_ASAP7_75t_L g238 ( .A(n_170), .Y(n_238) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g230 ( .A(n_176), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_179), .B(n_191), .Y(n_190) );
INVx5_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_179), .B(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_181), .Y(n_231) );
INVx1_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
INVx2_ASAP7_75t_L g224 ( .A(n_183), .Y(n_224) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_183), .A2(n_237), .B(n_246), .Y(n_236) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_183), .A2(n_465), .B(n_471), .Y(n_464) );
BUFx2_ASAP7_75t_L g254 ( .A(n_184), .Y(n_254) );
INVx1_ASAP7_75t_L g316 ( .A(n_184), .Y(n_316) );
INVx3_ASAP7_75t_L g341 ( .A(n_184), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_193), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_221), .Y(n_193) );
INVx1_ASAP7_75t_L g337 ( .A(n_194), .Y(n_337) );
OAI32xp33_ASAP7_75t_L g343 ( .A1(n_194), .A2(n_282), .A3(n_344), .B1(n_345), .B2(n_346), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_194), .A2(n_348), .B1(n_351), .B2(n_356), .Y(n_347) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g285 ( .A(n_195), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g363 ( .A(n_195), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g433 ( .A(n_195), .B(n_379), .Y(n_433) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
AND2x2_ASAP7_75t_L g248 ( .A(n_196), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g278 ( .A(n_196), .Y(n_278) );
INVx1_ASAP7_75t_L g297 ( .A(n_196), .Y(n_297) );
OR2x2_ASAP7_75t_L g305 ( .A(n_196), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g312 ( .A(n_196), .B(n_286), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_196), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_196), .B(n_251), .Y(n_333) );
INVx3_ASAP7_75t_L g355 ( .A(n_196), .Y(n_355) );
AND2x2_ASAP7_75t_L g380 ( .A(n_196), .B(n_252), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_196), .B(n_345), .Y(n_428) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_208), .Y(n_196) );
AOI21xp5_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_203), .B(n_204), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_202), .A2(n_262), .B(n_263), .C(n_264), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_202), .A2(n_242), .B1(n_508), .B2(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_202), .A2(n_519), .B(n_520), .C(n_521), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_204), .A2(n_215), .B(n_216), .Y(n_214) );
O2A1O1Ixp5_ASAP7_75t_L g455 ( .A1(n_204), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_204), .A2(n_457), .B(n_532), .C(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
INVx1_ASAP7_75t_L g217 ( .A(n_207), .Y(n_217) );
INVx2_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
AND2x2_ASAP7_75t_L g384 ( .A(n_210), .B(n_222), .Y(n_384) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_210) );
INVx1_ASAP7_75t_L g502 ( .A(n_217), .Y(n_502) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_217), .A2(n_555), .B(n_556), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_220), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_220), .B(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_220), .A2(n_452), .B(n_459), .Y(n_451) );
INVx2_ASAP7_75t_L g426 ( .A(n_221), .Y(n_426) );
OR2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_235), .Y(n_221) );
INVx1_ASAP7_75t_L g271 ( .A(n_222), .Y(n_271) );
AND2x2_ASAP7_75t_L g298 ( .A(n_222), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_222), .B(n_252), .Y(n_306) );
AND2x2_ASAP7_75t_L g364 ( .A(n_222), .B(n_287), .Y(n_364) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
AND2x2_ASAP7_75t_L g277 ( .A(n_223), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_223), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_223), .B(n_252), .Y(n_352) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_223) );
INVx1_ASAP7_75t_L g512 ( .A(n_224), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_224), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_231), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_230), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_235), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g299 ( .A(n_235), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_235), .B(n_252), .Y(n_345) );
AND2x2_ASAP7_75t_L g354 ( .A(n_235), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g379 ( .A(n_235), .Y(n_379) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g251 ( .A(n_236), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g287 ( .A(n_236), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_242), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_242), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_242), .B(n_488), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_247), .A2(n_257), .B1(n_416), .B2(n_419), .Y(n_415) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_249), .A2(n_360), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_250), .B(n_355), .Y(n_372) );
INVx1_ASAP7_75t_L g397 ( .A(n_250), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_251), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g324 ( .A(n_251), .B(n_277), .Y(n_324) );
INVx2_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
INVx1_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_253), .A2(n_405), .B1(n_422), .B2(n_425), .C(n_427), .Y(n_421) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_254), .B(n_303), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_255), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g346 ( .A(n_255), .B(n_292), .Y(n_346) );
INVx3_ASAP7_75t_SL g387 ( .A(n_255), .Y(n_387) );
AND2x2_ASAP7_75t_L g331 ( .A(n_256), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g360 ( .A(n_256), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_256), .B(n_269), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_256), .B(n_315), .Y(n_401) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx3_ASAP7_75t_L g303 ( .A(n_257), .Y(n_303) );
OAI322xp33_ASAP7_75t_L g398 ( .A1(n_257), .A2(n_329), .A3(n_351), .B1(n_399), .B2(n_401), .C1(n_402), .C2(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_268), .A2(n_271), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_269), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g370 ( .A(n_269), .B(n_282), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_269), .B(n_309), .Y(n_385) );
INVxp67_ASAP7_75t_L g336 ( .A(n_271), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g342 ( .A1(n_271), .A2(n_343), .B(n_347), .C(n_357), .Y(n_342) );
OAI221xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_281), .B1(n_284), .B2(n_288), .C(n_293), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g296 ( .A(n_280), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g413 ( .A(n_280), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_281), .A2(n_430), .B1(n_435), .B2(n_436), .C(n_438), .Y(n_429) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_282), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g329 ( .A(n_282), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_282), .B(n_360), .Y(n_367) );
AND2x2_ASAP7_75t_L g409 ( .A(n_282), .B(n_387), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_283), .B(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_283), .A2(n_295), .B1(n_405), .B2(n_406), .Y(n_404) );
OR2x2_ASAP7_75t_L g435 ( .A(n_283), .B(n_303), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g412 ( .A(n_286), .Y(n_412) );
AND2x2_ASAP7_75t_L g437 ( .A(n_286), .B(n_380), .Y(n_437) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g301 ( .A(n_291), .B(n_302), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_300), .B1(n_304), .B2(n_307), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g368 ( .A(n_296), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_296), .B(n_336), .Y(n_403) );
AOI322xp5_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_328), .A3(n_330), .B1(n_331), .B2(n_333), .C1(n_334), .C2(n_338), .Y(n_327) );
INVxp67_ASAP7_75t_L g321 ( .A(n_299), .Y(n_321) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_301), .A2(n_306), .B1(n_323), .B2(n_325), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_302), .B(n_315), .Y(n_402) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_303), .B(n_341), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_303), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g399 ( .A(n_305), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NAND3xp33_ASAP7_75t_SL g310 ( .A(n_311), .B(n_327), .C(n_342), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_318), .B2(n_320), .C(n_322), .Y(n_311) );
AND2x2_ASAP7_75t_L g318 ( .A(n_314), .B(n_319), .Y(n_318) );
INVx3_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g328 ( .A(n_319), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_321), .Y(n_400) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_326), .B(n_340), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_329), .B(n_387), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_330), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g405 ( .A(n_333), .Y(n_405) );
AND2x2_ASAP7_75t_L g420 ( .A(n_333), .B(n_397), .Y(n_420) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_344), .A2(n_415), .B(n_421), .C(n_429), .Y(n_414) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g383 ( .A(n_354), .B(n_384), .Y(n_383) );
NAND2x1_ASAP7_75t_SL g425 ( .A(n_355), .B(n_426), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g395 ( .A(n_358), .Y(n_395) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
AND2x2_ASAP7_75t_L g394 ( .A(n_364), .B(n_380), .Y(n_394) );
NOR5xp2_ASAP7_75t_L g365 ( .A(n_366), .B(n_381), .C(n_398), .D(n_404), .E(n_407), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_369), .B2(n_371), .C(n_373), .Y(n_366) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_370), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g396 ( .A(n_380), .B(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_385), .B1(n_386), .B2(n_388), .C(n_391), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
AOI211xp5_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_410), .B(n_412), .C(n_413), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
CKINVDCx14_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g714 ( .A(n_444), .Y(n_714) );
OR2x2_ASAP7_75t_SL g444 ( .A(n_445), .B(n_666), .Y(n_444) );
NAND5xp2_ASAP7_75t_L g445 ( .A(n_446), .B(n_578), .C(n_616), .D(n_637), .E(n_654), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_550), .C(n_571), .Y(n_446) );
OAI221xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_490), .B1(n_513), .B2(n_537), .C(n_541), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_461), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_450), .B(n_539), .Y(n_558) );
OR2x2_ASAP7_75t_L g585 ( .A(n_450), .B(n_473), .Y(n_585) );
AND2x2_ASAP7_75t_L g599 ( .A(n_450), .B(n_473), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_450), .B(n_464), .Y(n_613) );
AND2x2_ASAP7_75t_L g651 ( .A(n_450), .B(n_615), .Y(n_651) );
AND2x2_ASAP7_75t_L g680 ( .A(n_450), .B(n_590), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_450), .B(n_562), .Y(n_697) );
INVx4_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g577 ( .A(n_451), .B(n_472), .Y(n_577) );
BUFx3_ASAP7_75t_L g602 ( .A(n_451), .Y(n_602) );
AND2x2_ASAP7_75t_L g631 ( .A(n_451), .B(n_473), .Y(n_631) );
AND3x2_ASAP7_75t_L g644 ( .A(n_451), .B(n_645), .C(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g567 ( .A(n_461), .Y(n_567) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
AOI32xp33_ASAP7_75t_L g622 ( .A1(n_462), .A2(n_574), .A3(n_623), .B1(n_626), .B2(n_627), .Y(n_622) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g549 ( .A(n_463), .B(n_472), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_463), .B(n_577), .Y(n_620) );
AND2x2_ASAP7_75t_L g627 ( .A(n_463), .B(n_599), .Y(n_627) );
OR2x2_ASAP7_75t_L g633 ( .A(n_463), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_463), .B(n_588), .Y(n_658) );
OR2x2_ASAP7_75t_L g676 ( .A(n_463), .B(n_501), .Y(n_676) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g540 ( .A(n_464), .B(n_482), .Y(n_540) );
INVx2_ASAP7_75t_L g562 ( .A(n_464), .Y(n_562) );
OR2x2_ASAP7_75t_L g584 ( .A(n_464), .B(n_482), .Y(n_584) );
AND2x2_ASAP7_75t_L g589 ( .A(n_464), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_464), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g645 ( .A(n_464), .B(n_539), .Y(n_645) );
INVx1_ASAP7_75t_SL g696 ( .A(n_472), .Y(n_696) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
INVx1_ASAP7_75t_SL g539 ( .A(n_473), .Y(n_539) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_473), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_473), .B(n_625), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_473), .B(n_562), .C(n_680), .Y(n_691) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_474), .A2(n_483), .B(n_489), .Y(n_482) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_474), .A2(n_493), .B(n_499), .Y(n_492) );
INVx2_ASAP7_75t_L g590 ( .A(n_482), .Y(n_590) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_482), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_500), .Y(n_490) );
INVx1_ASAP7_75t_L g626 ( .A(n_491), .Y(n_626) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g544 ( .A(n_492), .B(n_526), .Y(n_544) );
INVx2_ASAP7_75t_L g561 ( .A(n_492), .Y(n_561) );
AND2x2_ASAP7_75t_L g566 ( .A(n_492), .B(n_527), .Y(n_566) );
AND2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_514), .Y(n_581) );
AND2x2_ASAP7_75t_L g593 ( .A(n_492), .B(n_565), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_500), .B(n_609), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_500), .B(n_566), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_500), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_500), .B(n_560), .Y(n_688) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g525 ( .A(n_501), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_501), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g570 ( .A(n_501), .B(n_514), .Y(n_570) );
AND2x2_ASAP7_75t_L g596 ( .A(n_501), .B(n_526), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_501), .B(n_636), .Y(n_635) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_511), .Y(n_501) );
INVx1_ASAP7_75t_L g555 ( .A(n_503), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_510), .Y(n_506) );
INVx2_ASAP7_75t_L g521 ( .A(n_510), .Y(n_521) );
INVx1_ASAP7_75t_L g556 ( .A(n_511), .Y(n_556) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_525), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_514), .B(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g560 ( .A(n_514), .B(n_561), .Y(n_560) );
INVx3_ASAP7_75t_SL g565 ( .A(n_514), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_514), .B(n_552), .Y(n_618) );
OR2x2_ASAP7_75t_L g628 ( .A(n_514), .B(n_554), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_514), .B(n_596), .Y(n_656) );
OR2x2_ASAP7_75t_L g686 ( .A(n_514), .B(n_526), .Y(n_686) );
AND2x2_ASAP7_75t_L g690 ( .A(n_514), .B(n_527), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_514), .B(n_566), .Y(n_703) );
AND2x2_ASAP7_75t_L g710 ( .A(n_514), .B(n_592), .Y(n_710) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
INVx1_ASAP7_75t_SL g653 ( .A(n_525), .Y(n_653) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_554), .Y(n_592) );
AND2x2_ASAP7_75t_L g606 ( .A(n_526), .B(n_561), .Y(n_606) );
AND2x2_ASAP7_75t_L g609 ( .A(n_526), .B(n_565), .Y(n_609) );
INVx1_ASAP7_75t_L g636 ( .A(n_526), .Y(n_636) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g548 ( .A(n_527), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_538), .A2(n_584), .B(n_708), .C(n_709), .Y(n_707) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g614 ( .A(n_539), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_540), .B(n_557), .Y(n_572) );
AND2x2_ASAP7_75t_L g598 ( .A(n_540), .B(n_599), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_545), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_543), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g569 ( .A(n_544), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_544), .B(n_565), .Y(n_610) );
AND2x2_ASAP7_75t_L g701 ( .A(n_544), .B(n_552), .Y(n_701) );
INVxp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g574 ( .A(n_548), .B(n_561), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_548), .B(n_559), .Y(n_575) );
OAI322xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_558), .A3(n_559), .B1(n_562), .B2(n_563), .C1(n_567), .C2(n_568), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_557), .Y(n_551) );
AND2x2_ASAP7_75t_L g662 ( .A(n_552), .B(n_574), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_552), .B(n_626), .Y(n_708) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g605 ( .A(n_554), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g671 ( .A(n_558), .B(n_584), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_559), .B(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_560), .B(n_592), .Y(n_649) );
AND2x2_ASAP7_75t_L g595 ( .A(n_561), .B(n_565), .Y(n_595) );
AND2x2_ASAP7_75t_L g603 ( .A(n_562), .B(n_604), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g700 ( .A1(n_562), .A2(n_641), .B(n_701), .C(n_702), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_563), .A2(n_576), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_565), .B(n_592), .Y(n_632) );
AND2x2_ASAP7_75t_L g638 ( .A(n_565), .B(n_606), .Y(n_638) );
AND2x2_ASAP7_75t_L g672 ( .A(n_565), .B(n_574), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_566), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g682 ( .A(n_566), .Y(n_682) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_570), .A2(n_598), .B1(n_600), .B2(n_605), .Y(n_597) );
OAI22xp5_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_573), .B1(n_575), .B2(n_576), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_572), .A2(n_608), .B1(n_610), .B2(n_611), .Y(n_607) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_577), .A2(n_679), .B1(n_681), .B2(n_683), .C(n_687), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B(n_586), .C(n_607), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OR2x2_ASAP7_75t_L g648 ( .A(n_584), .B(n_601), .Y(n_648) );
INVx1_ASAP7_75t_L g699 ( .A(n_584), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_585), .A2(n_587), .B1(n_591), .B2(n_594), .C(n_597), .Y(n_586) );
INVx2_ASAP7_75t_SL g641 ( .A(n_585), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g706 ( .A(n_588), .Y(n_706) );
AND2x2_ASAP7_75t_L g630 ( .A(n_589), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g615 ( .A(n_590), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g677 ( .A(n_593), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_601), .B(n_703), .Y(n_702) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_L g646 ( .A(n_604), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_605), .A2(n_617), .B(n_619), .C(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g694 ( .A(n_608), .Y(n_694) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_612), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx2_ASAP7_75t_L g625 ( .A(n_615), .Y(n_625) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_628), .B1(n_629), .B2(n_632), .C1(n_633), .C2(n_635), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g661 ( .A(n_625), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_628), .B(n_682), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_629), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g634 ( .A(n_631), .Y(n_634) );
AND2x2_ASAP7_75t_L g698 ( .A(n_631), .B(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g664 ( .A(n_634), .B(n_661), .Y(n_664) );
INVx1_ASAP7_75t_L g693 ( .A(n_635), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_642), .C(n_647), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_641), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_644), .A2(n_672), .A3(n_677), .B1(n_693), .B2(n_694), .C1(n_695), .C2(n_698), .Y(n_692) );
AND2x2_ASAP7_75t_L g679 ( .A(n_645), .B(n_680), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_650), .B2(n_652), .Y(n_647) );
INVxp33_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B1(n_659), .B2(n_662), .C(n_663), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND5xp2_ASAP7_75t_L g666 ( .A(n_667), .B(n_678), .C(n_692), .D(n_700), .E(n_704), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_672), .B(n_673), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVxp33_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_680), .A2(n_705), .B(n_706), .C(n_707), .Y(n_704) );
AOI31xp33_ASAP7_75t_L g687 ( .A1(n_682), .A2(n_688), .A3(n_689), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g705 ( .A(n_703), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_711), .Y(n_716) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
endmodule