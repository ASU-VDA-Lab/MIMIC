module real_jpeg_12014_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_3),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_40),
.B1(n_46),
.B2(n_50),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_33),
.B1(n_37),
.B2(n_135),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_135),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_46),
.B1(n_50),
.B2(n_135),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_6),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_6),
.A2(n_33),
.B1(n_37),
.B2(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_174),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_6),
.A2(n_46),
.B1(n_50),
.B2(n_174),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_8),
.A2(n_46),
.B1(n_50),
.B2(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_33),
.B1(n_37),
.B2(n_57),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_33),
.B1(n_37),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_46),
.B1(n_50),
.B2(n_69),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_30),
.B1(n_53),
.B2(n_54),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_30),
.B1(n_46),
.B2(n_50),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_12),
.A2(n_33),
.B1(n_37),
.B2(n_159),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_159),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_46),
.B1(n_50),
.B2(n_159),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_13),
.A2(n_33),
.B1(n_37),
.B2(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_93),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_13),
.A2(n_46),
.B1(n_50),
.B2(n_93),
.Y(n_229)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_15),
.A2(n_27),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_15),
.B(n_196),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_172),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_15),
.A2(n_49),
.B(n_53),
.C(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_15),
.B(n_70),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_86),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_15),
.B(n_44),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_15),
.A2(n_37),
.B(n_62),
.C(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_16),
.A2(n_33),
.B1(n_37),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_16),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_61),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_16),
.A2(n_46),
.B1(n_50),
.B2(n_61),
.Y(n_150)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_94),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_22),
.B(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_72),
.C(n_79),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_23),
.A2(n_72),
.B1(n_73),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_24),
.A2(n_25),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_43),
.C(n_59),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_27),
.A2(n_33),
.A3(n_36),
.B1(n_171),
.B2(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_28),
.B(n_172),
.Y(n_171)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_31),
.A2(n_32),
.B1(n_39),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_31),
.A2(n_32),
.B1(n_92),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_31),
.A2(n_32),
.B1(n_134),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_31),
.A2(n_32),
.B1(n_169),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_32),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_33),
.B(n_172),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_35),
.B(n_37),
.Y(n_189)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_37),
.A2(n_54),
.A3(n_64),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_58),
.B1(n_59),
.B2(n_71),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_43),
.A2(n_71),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_51),
.B1(n_56),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_51),
.B1(n_78),
.B2(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_44),
.A2(n_51),
.B1(n_90),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_44),
.A2(n_51),
.B1(n_153),
.B2(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_44),
.A2(n_51),
.B1(n_180),
.B2(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_44),
.A2(n_51),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_44),
.A2(n_51),
.B1(n_241),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_45),
.A2(n_130),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_45),
.A2(n_154),
.B1(n_221),
.B2(n_279),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_46),
.B(n_264),
.Y(n_263)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_48),
.A2(n_50),
.B(n_172),
.Y(n_243)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_51),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_53),
.B(n_65),
.Y(n_227)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_67),
.B2(n_70),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_62),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_62),
.A2(n_70),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_62),
.A2(n_70),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_68),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_66),
.A2(n_76),
.B1(n_102),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_66),
.A2(n_102),
.B1(n_132),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_66),
.A2(n_102),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_66),
.A2(n_193),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_91),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_81),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_87),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_84),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_84),
.A2(n_86),
.B1(n_150),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_84),
.A2(n_86),
.B1(n_186),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_84),
.A2(n_86),
.B1(n_198),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_84),
.A2(n_86),
.B1(n_229),
.B2(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_84),
.A2(n_86),
.B1(n_172),
.B2(n_262),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_84),
.A2(n_86),
.B1(n_255),
.B2(n_262),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_126),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_85),
.A2(n_148),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_136),
.B(n_309),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_109),
.B(n_112),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_131),
.C(n_133),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_122),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_295)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_162),
.B(n_308),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_160),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_139),
.B(n_160),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_144),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_140),
.B(n_143),
.Y(n_306)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_144),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.C(n_157),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_145),
.A2(n_146),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_151),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_155),
.B(n_157),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_303),
.B(n_307),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_213),
.B(n_291),
.C(n_302),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_199),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_165),
.B(n_199),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_183),
.C(n_190),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_166),
.A2(n_167),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_176),
.C(n_182),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_190),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.C(n_197),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_205),
.B(n_208),
.C(n_212),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_290),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_233),
.B(n_289),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_230),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_216),
.B(n_230),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_222),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_283),
.B(n_288),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_271),
.B(n_282),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_251),
.B(n_270),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_237),
.B(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_247),
.C(n_249),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_250),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_259),
.B(n_269),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_257),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_265),
.B(n_268),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_266),
.B(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_301),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_300),
.C(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);


endmodule