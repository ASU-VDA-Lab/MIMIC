module fake_jpeg_2938_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_9),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_50),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_32),
.B(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_44),
.B1(n_37),
.B2(n_46),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_53),
.B1(n_52),
.B2(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_36),
.B1(n_44),
.B2(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_1),
.B(n_2),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_69),
.B(n_4),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_2),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_26),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_74),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_96),
.C(n_84),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_5),
.B(n_6),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_3),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_30),
.C(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_3),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_24),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_79),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_84),
.B(n_25),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_112),
.B1(n_116),
.B2(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_114),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_23),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_115),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_8),
.C(n_11),
.Y(n_113)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_96),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_13),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_11),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_20),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_92),
.C(n_95),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_105),
.C(n_109),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_110),
.CI(n_115),
.CON(n_125),
.SN(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_121),
.C(n_122),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_131),
.B(n_132),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_129),
.C(n_128),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_127),
.B(n_125),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_129),
.B(n_125),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_120),
.B(n_18),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_16),
.CI(n_18),
.CON(n_137),
.SN(n_137)
);


endmodule