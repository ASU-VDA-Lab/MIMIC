module real_jpeg_16385_n_19 (n_17, n_8, n_0, n_141, n_2, n_132, n_139, n_142, n_10, n_137, n_9, n_12, n_135, n_134, n_6, n_136, n_133, n_11, n_14, n_131, n_138, n_7, n_18, n_3, n_5, n_4, n_1, n_140, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_141;
input n_2;
input n_132;
input n_139;
input n_142;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_134;
input n_6;
input n_136;
input n_133;
input n_11;
input n_14;
input n_131;
input n_138;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_140;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_3),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_4),
.B(n_76),
.C(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_6),
.B(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_7),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_72),
.C(n_96),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_74),
.B(n_85),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_13),
.B(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_14),
.Y(n_124)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_52),
.A3(n_64),
.B1(n_67),
.B2(n_105),
.C1(n_107),
.C2(n_142),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_17),
.Y(n_113)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_18),
.B(n_55),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_121),
.B(n_127),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_36),
.B(n_119),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_30),
.B(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_110),
.B(n_116),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI31xp67_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.A3(n_71),
.B(n_101),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_51),
.C(n_58),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_45),
.B(n_60),
.C(n_106),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_58),
.A3(n_102),
.B1(n_103),
.B2(n_104),
.C(n_141),
.Y(n_101)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_91),
.C(n_92),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_80),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_131),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_132),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_133),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_134),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_135),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_136),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_137),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_138),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_139),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_140),
.Y(n_97)
);


endmodule