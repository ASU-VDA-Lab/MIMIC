module fake_aes_8074_n_679 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_679);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_679;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_26), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_11), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_71), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_58), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_35), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_67), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_75), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_3), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_17), .B(n_64), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_13), .Y(n_92) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_48), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_72), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_54), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_29), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_56), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_25), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_24), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_42), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_53), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_37), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_55), .Y(n_105) );
BUFx2_ASAP7_75t_SL g106 ( .A(n_20), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_41), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_61), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_63), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_18), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_2), .Y(n_113) );
INVxp33_ASAP7_75t_L g114 ( .A(n_4), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_59), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_80), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_17), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_15), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_9), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_13), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_4), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_65), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_7), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_30), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
NOR2xp33_ASAP7_75t_R g132 ( .A(n_97), .B(n_36), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_125), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_125), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_92), .B(n_0), .Y(n_141) );
NOR2xp33_ASAP7_75t_R g142 ( .A(n_112), .B(n_38), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_112), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
NOR2xp33_ASAP7_75t_R g145 ( .A(n_89), .B(n_40), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_82), .B(n_1), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_93), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_90), .A2(n_94), .B(n_102), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_88), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_99), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_113), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_110), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_119), .B(n_1), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_106), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_92), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_106), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_123), .B(n_2), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_98), .B(n_5), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_98), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_120), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_101), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_102), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_101), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_117), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_109), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_117), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
BUFx4_ASAP7_75t_L g177 ( .A(n_166), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_150), .B(n_95), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_143), .B(n_100), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_161), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_139), .Y(n_185) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_137), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_137), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_133), .Y(n_191) );
INVxp67_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_172), .A2(n_129), .B1(n_122), .B2(n_107), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_164), .B(n_129), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_174), .B(n_130), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_164), .B(n_170), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_170), .B(n_122), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_159), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_153), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_158), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_155), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_131), .B(n_89), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_149), .B(n_81), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_163), .B(n_115), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_168), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_168), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_173), .Y(n_219) );
BUFx10_ASAP7_75t_L g220 ( .A(n_154), .Y(n_220) );
NAND3x1_ASAP7_75t_L g221 ( .A(n_157), .B(n_128), .C(n_118), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_156), .B(n_116), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_173), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_157), .B(n_127), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_173), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_131), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_134), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_134), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_135), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_135), .B(n_128), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_136), .B(n_83), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_136), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_138), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_138), .B(n_111), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_142), .Y(n_236) );
OR2x2_ASAP7_75t_SL g237 ( .A(n_146), .B(n_124), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_144), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_148), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_148), .A2(n_124), .B(n_121), .C(n_118), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_233), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_204), .B(n_175), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_179), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g245 ( .A(n_192), .B(n_213), .C(n_222), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_204), .B(n_171), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_196), .B(n_162), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
BUFx8_ASAP7_75t_SL g251 ( .A(n_208), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_178), .B(n_162), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_196), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_211), .B(n_160), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_233), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_215), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_220), .Y(n_257) );
INVx6_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
CKINVDCx11_ASAP7_75t_R g260 ( .A(n_220), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_180), .B(n_160), .Y(n_261) );
AND3x1_ASAP7_75t_L g262 ( .A(n_180), .B(n_152), .C(n_169), .Y(n_262) );
AO22x1_ASAP7_75t_L g263 ( .A1(n_176), .A2(n_105), .B1(n_103), .B2(n_121), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_181), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_184), .B(n_145), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
NOR2xp33_ASAP7_75t_R g267 ( .A(n_185), .B(n_104), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_214), .A2(n_167), .B1(n_132), .B2(n_8), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_220), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_184), .B(n_45), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_187), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
AOI22xp5_ASAP7_75t_SL g274 ( .A1(n_208), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_211), .B(n_6), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_186), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_214), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_195), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
OR2x2_ASAP7_75t_SL g280 ( .A(n_177), .B(n_9), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_181), .Y(n_281) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_214), .B(n_10), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_211), .B(n_10), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_233), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_181), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_182), .B(n_49), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_194), .A2(n_191), .B1(n_197), .B2(n_231), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_191), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_218), .Y(n_291) );
OR2x6_ASAP7_75t_L g292 ( .A(n_221), .B(n_14), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_187), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_188), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_207), .Y(n_295) );
AOI22x1_ASAP7_75t_L g296 ( .A1(n_213), .A2(n_50), .B1(n_77), .B2(n_74), .Y(n_296) );
NOR2xp33_ASAP7_75t_R g297 ( .A(n_210), .B(n_46), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_188), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_221), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_210), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_224), .Y(n_301) );
INVx5_ASAP7_75t_L g302 ( .A(n_197), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_225), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_197), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_225), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_236), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_189), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_189), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_258), .Y(n_309) );
BUFx5_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_273), .B(n_278), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_249), .B(n_206), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_258), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_243), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_246), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_243), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_248), .B(n_230), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_247), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_248), .B(n_230), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_244), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_273), .B(n_212), .Y(n_326) );
OR2x2_ASAP7_75t_SL g327 ( .A(n_272), .B(n_177), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_261), .B(n_228), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_261), .B(n_228), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_278), .B(n_198), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_244), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_253), .B(n_238), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_246), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_244), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_266), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_260), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_304), .A2(n_205), .B(n_207), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_292), .B(n_213), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_253), .Y(n_339) );
BUFx12f_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_292), .A2(n_226), .B1(n_239), .B2(n_229), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_246), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_252), .B(n_239), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_242), .A2(n_205), .B(n_226), .Y(n_344) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_245), .B(n_240), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_276), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_282), .B(n_234), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_256), .B(n_223), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_301), .B(n_238), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_254), .B(n_235), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_257), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_256), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_266), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_244), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_256), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_244), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_264), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_271), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_264), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_263), .B(n_235), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_310), .B(n_269), .Y(n_362) );
AND2x6_ASAP7_75t_L g363 ( .A(n_319), .B(n_284), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_289), .B1(n_262), .B2(n_299), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
OAI222xp33_ASAP7_75t_L g366 ( .A1(n_338), .A2(n_274), .B1(n_300), .B2(n_269), .C1(n_290), .C2(n_268), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_312), .B(n_301), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_308), .B(n_307), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_312), .B(n_277), .Y(n_370) );
BUFx4f_ASAP7_75t_SL g371 ( .A(n_340), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_349), .B(n_271), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_346), .B(n_290), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_300), .B1(n_306), .B2(n_275), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_319), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_340), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_337), .A2(n_281), .B(n_264), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_341), .A2(n_307), .B1(n_293), .B2(n_298), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_316), .A2(n_283), .B1(n_306), .B2(n_284), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_358), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_316), .A2(n_265), .B(n_259), .Y(n_383) );
AND2x4_ASAP7_75t_SL g384 ( .A(n_338), .B(n_293), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_348), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_320), .B(n_263), .Y(n_386) );
HB1xp67_ASAP7_75t_SL g387 ( .A(n_336), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_321), .A2(n_325), .B1(n_347), .B2(n_338), .Y(n_388) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_321), .A2(n_280), .B1(n_296), .B2(n_298), .C1(n_294), .C2(n_270), .Y(n_389) );
NAND2xp33_ASAP7_75t_R g390 ( .A(n_351), .B(n_267), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_349), .B(n_294), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_361), .A2(n_259), .B(n_295), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
INVx4_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_347), .B1(n_251), .B2(n_326), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_394), .B(n_335), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_394), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_367), .A2(n_323), .B1(n_329), .B2(n_328), .C(n_347), .Y(n_398) );
AOI21x1_ASAP7_75t_L g399 ( .A1(n_377), .A2(n_360), .B(n_334), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_360), .B(n_356), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_370), .B(n_347), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_375), .B(n_327), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_372), .B(n_353), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_326), .B1(n_330), .B2(n_343), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_373), .A2(n_326), .B1(n_330), .B2(n_311), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_373), .A2(n_326), .B1(n_330), .B2(n_311), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_330), .B1(n_311), .B2(n_359), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_372), .B(n_353), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_394), .A2(n_327), .B1(n_280), .B2(n_359), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_380), .B(n_339), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_380), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_391), .B(n_332), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_311), .B1(n_345), .B2(n_332), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_350), .B(n_348), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_342), .B1(n_333), .B2(n_352), .Y(n_420) );
OR2x6_ASAP7_75t_L g421 ( .A(n_385), .B(n_324), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_391), .B(n_288), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_371), .A2(n_342), .B1(n_333), .B2(n_352), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_422), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_402), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_411), .A2(n_381), .B1(n_388), .B2(n_379), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_403), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_395), .B(n_296), .C(n_383), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_398), .A2(n_369), .B1(n_365), .B2(n_384), .Y(n_430) );
NAND4xp25_ASAP7_75t_L g431 ( .A(n_406), .B(n_366), .C(n_365), .D(n_369), .Y(n_431) );
INVx4_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
NOR2xp33_ASAP7_75t_R g433 ( .A(n_417), .B(n_376), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g434 ( .A(n_407), .B(n_190), .C(n_193), .D(n_200), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_415), .B(n_382), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_409), .A2(n_368), .B1(n_393), .B2(n_382), .C(n_385), .Y(n_436) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_401), .A2(n_382), .B1(n_362), .B2(n_342), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_399), .A2(n_400), .B(n_418), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_396), .A2(n_384), .B1(n_363), .B2(n_297), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_396), .A2(n_384), .B1(n_363), .B2(n_392), .Y(n_441) );
AND2x6_ASAP7_75t_L g442 ( .A(n_397), .B(n_363), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_397), .B(n_310), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_410), .B(n_16), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_412), .A2(n_342), .B1(n_389), .B2(n_318), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_412), .B(n_237), .Y(n_447) );
OAI21x1_ASAP7_75t_L g448 ( .A1(n_399), .A2(n_360), .B(n_356), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_408), .A2(n_314), .B1(n_309), .B2(n_313), .C(n_317), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_416), .A2(n_314), .B1(n_309), .B2(n_313), .C(n_317), .Y(n_450) );
AOI31xp33_ASAP7_75t_L g451 ( .A1(n_396), .A2(n_387), .A3(n_223), .B(n_217), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_419), .B(n_237), .Y(n_452) );
NOR3xp33_ASAP7_75t_SL g453 ( .A(n_423), .B(n_287), .C(n_217), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_404), .B(n_219), .C(n_190), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_419), .B(n_313), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_396), .A2(n_363), .B1(n_310), .B2(n_318), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_404), .A2(n_324), .B1(n_357), .B2(n_331), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_427), .B(n_422), .C(n_419), .D(n_209), .Y(n_458) );
AOI33xp33_ASAP7_75t_L g459 ( .A1(n_444), .A2(n_420), .A3(n_216), .B1(n_405), .B2(n_414), .B3(n_413), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_428), .B(n_414), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_433), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_432), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_431), .A2(n_397), .B1(n_363), .B2(n_405), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_430), .B(n_413), .C(n_227), .D(n_232), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_439), .B(n_397), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_445), .B(n_421), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_442), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_448), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_425), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_424), .A2(n_363), .B1(n_421), .B2(n_313), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_426), .B(n_421), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_451), .B(n_18), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_442), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_442), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_436), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_440), .A2(n_421), .B1(n_352), .B2(n_318), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_452), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_447), .B(n_400), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_457), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_434), .B(n_19), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_455), .B(n_19), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_442), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_454), .B(n_291), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_441), .B(n_291), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_456), .B(n_288), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_429), .B(n_317), .C(n_227), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_443), .B(n_303), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_449), .B(n_305), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_453), .B(n_305), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_437), .B(n_21), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_425), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_431), .A2(n_232), .B1(n_201), .B2(n_203), .C(n_202), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_424), .Y(n_503) );
INVx6_ASAP7_75t_L g504 ( .A(n_432), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_428), .B(n_23), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_428), .B(n_355), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_484), .B(n_28), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_503), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_476), .B(n_183), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_484), .B(n_31), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_476), .B(n_355), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_501), .B(n_183), .Y(n_512) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_458), .B(n_355), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_471), .B(n_355), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_468), .Y(n_515) );
NOR3xp33_ASAP7_75t_SL g516 ( .A(n_461), .B(n_32), .C(n_34), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_500), .B(n_183), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_500), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_465), .B(n_44), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_465), .B(n_47), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_466), .B(n_51), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_466), .B(n_181), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_474), .B(n_52), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_483), .B(n_183), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_473), .B(n_57), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_493), .B(n_60), .Y(n_528) );
NAND2xp33_ASAP7_75t_R g529 ( .A(n_486), .B(n_62), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_486), .B(n_66), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_478), .B(n_68), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_493), .B(n_69), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_468), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_477), .B(n_70), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_481), .B(n_73), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_504), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_477), .B(n_78), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_504), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_480), .B(n_183), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_481), .B(n_354), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_504), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_504), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_485), .B(n_354), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_467), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_479), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_480), .B(n_310), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_469), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_459), .B(n_310), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_470), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_491), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_485), .B(n_354), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_488), .B(n_334), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_488), .B(n_334), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_470), .Y(n_556) );
NOR3xp33_ASAP7_75t_L g557 ( .A(n_487), .B(n_259), .C(n_250), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_489), .B(n_356), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_491), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_489), .B(n_241), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_513), .A2(n_496), .B1(n_464), .B2(n_498), .Y(n_561) );
INVxp33_ASAP7_75t_L g562 ( .A(n_541), .Y(n_562) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_508), .Y(n_563) );
A2O1A1O1Ixp25_ASAP7_75t_L g564 ( .A1(n_524), .A2(n_482), .B(n_463), .C(n_467), .D(n_475), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_526), .A2(n_499), .B(n_498), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_522), .B(n_505), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_518), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_515), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_557), .A2(n_494), .B1(n_505), .B2(n_499), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_543), .A2(n_472), .B1(n_502), .B2(n_492), .C(n_495), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_545), .B(n_475), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_545), .B(n_475), .Y(n_573) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_529), .A2(n_497), .B(n_495), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_515), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_533), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_552), .B(n_497), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_514), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_533), .Y(n_579) );
OAI311xp33_ASAP7_75t_L g580 ( .A1(n_528), .A2(n_490), .A3(n_302), .B1(n_310), .C1(n_264), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_530), .A2(n_310), .B1(n_302), .B2(n_286), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_546), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_559), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_511), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_524), .A2(n_241), .A3(n_250), .B(n_255), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_510), .B(n_357), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_536), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_538), .B(n_302), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_542), .Y(n_589) );
INVxp67_ASAP7_75t_SL g590 ( .A(n_546), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_507), .B(n_302), .Y(n_591) );
XNOR2x1_ASAP7_75t_L g592 ( .A(n_521), .B(n_255), .Y(n_592) );
OAI222xp33_ASAP7_75t_L g593 ( .A1(n_510), .A2(n_302), .B1(n_279), .B2(n_285), .C1(n_331), .C2(n_324), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_517), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_528), .B(n_357), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_550), .A2(n_264), .B1(n_281), .B2(n_286), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_532), .A2(n_324), .B(n_331), .Y(n_597) );
OAI322xp33_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_279), .A3(n_285), .B1(n_281), .B2(n_286), .C1(n_324), .C2(n_331), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_516), .A2(n_331), .B(n_281), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_532), .B(n_281), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_507), .A2(n_286), .B1(n_547), .B2(n_548), .C(n_535), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_540), .B(n_544), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_509), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_527), .B(n_521), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_549), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_563), .B(n_523), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_561), .B(n_527), .C(n_537), .D(n_534), .Y(n_607) );
XNOR2xp5_ASAP7_75t_L g608 ( .A(n_592), .B(n_519), .Y(n_608) );
OAI21xp33_ASAP7_75t_SL g609 ( .A1(n_567), .A2(n_535), .B(n_519), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_569), .B(n_551), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_569), .B(n_551), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_583), .B(n_553), .Y(n_612) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_572), .B(n_520), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_602), .B(n_553), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_575), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_574), .B(n_531), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_568), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_584), .B(n_544), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_572), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_578), .B(n_554), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_587), .Y(n_621) );
NAND2xp33_ASAP7_75t_R g622 ( .A(n_604), .B(n_555), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_589), .B(n_539), .Y(n_623) );
NOR2x1_ASAP7_75t_L g624 ( .A(n_573), .B(n_512), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_594), .B(n_556), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_566), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_570), .A2(n_558), .B1(n_556), .B2(n_560), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_590), .B(n_560), .Y(n_628) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_593), .B(n_558), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_590), .B(n_605), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_603), .B(n_577), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_579), .B(n_582), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_565), .B(n_605), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_581), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_621), .B(n_562), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_607), .B(n_588), .C(n_571), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_619), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_609), .A2(n_570), .B(n_601), .Y(n_639) );
AND3x2_ASAP7_75t_L g640 ( .A(n_629), .B(n_585), .C(n_564), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_627), .B(n_597), .C(n_591), .D(n_595), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_631), .B(n_576), .Y(n_642) );
NAND4xp25_ASAP7_75t_L g643 ( .A(n_616), .B(n_595), .C(n_596), .D(n_600), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_624), .B(n_596), .Y(n_644) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_626), .B(n_580), .C(n_586), .D(n_599), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_614), .B(n_600), .Y(n_646) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_630), .Y(n_647) );
OA21x2_ASAP7_75t_L g648 ( .A1(n_633), .A2(n_598), .B(n_632), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_608), .B(n_634), .Y(n_649) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_613), .B(n_622), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_639), .A2(n_617), .B1(n_623), .B2(n_616), .C(n_612), .Y(n_651) );
AOI31xp33_ASAP7_75t_L g652 ( .A1(n_649), .A2(n_622), .A3(n_606), .B(n_628), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_640), .A2(n_623), .B(n_610), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_638), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_650), .B(n_615), .Y(n_655) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_644), .B(n_611), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_647), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_637), .B(n_611), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_640), .A2(n_620), .B(n_618), .Y(n_659) );
NOR2xp33_ASAP7_75t_R g660 ( .A(n_645), .B(n_625), .Y(n_660) );
OAI22xp5_ASAP7_75t_SL g661 ( .A1(n_648), .A2(n_635), .B1(n_636), .B2(n_646), .Y(n_661) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_641), .B(n_643), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_648), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_650), .A2(n_639), .B(n_644), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_642), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_654), .Y(n_666) );
NOR2xp67_ASAP7_75t_L g667 ( .A(n_653), .B(n_659), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_662), .B(n_658), .Y(n_668) );
NOR2x1p5_ASAP7_75t_L g669 ( .A(n_663), .B(n_661), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_651), .B(n_664), .Y(n_670) );
NOR2x1p5_ASAP7_75t_L g671 ( .A(n_668), .B(n_665), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_666), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_670), .Y(n_673) );
AOI22xp33_ASAP7_75t_R g674 ( .A1(n_672), .A2(n_660), .B1(n_657), .B2(n_669), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_671), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_675), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_674), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_667), .B1(n_673), .B2(n_655), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_673), .B1(n_676), .B2(n_652), .C(n_656), .Y(n_679) );
endmodule