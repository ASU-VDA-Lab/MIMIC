module fake_jpeg_2603_n_708 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_708);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_708;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_65),
.Y(n_212)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_70),
.A2(n_58),
.B1(n_56),
.B2(n_53),
.Y(n_168)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_76),
.B(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_18),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_80),
.Y(n_207)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_88),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx6p67_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_86),
.Y(n_231)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_87),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_89),
.B(n_94),
.Y(n_228)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_90),
.Y(n_177)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_27),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g144 ( 
.A(n_92),
.Y(n_144)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_93),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_37),
.B(n_17),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_37),
.B(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_96),
.B(n_118),
.Y(n_161)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_35),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_105),
.B(n_40),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_108),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_109),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_39),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_35),
.B(n_16),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_41),
.B(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_120),
.B(n_125),
.Y(n_185)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_49),
.B(n_14),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_59),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_47),
.Y(n_165)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_38),
.Y(n_128)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g129 ( 
.A(n_43),
.Y(n_129)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_13),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_130),
.B(n_133),
.Y(n_189)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_24),
.Y(n_132)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_51),
.B(n_13),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_134),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_93),
.C(n_108),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_159),
.B(n_160),
.C(n_170),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_34),
.C(n_29),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_165),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_85),
.A2(n_43),
.B1(n_48),
.B2(n_23),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_167),
.A2(n_196),
.B1(n_202),
.B2(n_214),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_168),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_29),
.C(n_26),
.Y(n_170)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_88),
.B(n_56),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_181),
.B(n_197),
.Y(n_278)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_64),
.Y(n_184)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_70),
.A2(n_85),
.B(n_114),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g254 ( 
.A(n_192),
.B(n_77),
.Y(n_254)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_65),
.A2(n_43),
.B1(n_48),
.B2(n_23),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_67),
.B(n_49),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_198),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_73),
.B(n_53),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_205),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_86),
.A2(n_48),
.B1(n_47),
.B2(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_100),
.B(n_48),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_99),
.B(n_54),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_124),
.B(n_33),
.C(n_54),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_210),
.B(n_68),
.C(n_11),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_213),
.B(n_11),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_91),
.A2(n_47),
.B1(n_40),
.B2(n_28),
.Y(n_214)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_71),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_127),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_131),
.A2(n_47),
.B1(n_79),
.B2(n_97),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_229),
.B1(n_132),
.B2(n_95),
.Y(n_238)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_92),
.A2(n_28),
.B1(n_26),
.B2(n_59),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_225),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_113),
.B(n_128),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_72),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_81),
.A2(n_59),
.B1(n_13),
.B2(n_11),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_232),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_135),
.A2(n_122),
.B1(n_112),
.B2(n_87),
.Y(n_233)
);

AO21x2_ASAP7_75t_L g325 ( 
.A1(n_233),
.A2(n_254),
.B(n_290),
.Y(n_325)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_234),
.Y(n_329)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_238),
.A2(n_300),
.B1(n_307),
.B2(n_312),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_143),
.B(n_109),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_241),
.B(n_248),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_153),
.A2(n_110),
.B1(n_83),
.B2(n_104),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_244),
.A2(n_256),
.B1(n_275),
.B2(n_276),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_247),
.B(n_295),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_155),
.B(n_0),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_255),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_194),
.A2(n_101),
.B1(n_98),
.B2(n_75),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_257),
.B(n_281),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_0),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_258),
.B(n_297),
.Y(n_353)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_139),
.Y(n_259)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_177),
.B(n_0),
.Y(n_260)
);

NAND2x1_ASAP7_75t_L g368 ( 
.A(n_260),
.B(n_187),
.Y(n_368)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_262),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_263),
.Y(n_373)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_141),
.Y(n_264)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_179),
.Y(n_268)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_268),
.Y(n_348)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_157),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_269),
.Y(n_370)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_156),
.Y(n_270)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_144),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_271),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_279),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_211),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_277),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_164),
.B(n_123),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_280),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_162),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_182),
.Y(n_282)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_156),
.Y(n_283)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_152),
.Y(n_285)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_285),
.Y(n_374)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_137),
.Y(n_287)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_169),
.Y(n_288)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_298),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_189),
.A2(n_185),
.B1(n_161),
.B2(n_167),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_166),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_291),
.B(n_301),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_292),
.A2(n_302),
.B1(n_229),
.B2(n_214),
.Y(n_322)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_145),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_154),
.B(n_3),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_158),
.B(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_221),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_223),
.B(n_123),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_216),
.C(n_218),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_196),
.A2(n_106),
.B1(n_6),
.B2(n_7),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_207),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_211),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_302)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_306),
.Y(n_362)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_201),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_230),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_308),
.B(n_309),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_146),
.B(n_6),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_149),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_315),
.Y(n_320)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_227),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_314),
.Y(n_377)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_136),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_6),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_8),
.Y(n_356)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_147),
.B(n_8),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_202),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_231),
.Y(n_369)
);

AO22x1_ASAP7_75t_SL g321 ( 
.A1(n_237),
.A2(n_218),
.B1(n_136),
.B2(n_144),
.Y(n_321)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_321),
.A2(n_215),
.B(n_217),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_322),
.A2(n_331),
.B1(n_349),
.B2(n_234),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_254),
.A2(n_169),
.B(n_216),
.C(n_212),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_327),
.A2(n_289),
.B(n_217),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_272),
.A2(n_142),
.B1(n_188),
.B2(n_200),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_339),
.C(n_344),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_253),
.B(n_172),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_304),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_343),
.B(n_352),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_253),
.B(n_151),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_232),
.B(n_187),
.C(n_138),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_378),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_241),
.A2(n_142),
.B1(n_188),
.B2(n_200),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_255),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_356),
.B(n_375),
.Y(n_423)
);

OAI32xp33_ASAP7_75t_L g358 ( 
.A1(n_240),
.A2(n_171),
.A3(n_212),
.B1(n_190),
.B2(n_140),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_361),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_248),
.B(n_297),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_279),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_365),
.B(n_284),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_140),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_379),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_280),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_369),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_242),
.A2(n_178),
.B(n_183),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_262),
.B(n_269),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_278),
.B(n_231),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_274),
.B(n_149),
.C(n_215),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_258),
.B(n_260),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_380),
.Y(n_381)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_325),
.A2(n_292),
.B1(n_271),
.B2(n_314),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_385),
.A2(n_331),
.B1(n_373),
.B2(n_327),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_386),
.A2(n_389),
.B(n_428),
.Y(n_441)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_388),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_373),
.A2(n_235),
.B1(n_299),
.B2(n_233),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_325),
.A2(n_280),
.B1(n_260),
.B2(n_183),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_390),
.A2(n_392),
.B1(n_395),
.B2(n_396),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_325),
.A2(n_151),
.B1(n_191),
.B2(n_145),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_334),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_393),
.B(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_325),
.A2(n_191),
.B1(n_171),
.B2(n_190),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_325),
.A2(n_286),
.B1(n_296),
.B2(n_287),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_259),
.B1(n_266),
.B2(n_311),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_397),
.A2(n_406),
.B1(n_416),
.B2(n_424),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_407),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_326),
.A2(n_174),
.B1(n_294),
.B2(n_268),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_326),
.A2(n_174),
.B1(n_282),
.B2(n_261),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_333),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_261),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_411),
.Y(n_434)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_322),
.A2(n_252),
.B1(n_293),
.B2(n_273),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_372),
.A2(n_252),
.B1(n_267),
.B2(n_265),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_409),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_363),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_413),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_264),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_353),
.B(n_249),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_418),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_330),
.A2(n_245),
.B1(n_277),
.B2(n_285),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_415),
.A2(n_421),
.B1(n_431),
.B2(n_364),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_344),
.A2(n_245),
.B1(n_250),
.B2(n_270),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_345),
.B(n_246),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_417),
.B(n_375),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_366),
.B(n_243),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_362),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_422),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_420),
.B(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_354),
.A2(n_283),
.B1(n_239),
.B2(n_251),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_339),
.A2(n_251),
.B1(n_243),
.B2(n_236),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_367),
.B1(n_318),
.B2(n_328),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_379),
.B(n_310),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_368),
.Y(n_457)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_430),
.A2(n_364),
.B1(n_329),
.B2(n_370),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_369),
.A2(n_305),
.B1(n_288),
.B2(n_312),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_432),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_436),
.A2(n_421),
.B(n_406),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_338),
.C(n_378),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_443),
.C(n_454),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_383),
.A2(n_323),
.B1(n_320),
.B2(n_321),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_439),
.A2(n_449),
.B1(n_451),
.B2(n_453),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_323),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_384),
.B(n_371),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_388),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_383),
.A2(n_320),
.B1(n_321),
.B2(n_358),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_393),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_356),
.B1(n_347),
.B2(n_377),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_368),
.C(n_328),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_426),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_457),
.Y(n_475)
);

OAI21xp33_ASAP7_75t_SL g501 ( 
.A1(n_456),
.A2(n_421),
.B(n_424),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_414),
.B(n_404),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_464),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_395),
.A2(n_349),
.B1(n_346),
.B2(n_317),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_461),
.A2(n_468),
.B1(n_472),
.B2(n_392),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_357),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_398),
.A2(n_359),
.B1(n_346),
.B2(n_351),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_402),
.B(n_324),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_427),
.C(n_416),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_402),
.B(n_374),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_388),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_396),
.A2(n_329),
.B1(n_374),
.B2(n_351),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_418),
.B(n_336),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_474),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_429),
.B(n_423),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_449),
.A2(n_439),
.B(n_456),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_512),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_441),
.A2(n_412),
.B(n_428),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_479),
.A2(n_494),
.B(n_497),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_462),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_480),
.B(n_500),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_510),
.Y(n_516)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_483),
.B(n_485),
.Y(n_525)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_486),
.Y(n_530)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_489),
.C(n_432),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_447),
.A2(n_423),
.B(n_388),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_460),
.Y(n_491)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_492),
.A2(n_498),
.B1(n_508),
.B2(n_461),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_441),
.A2(n_412),
.B(n_386),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_426),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_444),
.C(n_454),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_496),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_455),
.A2(n_410),
.B1(n_442),
.B2(n_459),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_460),
.Y(n_499)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_440),
.B1(n_446),
.B2(n_468),
.Y(n_515)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_502),
.Y(n_537)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_503),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_514),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_458),
.B(n_399),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_505),
.B(n_507),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_450),
.B(n_387),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_440),
.A2(n_390),
.B1(n_446),
.B2(n_442),
.Y(n_508)
);

OAI32xp33_ASAP7_75t_L g509 ( 
.A1(n_450),
.A2(n_382),
.A3(n_422),
.B1(n_394),
.B2(n_405),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_511),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_443),
.B(n_415),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_466),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_448),
.A2(n_421),
.B(n_413),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_513),
.A2(n_436),
.B(n_457),
.Y(n_518)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_467),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_515),
.A2(n_526),
.B1(n_529),
.B2(n_538),
.Y(n_554)
);

AND2x2_ASAP7_75t_SL g517 ( 
.A(n_475),
.B(n_448),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_517),
.B(n_543),
.Y(n_555)
);

AO21x1_ASAP7_75t_L g588 ( 
.A1(n_518),
.A2(n_523),
.B(n_539),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_524),
.C(n_533),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_496),
.B(n_469),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_522),
.B(n_551),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_474),
.B(n_434),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_478),
.B(n_471),
.C(n_453),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_495),
.B(n_470),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g581 ( 
.A(n_527),
.B(n_319),
.Y(n_581)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_506),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_528),
.B(n_542),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_478),
.B(n_434),
.C(n_464),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_476),
.A2(n_451),
.B1(n_447),
.B2(n_407),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_491),
.A2(n_499),
.B1(n_475),
.B2(n_484),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_473),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_511),
.Y(n_573)
);

NOR2x1_ASAP7_75t_L g542 ( 
.A(n_507),
.B(n_467),
.Y(n_542)
);

AOI32xp33_ASAP7_75t_L g543 ( 
.A1(n_479),
.A2(n_409),
.A3(n_381),
.B1(n_417),
.B2(n_438),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_510),
.B(n_400),
.C(n_355),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_548),
.B(n_550),
.C(n_527),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_508),
.A2(n_397),
.B1(n_472),
.B2(n_438),
.Y(n_549)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_485),
.B(n_337),
.C(n_355),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_500),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_476),
.Y(n_552)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_552),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_477),
.A2(n_431),
.B1(n_445),
.B2(n_403),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_553),
.A2(n_445),
.B1(n_403),
.B2(n_430),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_538),
.A2(n_477),
.B1(n_513),
.B2(n_493),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_556),
.A2(n_557),
.B1(n_558),
.B2(n_572),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_546),
.A2(n_493),
.B1(n_505),
.B2(n_490),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_546),
.A2(n_535),
.B1(n_515),
.B2(n_518),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_542),
.B(n_509),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_SL g603 ( 
.A(n_559),
.B(n_561),
.C(n_576),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_480),
.Y(n_560)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_560),
.Y(n_589)
);

XOR2x1_ASAP7_75t_SL g561 ( 
.A(n_535),
.B(n_497),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_521),
.A2(n_484),
.B(n_490),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_563),
.A2(n_569),
.B(n_532),
.Y(n_594)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_536),
.Y(n_564)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_564),
.Y(n_592)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_537),
.Y(n_565)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_537),
.Y(n_567)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_521),
.A2(n_514),
.B(n_512),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_547),
.Y(n_570)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_570),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_517),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_571),
.B(n_587),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_535),
.A2(n_492),
.B1(n_481),
.B2(n_503),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_573),
.B(n_575),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_502),
.B1(n_487),
.B2(n_486),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_574),
.A2(n_583),
.B1(n_531),
.B2(n_530),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_547),
.B(n_482),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_337),
.C(n_336),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_577),
.B(n_540),
.C(n_550),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_324),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_581),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_534),
.B(n_504),
.Y(n_580)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_519),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_584),
.Y(n_600)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_519),
.Y(n_584)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_530),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_586),
.B(n_560),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_517),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_590),
.B(n_574),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_577),
.B(n_520),
.C(n_524),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_591),
.B(n_593),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_566),
.B(n_533),
.C(n_525),
.Y(n_593)
);

XNOR2x1_ASAP7_75t_L g637 ( 
.A(n_594),
.B(n_561),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_596),
.A2(n_616),
.B1(n_558),
.B2(n_564),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_566),
.B(n_525),
.C(n_548),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_602),
.C(n_605),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_575),
.B(n_539),
.C(n_545),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_578),
.B(n_532),
.C(n_545),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_562),
.Y(n_606)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_606),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_585),
.B(n_523),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_615),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_541),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_569),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_581),
.B(n_553),
.C(n_541),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_567),
.C(n_565),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_559),
.A2(n_531),
.B(n_544),
.C(n_445),
.Y(n_613)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_613),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_614),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_588),
.B(n_360),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_554),
.A2(n_430),
.B1(n_401),
.B2(n_341),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_619),
.B(n_628),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_622),
.B(n_639),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_623),
.B(n_625),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_602),
.A2(n_588),
.B(n_563),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_624),
.A2(n_638),
.B(n_603),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_601),
.B(n_570),
.C(n_572),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_626),
.A2(n_616),
.B1(n_600),
.B2(n_401),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_555),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_557),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_629),
.B(n_604),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_605),
.Y(n_630)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_630),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_608),
.A2(n_568),
.B1(n_583),
.B2(n_556),
.Y(n_632)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_632),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_601),
.B(n_555),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_633),
.B(n_635),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_591),
.B(n_560),
.C(n_580),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_634),
.B(n_640),
.C(n_612),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_593),
.B(n_579),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_576),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_598),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_637),
.B(n_609),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_597),
.A2(n_586),
.B(n_584),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_599),
.B(n_582),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_607),
.B(n_594),
.C(n_589),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_631),
.A2(n_592),
.B1(n_609),
.B2(n_589),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_641),
.B(n_650),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_645),
.A2(n_657),
.B(n_640),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_637),
.A2(n_621),
.B(n_592),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_647),
.A2(n_654),
.B(n_656),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g661 ( 
.A(n_649),
.B(n_651),
.Y(n_661)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_620),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_627),
.B(n_604),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_651),
.B(n_655),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_652),
.B(n_659),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_653),
.B(n_619),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_634),
.A2(n_595),
.B(n_598),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g656 ( 
.A1(n_618),
.A2(n_614),
.B(n_595),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_622),
.A2(n_613),
.B(n_596),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_SL g658 ( 
.A(n_633),
.B(n_607),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_628),
.Y(n_672)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_661),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_646),
.B(n_639),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_662),
.B(n_665),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_643),
.B(n_635),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_646),
.B(n_617),
.C(n_623),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_666),
.B(n_667),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_648),
.B(n_617),
.Y(n_667)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_669),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_625),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_670),
.A2(n_672),
.B(n_674),
.Y(n_687)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_651),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_671),
.B(n_627),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_652),
.B(n_636),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_647),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g679 ( 
.A(n_675),
.B(n_648),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_676),
.B(n_642),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_679),
.B(n_683),
.Y(n_696)
);

AOI21xp33_ASAP7_75t_SL g693 ( 
.A1(n_681),
.A2(n_684),
.B(n_664),
.Y(n_693)
);

AOI21xp33_ASAP7_75t_L g682 ( 
.A1(n_668),
.A2(n_649),
.B(n_660),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_682),
.A2(n_688),
.B(n_662),
.Y(n_694)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_666),
.B(n_642),
.C(n_659),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_663),
.B(n_641),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_685),
.A2(n_673),
.B(n_661),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_SL g688 ( 
.A1(n_671),
.A2(n_649),
.B1(n_657),
.B2(n_658),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_679),
.B(n_663),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_689),
.A2(n_690),
.B(n_691),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_SL g690 ( 
.A1(n_678),
.A2(n_687),
.B(n_686),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_680),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_SL g701 ( 
.A1(n_692),
.A2(n_694),
.B(n_319),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_SL g697 ( 
.A1(n_693),
.A2(n_677),
.B(n_684),
.C(n_688),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_683),
.B(n_600),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_335),
.Y(n_700)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_697),
.Y(n_703)
);

NOR3x1_ASAP7_75t_SL g699 ( 
.A(n_696),
.B(n_380),
.C(n_335),
.Y(n_699)
);

OAI311xp33_ASAP7_75t_L g702 ( 
.A1(n_699),
.A2(n_698),
.A3(n_341),
.B1(n_303),
.C1(n_178),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_700),
.B(n_701),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_702),
.A2(n_178),
.B(n_360),
.Y(n_705)
);

MAJx2_ASAP7_75t_L g706 ( 
.A(n_705),
.B(n_703),
.C(n_704),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_706),
.A2(n_8),
.B(n_9),
.Y(n_707)
);

MAJIxp5_ASAP7_75t_L g708 ( 
.A(n_707),
.B(n_10),
.C(n_234),
.Y(n_708)
);


endmodule