module real_jpeg_26264_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_105)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_7),
.A2(n_22),
.B1(n_26),
.B2(n_28),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_9),
.A2(n_34),
.B1(n_52),
.B2(n_53),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_9),
.B(n_22),
.C(n_25),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_9),
.B(n_21),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_47),
.C(n_59),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_9),
.B(n_49),
.C(n_52),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_9),
.B(n_85),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_9),
.B(n_72),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_9),
.B(n_77),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_11),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_112),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_111),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_96),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_15),
.B(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_78),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_16),
.A2(n_17),
.B1(n_68),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_37),
.B2(n_38),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_40),
.C(n_56),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_18),
.A2(n_19),
.B1(n_101),
.B2(n_110),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_18),
.B(n_129),
.C(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_18),
.A2(n_19),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_18),
.A2(n_19),
.B1(n_151),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_19),
.B(n_143),
.C(n_151),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_31),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_21),
.B(n_35),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_21),
.A2(n_32),
.B1(n_35),
.B2(n_107),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_23),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_23),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_29),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_56),
.B2(n_67),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_39),
.A2(n_40),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_54),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_42),
.B(n_91),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_44),
.A2(n_72),
.B1(n_91),
.B2(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_47),
.B(n_219),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_71),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_51),
.A2(n_90),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_52),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_63),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_63),
.B(n_76),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_57),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_64),
.B1(n_77),
.B2(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_66),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_64),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_68),
.A2(n_69),
.B(n_74),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_74),
.A2(n_106),
.B1(n_109),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_74),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_74),
.B(n_190),
.C(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_74),
.A2(n_180),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_74),
.B(n_106),
.C(n_170),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_132),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_92),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_92),
.B1(n_93),
.B2(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_89),
.B1(n_118),
.B2(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_81),
.B(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_87),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_86),
.A2(n_123),
.B(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_89),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_121),
.C(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_109),
.B1(n_129),
.B2(n_130),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_134),
.B(n_272),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_131),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_115),
.B(n_131),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.C(n_120),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_119),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_122),
.Y(n_263)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_126),
.A2(n_127),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_126),
.A2(n_127),
.B1(n_203),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_197),
.C(n_203),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_127),
.B(n_175),
.C(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_129),
.A2(n_130),
.B1(n_166),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_129),
.A2(n_130),
.B1(n_149),
.B2(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_130),
.B(n_149),
.C(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_156),
.B(n_271),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_154),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_137),
.B(n_154),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_138),
.B(n_140),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_142),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_143),
.A2(n_144),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_149),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_177),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_149),
.A2(n_163),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_149),
.B(n_220),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_266),
.B(n_270),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_193),
.B(n_252),
.C(n_265),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_182),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_159),
.B(n_182),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_169),
.B2(n_181),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_162),
.B(n_168),
.C(n_181),
.Y(n_253)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_174),
.A2(n_175),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_226),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.C(n_189),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_184),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_189),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_192),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_190),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_251),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_212),
.B(n_250),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_209),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_196),
.B(n_209),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_198),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_243),
.B(n_249),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_237),
.B(n_242),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_229),
.B(n_236),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_221),
.B(n_228),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_218),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B(n_227),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_254),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_262),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);


endmodule