module fake_jpeg_24194_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_8),
.Y(n_11)
);

BUFx2_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_9),
.B(n_14),
.C(n_16),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_31),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_32),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_19),
.B(n_18),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_9),
.C(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_40),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_4),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_26),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_6),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_33),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_39),
.B1(n_37),
.B2(n_34),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_45),
.B1(n_44),
.B2(n_46),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_33),
.B(n_32),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_34),
.B1(n_48),
.B2(n_50),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_53),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_22),
.B1(n_7),
.B2(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B1(n_57),
.B2(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_58),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_67),
.B(n_70),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_60),
.B(n_22),
.Y(n_73)
);


endmodule