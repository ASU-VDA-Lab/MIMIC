module fake_aes_50_n_16 (n_3, n_1, n_2, n_0, n_16);
input n_3;
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g4 ( .A(n_3), .Y(n_4) );
INVx2_ASAP7_75t_SL g5 ( .A(n_2), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
BUFx12f_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx2_ASAP7_75t_SL g10 ( .A(n_9), .Y(n_10) );
OAI221xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_8), .B1(n_4), .B2(n_5), .C(n_9), .Y(n_11) );
OAI32xp33_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_8), .A3(n_4), .B1(n_9), .B2(n_3), .Y(n_12) );
NAND4xp75_ASAP7_75t_L g13 ( .A(n_12), .B(n_8), .C(n_1), .D(n_2), .Y(n_13) );
AND3x2_ASAP7_75t_L g14 ( .A(n_11), .B(n_0), .C(n_1), .Y(n_14) );
OAI22x1_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_15) );
OAI21xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_14), .B(n_9), .Y(n_16) );
endmodule