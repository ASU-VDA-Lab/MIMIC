module real_jpeg_18905_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_570),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_0),
.B(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_1),
.Y(n_571)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_2),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_3),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_4),
.A2(n_31),
.B1(n_115),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_4),
.A2(n_115),
.B1(n_247),
.B2(n_251),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_4),
.A2(n_115),
.B1(n_268),
.B2(n_273),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_36),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_5),
.A2(n_36),
.B1(n_223),
.B2(n_226),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_5),
.A2(n_36),
.B1(n_280),
.B2(n_284),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_5),
.A2(n_36),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_60),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_6),
.A2(n_60),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_6),
.A2(n_60),
.B1(n_310),
.B2(n_313),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_7),
.A2(n_58),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_7),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_7),
.A2(n_182),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_7),
.A2(n_182),
.B1(n_247),
.B2(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_7),
.A2(n_182),
.B1(n_462),
.B2(n_465),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_8),
.Y(n_221)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_8),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_8),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g469 ( 
.A(n_8),
.Y(n_469)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_9),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_9),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_9),
.Y(n_441)
);

BUFx5_ASAP7_75t_L g496 ( 
.A(n_9),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_89),
.B1(n_106),
.B2(n_109),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_10),
.A2(n_89),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_10),
.A2(n_62),
.B1(n_89),
.B2(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_148),
.B1(n_192),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_11),
.A2(n_195),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_11),
.A2(n_195),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_11),
.A2(n_195),
.B1(n_490),
.B2(n_492),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_13),
.A2(n_57),
.A3(n_198),
.B1(n_200),
.B2(n_206),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_13),
.A2(n_62),
.B1(n_205),
.B2(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_13),
.B(n_38),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_13),
.B(n_97),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_13),
.B(n_65),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_13),
.B(n_479),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_13),
.A2(n_201),
.B1(n_205),
.B2(n_259),
.Y(n_498)
);

OAI32xp33_ASAP7_75t_L g500 ( 
.A1(n_13),
.A2(n_501),
.A3(n_504),
.B1(n_507),
.B2(n_508),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_15),
.Y(n_135)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_16),
.Y(n_272)
);

BUFx4f_ASAP7_75t_L g477 ( 
.A(n_16),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g143 ( 
.A(n_17),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_167),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_165),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_158),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_22),
.B(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_137),
.C(n_145),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_24),
.A2(n_137),
.B1(n_549),
.B2(n_550),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_24),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_63),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_25),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g137 ( 
.A1(n_26),
.A2(n_55),
.B(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_28),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_30),
.Y(n_322)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_34),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_35),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_37),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_37),
.A2(n_56),
.B(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_37),
.A2(n_55),
.B1(n_179),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_37),
.A2(n_55),
.B1(n_184),
.B2(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_37),
.A2(n_319),
.B(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_37),
.A2(n_160),
.B(n_394),
.Y(n_393)
);

OR2x6_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_38),
.B(n_139),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_38),
.A2(n_144),
.B1(n_178),
.B2(n_183),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_38),
.B(n_370),
.Y(n_369)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_40),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_42),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_44),
.Y(n_503)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_92),
.B1(n_93),
.B2(n_136),
.Y(n_63)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_64),
.B(n_137),
.C(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_64),
.B(n_146),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_75),
.B(n_86),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_65),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_65),
.B(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_65),
.A2(n_75),
.B1(n_417),
.B2(n_422),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_65),
.A2(n_75),
.B1(n_422),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_66),
.A2(n_243),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_66),
.B(n_87),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_66),
.A2(n_243),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_68),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_72),
.Y(n_428)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_73),
.Y(n_228)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_73),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_73),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_73),
.Y(n_453)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_73),
.Y(n_464)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_74),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_75),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_75),
.B(n_246),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_75),
.A2(n_388),
.B(n_530),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_97)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_79),
.Y(n_253)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_79),
.Y(n_283)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_84),
.Y(n_424)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_85),
.Y(n_407)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_86),
.Y(n_244)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_91),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_136),
.C(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_111),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_95),
.A2(n_119),
.B(n_190),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_96),
.A2(n_120),
.B1(n_191),
.B2(n_258),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_96),
.A2(n_120),
.B1(n_258),
.B2(n_333),
.Y(n_332)
);

OAI22x1_ASAP7_75t_L g361 ( 
.A1(n_96),
.A2(n_120),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_96),
.A2(n_120),
.B1(n_333),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_112),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_119),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_97),
.A2(n_119),
.B1(n_147),
.B2(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_105),
.A2(n_120),
.B(n_157),
.Y(n_323)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_112),
.Y(n_362)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_114),
.Y(n_335)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21x1_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_147),
.B(n_156),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_127),
.B2(n_132),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_135),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_135),
.Y(n_511)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_137),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_137),
.A2(n_550),
.B1(n_554),
.B2(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_143),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_145),
.B(n_548),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_149),
.Y(n_364)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_155),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_155),
.Y(n_367)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g573 ( 
.A(n_158),
.Y(n_573)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.CI(n_163),
.CON(n_158),
.SN(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_545),
.B(n_567),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_539),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_397),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_347),
.C(n_377),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_325),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_289),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_174),
.B(n_289),
.C(n_541),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_241),
.C(n_262),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_175),
.B(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_196),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_177),
.B(n_189),
.C(n_196),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_187),
.A2(n_188),
.B1(n_438),
.B2(n_440),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_187),
.A2(n_188),
.B1(n_448),
.B2(n_452),
.Y(n_447)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_212),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_197),
.B(n_212),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_204),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_205),
.B(n_247),
.Y(n_412)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_205),
.A2(n_412),
.B(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_205),
.A2(n_214),
.B1(n_461),
.B2(n_468),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_205),
.B(n_404),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_210),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_222),
.B1(n_229),
.B2(n_234),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_213),
.A2(n_234),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_213),
.A2(n_446),
.B1(n_454),
.B2(n_455),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_213),
.A2(n_264),
.B(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_214),
.B(n_267),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_214),
.A2(n_298),
.B(n_354),
.Y(n_353)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_214),
.A2(n_427),
.B(n_434),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_214),
.A2(n_447),
.B1(n_461),
.B2(n_466),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_215),
.Y(n_465)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_217),
.Y(n_451)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_218),
.Y(n_354)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_221),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_222),
.A2(n_306),
.B(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_241),
.B(n_262),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_254),
.C(n_257),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_242),
.B(n_257),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_243),
.A2(n_245),
.B(n_309),
.Y(n_356)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_277),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_277),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_271),
.Y(n_433)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_288),
.Y(n_277)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_283),
.Y(n_506)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_314),
.C(n_324),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_314),
.B1(n_315),
.B2(n_324),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_307),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_307),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_306),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_294),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_298),
.Y(n_518)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_305),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_R g374 ( 
.A(n_316),
.B(n_318),
.C(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_345),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_326),
.B(n_345),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.C(n_331),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_327),
.B(n_535),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_331),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_338),
.C(n_340),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_332),
.B(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_340),
.Y(n_526)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_344),
.Y(n_455)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g539 ( 
.A1(n_348),
.A2(n_540),
.B(n_542),
.C(n_543),
.D(n_544),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_349),
.B(n_350),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_373),
.B1(n_374),
.B2(n_376),
.Y(n_350)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_358),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_358),
.C(n_373),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_353),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_357),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_356),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI21xp33_ASAP7_75t_L g558 ( 
.A1(n_357),
.A2(n_395),
.B(n_559),
.Y(n_558)
);

XNOR2x1_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_368),
.C(n_381),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_368),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_377),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_378),
.B(n_379),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_380),
.B(n_383),
.C(n_391),
.Y(n_562)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_391),
.Y(n_382)
);

OA21x2_ASAP7_75t_SL g383 ( 
.A1(n_384),
.A2(n_387),
.B(n_390),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_387),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_390),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_390),
.A2(n_553),
.B1(n_556),
.B2(n_566),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_396),
.Y(n_391)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_396),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_533),
.B(n_538),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_520),
.B(n_532),
.Y(n_398)
);

OAI21x1_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_483),
.B(n_519),
.Y(n_399)
);

AOI21x1_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_443),
.B(n_482),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_425),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_402),
.B(n_425),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_415),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_403),
.A2(n_415),
.B1(n_416),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_408),
.A3(n_410),
.B1(n_412),
.B2(n_413),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_414),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_435),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_436),
.C(n_442),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_442),
.Y(n_435)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_458),
.B(n_481),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_456),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_456),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_471),
.B(n_480),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_470),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_470),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

BUFx12f_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_478),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_484),
.B(n_485),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_499),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_497),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_497),
.C(n_499),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_517),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_500),
.B(n_517),
.Y(n_528)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_512),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_SL g532 ( 
.A(n_521),
.B(n_522),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_523),
.A2(n_524),
.B1(n_527),
.B2(n_531),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_523),
.B(n_528),
.C(n_529),
.Y(n_537)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_527),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_SL g533 ( 
.A(n_534),
.B(n_537),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_534),
.B(n_537),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_561),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_546),
.A2(n_568),
.B(n_569),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_551),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_547),
.B(n_551),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_556),
.C(n_557),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_553),
.Y(n_566)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_554),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_557),
.A2(n_558),
.B1(n_564),
.B2(n_565),
.Y(n_563)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_SL g561 ( 
.A(n_562),
.B(n_563),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_562),
.B(n_563),
.Y(n_568)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);


endmodule