module real_aes_6211_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g483 ( .A1(n_0), .A2(n_166), .B(n_484), .C(n_487), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_1), .B(n_478), .Y(n_489) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g128 ( .A(n_2), .Y(n_128) );
INVx1_ASAP7_75t_L g204 ( .A(n_3), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_4), .B(n_167), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g144 ( .A1(n_5), .A2(n_145), .B1(n_146), .B2(n_452), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_5), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_5), .A2(n_98), .B1(n_452), .B2(n_751), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_6), .A2(n_463), .B(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_7), .A2(n_173), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_8), .A2(n_38), .B1(n_170), .B2(n_222), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_9), .B(n_173), .Y(n_190) );
AND2x6_ASAP7_75t_L g175 ( .A(n_10), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_11), .A2(n_175), .B(n_466), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_12), .B(n_39), .Y(n_129) );
INVx1_ASAP7_75t_L g157 ( .A(n_13), .Y(n_157) );
INVx1_ASAP7_75t_L g196 ( .A(n_14), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_15), .B(n_163), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_16), .A2(n_41), .B1(n_538), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_16), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_17), .B(n_167), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_18), .B(n_153), .Y(n_152) );
AO32x2_ASAP7_75t_L g233 ( .A1(n_19), .A2(n_173), .A3(n_174), .B1(n_193), .B2(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_20), .B(n_170), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_21), .B(n_153), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_22), .A2(n_54), .B1(n_170), .B2(n_222), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g230 ( .A1(n_23), .A2(n_83), .B1(n_163), .B2(n_170), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_24), .B(n_170), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_25), .A2(n_174), .B(n_466), .C(n_468), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_26), .A2(n_174), .B(n_466), .C(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_27), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_28), .A2(n_99), .B1(n_138), .B2(n_139), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_28), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_29), .B(n_212), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_30), .A2(n_463), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_31), .B(n_212), .Y(n_249) );
INVx2_ASAP7_75t_L g165 ( .A(n_32), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_33), .A2(n_498), .B(n_499), .C(n_503), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_34), .B(n_170), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_35), .B(n_212), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_36), .A2(n_137), .B1(n_140), .B2(n_141), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_36), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_37), .B(n_218), .Y(n_545) );
INVx1_ASAP7_75t_L g111 ( .A(n_39), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_40), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_41), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_42), .B(n_167), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_43), .B(n_463), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_44), .A2(n_498), .B(n_503), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_45), .B(n_170), .Y(n_183) );
INVx1_ASAP7_75t_L g485 ( .A(n_46), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_47), .A2(n_753), .B1(n_754), .B2(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g756 ( .A(n_47), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_48), .A2(n_92), .B1(n_222), .B2(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g524 ( .A(n_49), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_50), .B(n_170), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_51), .B(n_170), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_52), .B(n_463), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_53), .B(n_188), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g169 ( .A1(n_55), .A2(n_60), .B1(n_163), .B2(n_170), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_56), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_56), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_57), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_58), .B(n_170), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_59), .B(n_170), .Y(n_269) );
INVx1_ASAP7_75t_L g176 ( .A(n_61), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_62), .B(n_463), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_63), .B(n_478), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_64), .A2(n_188), .B(n_199), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_65), .B(n_170), .Y(n_205) );
INVx1_ASAP7_75t_L g156 ( .A(n_66), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_67), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_68), .B(n_167), .Y(n_501) );
AO32x2_ASAP7_75t_L g226 ( .A1(n_69), .A2(n_173), .A3(n_174), .B1(n_227), .B2(n_231), .Y(n_226) );
AOI222xp33_ASAP7_75t_SL g131 ( .A1(n_70), .A2(n_132), .B1(n_133), .B2(n_142), .C1(n_736), .C2(n_742), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_71), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_72), .B(n_168), .Y(n_535) );
INVx1_ASAP7_75t_L g268 ( .A(n_73), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_74), .A2(n_106), .B1(n_117), .B2(n_758), .Y(n_105) );
INVx1_ASAP7_75t_L g244 ( .A(n_75), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_76), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_77), .B(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_78), .A2(n_466), .B(n_503), .C(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_79), .B(n_163), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_80), .Y(n_511) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_82), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_84), .B(n_222), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_85), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_86), .B(n_163), .Y(n_248) );
INVx2_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_88), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_89), .B(n_160), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_90), .B(n_163), .Y(n_184) );
INVx2_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_91), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g453 ( .A(n_91), .B(n_127), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_93), .A2(n_104), .B1(n_163), .B2(n_164), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_94), .B(n_463), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_95), .Y(n_500) );
INVxp67_ASAP7_75t_L g514 ( .A(n_96), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_97), .B(n_163), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_98), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_99), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g531 ( .A(n_101), .Y(n_531) );
INVx1_ASAP7_75t_L g560 ( .A(n_102), .Y(n_560) );
AND2x2_ASAP7_75t_L g526 ( .A(n_103), .B(n_212), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx12_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g759 ( .A(n_109), .Y(n_759) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
OR2x2_ASAP7_75t_L g735 ( .A(n_113), .B(n_127), .Y(n_735) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_113), .B(n_126), .Y(n_744) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AOI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_131), .B1(n_745), .B2(n_746), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g745 ( .A(n_120), .Y(n_745) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_122), .A2(n_747), .B(n_757), .Y(n_746) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_130), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_125), .Y(n_757) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g140 ( .A(n_137), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_453), .B1(n_454), .B2(n_735), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_144), .A2(n_737), .B1(n_739), .B2(n_740), .Y(n_736) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_146), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_386), .Y(n_146) );
NOR5xp2_ASAP7_75t_L g147 ( .A(n_148), .B(n_299), .C(n_345), .D(n_358), .E(n_370), .Y(n_147) );
OAI211xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_207), .B(n_253), .C(n_280), .Y(n_148) );
INVx1_ASAP7_75t_SL g381 ( .A(n_149), .Y(n_381) );
OR2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_177), .Y(n_149) );
AND2x2_ASAP7_75t_L g305 ( .A(n_150), .B(n_178), .Y(n_305) );
AND2x2_ASAP7_75t_L g333 ( .A(n_150), .B(n_279), .Y(n_333) );
AND2x2_ASAP7_75t_L g341 ( .A(n_150), .B(n_284), .Y(n_341) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g271 ( .A(n_151), .B(n_179), .Y(n_271) );
INVx2_ASAP7_75t_L g283 ( .A(n_151), .Y(n_283) );
AND2x2_ASAP7_75t_L g408 ( .A(n_151), .B(n_350), .Y(n_408) );
OR2x2_ASAP7_75t_L g410 ( .A(n_151), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_158), .Y(n_151) );
INVx1_ASAP7_75t_L g277 ( .A(n_152), .Y(n_277) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
INVx1_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_154), .B(n_155), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NAND3xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_172), .C(n_174), .Y(n_158) );
AO21x1_ASAP7_75t_L g276 ( .A1(n_159), .A2(n_172), .B(n_277), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B1(n_166), .B2(n_169), .Y(n_159) );
INVx2_ASAP7_75t_L g223 ( .A(n_160), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g227 ( .A1(n_160), .A2(n_168), .B1(n_228), .B2(n_230), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_160), .A2(n_166), .B1(n_235), .B2(n_236), .Y(n_234) );
INVx4_ASAP7_75t_L g486 ( .A(n_160), .Y(n_486) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_161), .Y(n_201) );
INVx1_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
AND2x2_ASAP7_75t_L g464 ( .A(n_161), .B(n_189), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_161), .Y(n_467) );
INVx2_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
INVx1_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_166), .A2(n_186), .B(n_187), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_166), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_167), .A2(n_183), .B(n_184), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_SL g242 ( .A1(n_167), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_167), .A2(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_167), .B(n_514), .Y(n_513) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g243 ( .A(n_170), .Y(n_243) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_170), .Y(n_562) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
BUFx3_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
AND2x6_ASAP7_75t_L g466 ( .A(n_171), .B(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g478 ( .A(n_172), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_172), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_172), .A2(n_530), .B(n_537), .Y(n_529) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_172), .A2(n_557), .B(n_564), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_172), .B(n_565), .Y(n_564) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_173), .A2(n_181), .B(n_190), .Y(n_180) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_173), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_173), .A2(n_542), .B(n_543), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_174), .A2(n_264), .B(n_267), .Y(n_263) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_175), .A2(n_182), .B(n_185), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_175), .A2(n_195), .B(n_202), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_175), .A2(n_214), .B(n_219), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_175), .A2(n_242), .B(n_246), .Y(n_241) );
AND2x4_ASAP7_75t_L g463 ( .A(n_175), .B(n_464), .Y(n_463) );
INVx4_ASAP7_75t_SL g488 ( .A(n_175), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_175), .B(n_464), .Y(n_532) );
INVx2_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g321 ( .A(n_178), .B(n_293), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_178), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g435 ( .A(n_178), .B(n_275), .Y(n_435) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_191), .Y(n_178) );
AND2x2_ASAP7_75t_L g278 ( .A(n_179), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g325 ( .A(n_179), .Y(n_325) );
AND2x2_ASAP7_75t_L g350 ( .A(n_179), .B(n_262), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_179), .B(n_383), .Y(n_420) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g284 ( .A(n_180), .B(n_262), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_180), .B(n_261), .Y(n_298) );
AND2x2_ASAP7_75t_L g315 ( .A(n_180), .B(n_191), .Y(n_315) );
AND2x2_ASAP7_75t_L g372 ( .A(n_180), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_180), .B(n_279), .Y(n_385) );
AND2x2_ASAP7_75t_L g437 ( .A(n_180), .B(n_362), .Y(n_437) );
INVx2_ASAP7_75t_L g203 ( .A(n_188), .Y(n_203) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g260 ( .A(n_191), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g279 ( .A(n_191), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_191), .B(n_262), .Y(n_356) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_206), .Y(n_191) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_192), .A2(n_263), .B(n_270), .Y(n_262) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_193), .B(n_538), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_197), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_197), .A2(n_545), .B(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_199), .A2(n_560), .B(n_561), .C(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_200), .A2(n_247), .B(n_248), .Y(n_246) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g470 ( .A(n_201), .Y(n_470) );
O2A1O1Ixp5_ASAP7_75t_L g267 ( .A1(n_203), .A2(n_223), .B(n_268), .C(n_269), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_203), .A2(n_469), .B(n_471), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_237), .B(n_250), .Y(n_207) );
INVx1_ASAP7_75t_SL g369 ( .A(n_208), .Y(n_369) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_225), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_SL g257 ( .A(n_210), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
INVx1_ASAP7_75t_L g289 ( .A(n_211), .Y(n_289) );
AND2x2_ASAP7_75t_L g310 ( .A(n_211), .B(n_232), .Y(n_310) );
AND2x2_ASAP7_75t_L g344 ( .A(n_211), .B(n_233), .Y(n_344) );
OR2x2_ASAP7_75t_L g363 ( .A(n_211), .B(n_239), .Y(n_363) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_211), .Y(n_377) );
AND2x2_ASAP7_75t_L g390 ( .A(n_211), .B(n_391), .Y(n_390) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_224), .Y(n_211) );
INVx2_ASAP7_75t_L g231 ( .A(n_212), .Y(n_231) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_212), .A2(n_241), .B(n_249), .Y(n_240) );
INVx1_ASAP7_75t_L g476 ( .A(n_212), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_212), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_212), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_223), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_225), .A2(n_312), .B1(n_313), .B2(n_322), .Y(n_311) );
AND2x2_ASAP7_75t_L g395 ( .A(n_225), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_232), .Y(n_225) );
INVx1_ASAP7_75t_L g256 ( .A(n_226), .Y(n_256) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_226), .Y(n_293) );
INVx1_ASAP7_75t_L g304 ( .A(n_226), .Y(n_304) );
AND2x2_ASAP7_75t_L g319 ( .A(n_226), .B(n_233), .Y(n_319) );
INVx2_ASAP7_75t_L g487 ( .A(n_229), .Y(n_487) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_229), .Y(n_502) );
INVx1_ASAP7_75t_L g473 ( .A(n_231), .Y(n_473) );
OR2x2_ASAP7_75t_L g273 ( .A(n_232), .B(n_258), .Y(n_273) );
AND2x2_ASAP7_75t_L g303 ( .A(n_232), .B(n_304), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_232), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g251 ( .A(n_233), .B(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g360 ( .A(n_233), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_237), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g338 ( .A(n_238), .B(n_304), .Y(n_338) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g250 ( .A(n_239), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g309 ( .A(n_239), .Y(n_309) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g258 ( .A(n_240), .Y(n_258) );
OR2x2_ASAP7_75t_L g288 ( .A(n_240), .B(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_240), .Y(n_343) );
AOI32xp33_ASAP7_75t_L g380 ( .A1(n_250), .A2(n_310), .A3(n_381), .B1(n_382), .B2(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g306 ( .A(n_251), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_251), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_251), .B(n_338), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_251), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_259), .B1(n_272), .B2(n_274), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
AND2x2_ASAP7_75t_L g359 ( .A(n_255), .B(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_256), .B(n_258), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_257), .A2(n_281), .B1(n_285), .B2(n_295), .Y(n_280) );
AND2x2_ASAP7_75t_L g302 ( .A(n_257), .B(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_257), .A2(n_271), .B(n_319), .C(n_354), .Y(n_353) );
OAI332xp33_ASAP7_75t_L g358 ( .A1(n_257), .A2(n_359), .A3(n_361), .B1(n_363), .B2(n_364), .B3(n_366), .C1(n_367), .C2(n_369), .Y(n_358) );
INVx2_ASAP7_75t_L g399 ( .A(n_257), .Y(n_399) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
INVx1_ASAP7_75t_L g392 ( .A(n_258), .Y(n_392) );
AND2x2_ASAP7_75t_L g446 ( .A(n_258), .B(n_310), .Y(n_446) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_271), .Y(n_259) );
AND2x2_ASAP7_75t_L g326 ( .A(n_261), .B(n_276), .Y(n_326) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g275 ( .A(n_262), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g374 ( .A(n_262), .B(n_276), .Y(n_374) );
INVx1_ASAP7_75t_L g383 ( .A(n_262), .Y(n_383) );
INVx1_ASAP7_75t_L g357 ( .A(n_271), .Y(n_357) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g441 ( .A(n_273), .B(n_293), .Y(n_441) );
INVx1_ASAP7_75t_SL g352 ( .A(n_274), .Y(n_352) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
AND2x2_ASAP7_75t_L g379 ( .A(n_275), .B(n_337), .Y(n_379) );
INVx1_ASAP7_75t_L g398 ( .A(n_275), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_275), .B(n_365), .Y(n_400) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
AND2x2_ASAP7_75t_L g301 ( .A(n_278), .B(n_282), .Y(n_301) );
AND2x2_ASAP7_75t_L g368 ( .A(n_278), .B(n_326), .Y(n_368) );
INVx2_ASAP7_75t_L g411 ( .A(n_278), .Y(n_411) );
INVx2_ASAP7_75t_L g294 ( .A(n_279), .Y(n_294) );
AND2x2_ASAP7_75t_L g296 ( .A(n_279), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g312 ( .A(n_282), .Y(n_312) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_283), .B(n_356), .Y(n_362) );
OR2x2_ASAP7_75t_L g426 ( .A(n_283), .B(n_385), .Y(n_426) );
INVx1_ASAP7_75t_L g450 ( .A(n_283), .Y(n_450) );
INVx1_ASAP7_75t_L g406 ( .A(n_284), .Y(n_406) );
AND2x2_ASAP7_75t_L g451 ( .A(n_284), .B(n_294), .Y(n_451) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_288), .A2(n_314), .B1(n_316), .B2(n_320), .Y(n_313) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI322xp33_ASAP7_75t_SL g397 ( .A1(n_291), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_401), .C1(n_404), .C2(n_406), .Y(n_397) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
AND2x2_ASAP7_75t_L g394 ( .A(n_292), .B(n_310), .Y(n_394) );
OR2x2_ASAP7_75t_L g428 ( .A(n_292), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g431 ( .A(n_292), .B(n_363), .Y(n_431) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g376 ( .A(n_293), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g432 ( .A(n_293), .B(n_363), .Y(n_432) );
INVx3_ASAP7_75t_L g365 ( .A(n_294), .Y(n_365) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g421 ( .A(n_296), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g300 ( .A1(n_298), .A2(n_301), .B1(n_302), .B2(n_305), .C1(n_306), .C2(n_308), .Y(n_300) );
INVx1_ASAP7_75t_L g331 ( .A(n_298), .Y(n_331) );
NAND3xp33_ASAP7_75t_SL g299 ( .A(n_300), .B(n_311), .C(n_328), .Y(n_299) );
AND2x2_ASAP7_75t_L g416 ( .A(n_303), .B(n_317), .Y(n_416) );
BUFx2_ASAP7_75t_L g307 ( .A(n_304), .Y(n_307) );
INVx1_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_305), .A2(n_341), .B1(n_394), .B2(n_395), .C(n_397), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_307), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
AND2x2_ASAP7_75t_L g347 ( .A(n_310), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_315), .B(n_326), .Y(n_327) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OAI21xp33_ASAP7_75t_L g322 ( .A1(n_317), .A2(n_323), .B(n_327), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_317), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g414 ( .A(n_319), .B(n_396), .Y(n_414) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g337 ( .A(n_325), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_326), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g443 ( .A(n_326), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_334), .B1(n_335), .B2(n_338), .C(n_339), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_330), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g439 ( .A(n_338), .B(n_344), .Y(n_439) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OAI31xp33_ASAP7_75t_SL g407 ( .A1(n_342), .A2(n_381), .A3(n_408), .B(n_409), .Y(n_407) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g396 ( .A(n_343), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_344), .B(n_348), .Y(n_447) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_349), .B1(n_351), .B2(n_352), .C(n_353), .Y(n_345) );
INVx1_ASAP7_75t_L g351 ( .A(n_347), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_350), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g366 ( .A(n_359), .Y(n_366) );
INVx2_ASAP7_75t_L g402 ( .A(n_360), .Y(n_402) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g388 ( .A(n_365), .B(n_374), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_365), .A2(n_382), .B(n_439), .C(n_440), .Y(n_438) );
OAI221xp5_ASAP7_75t_SL g370 ( .A1(n_366), .A2(n_371), .B1(n_375), .B2(n_378), .C(n_380), .Y(n_370) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_369), .A2(n_434), .B(n_436), .C(n_438), .Y(n_433) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_372), .A2(n_423), .B1(n_425), .B2(n_427), .C(n_430), .Y(n_422) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NOR4xp25_ASAP7_75t_L g386 ( .A(n_387), .B(n_412), .C(n_433), .D(n_444), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .B(n_393), .C(n_407), .Y(n_387) );
INVx1_ASAP7_75t_SL g442 ( .A(n_394), .Y(n_442) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_403), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_410), .A2(n_419), .B1(n_431), .B2(n_432), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B(n_417), .C(n_422), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI31xp33_ASAP7_75t_L g444 ( .A1(n_415), .A2(n_445), .A3(n_447), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g738 ( .A(n_453), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_454), .Y(n_739) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_455), .B(n_671), .Y(n_454) );
NOR5xp2_ASAP7_75t_L g455 ( .A(n_456), .B(n_602), .C(n_631), .D(n_651), .E(n_658), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_490), .B(n_547), .C(n_589), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_458), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_673) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_477), .Y(n_458) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_459), .Y(n_550) );
AND2x4_ASAP7_75t_L g582 ( .A(n_459), .B(n_583), .Y(n_582) );
INVx5_ASAP7_75t_L g600 ( .A(n_459), .Y(n_600) );
AND2x2_ASAP7_75t_L g609 ( .A(n_459), .B(n_601), .Y(n_609) );
AND2x2_ASAP7_75t_L g621 ( .A(n_459), .B(n_494), .Y(n_621) );
AND2x2_ASAP7_75t_L g717 ( .A(n_459), .B(n_585), .Y(n_717) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
AOI21xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_465), .B(n_473), .Y(n_460) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx5_ASAP7_75t_L g482 ( .A(n_466), .Y(n_482) );
INVx2_ASAP7_75t_L g472 ( .A(n_470), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_472), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_472), .A2(n_502), .B(n_524), .C(n_525), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx2_ASAP7_75t_L g583 ( .A(n_477), .Y(n_583) );
AND2x2_ASAP7_75t_L g601 ( .A(n_477), .B(n_556), .Y(n_601) );
AND2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_555), .Y(n_620) );
AND2x2_ASAP7_75t_L g660 ( .A(n_477), .B(n_600), .Y(n_660) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_489), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_482), .B(n_483), .C(n_488), .Y(n_480) );
INVx2_ASAP7_75t_L g498 ( .A(n_482), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_482), .A2(n_488), .B(n_511), .C(n_512), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g503 ( .A(n_488), .Y(n_503) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_516), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI322xp5_ASAP7_75t_L g719 ( .A1(n_493), .A2(n_527), .A3(n_574), .B1(n_582), .B2(n_636), .C1(n_720), .C2(n_723), .Y(n_719) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .Y(n_493) );
INVx5_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
AND2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_554), .Y(n_568) );
BUFx2_ASAP7_75t_L g646 ( .A(n_494), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_494), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g723 ( .A(n_494), .B(n_630), .Y(n_723) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_506), .B(n_518), .Y(n_577) );
INVx1_ASAP7_75t_L g604 ( .A(n_506), .Y(n_604) );
AND2x2_ASAP7_75t_L g617 ( .A(n_506), .B(n_539), .Y(n_617) );
AND2x2_ASAP7_75t_L g718 ( .A(n_506), .B(n_636), .Y(n_718) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g572 ( .A(n_507), .B(n_518), .Y(n_572) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_507), .Y(n_580) );
OR2x2_ASAP7_75t_L g587 ( .A(n_507), .B(n_539), .Y(n_587) );
AND2x2_ASAP7_75t_L g597 ( .A(n_507), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_507), .B(n_529), .Y(n_626) );
INVxp67_ASAP7_75t_L g650 ( .A(n_507), .Y(n_650) );
AND2x2_ASAP7_75t_L g657 ( .A(n_507), .B(n_527), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_507), .B(n_539), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_507), .B(n_528), .Y(n_683) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_507) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_518), .B(n_540), .Y(n_627) );
OR2x2_ASAP7_75t_L g649 ( .A(n_518), .B(n_528), .Y(n_649) );
AND2x2_ASAP7_75t_L g662 ( .A(n_518), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_518), .B(n_617), .Y(n_668) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_518), .A2(n_673), .B(n_678), .C(n_687), .Y(n_672) );
AND2x2_ASAP7_75t_L g733 ( .A(n_518), .B(n_539), .Y(n_733) );
INVx5_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g586 ( .A(n_519), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_519), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_519), .B(n_581), .Y(n_593) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_519), .Y(n_595) );
OR2x2_ASAP7_75t_L g606 ( .A(n_519), .B(n_528), .Y(n_606) );
AND2x2_ASAP7_75t_SL g611 ( .A(n_519), .B(n_597), .Y(n_611) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_528), .Y(n_636) );
AND2x2_ASAP7_75t_L g656 ( .A(n_519), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g694 ( .A(n_519), .B(n_527), .Y(n_694) );
OR2x2_ASAP7_75t_L g697 ( .A(n_519), .B(n_683), .Y(n_697) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_526), .Y(n_519) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_528), .A2(n_641), .B(n_644), .C(n_650), .Y(n_640) );
INVx5_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_529), .B(n_539), .Y(n_571) );
AND2x2_ASAP7_75t_L g575 ( .A(n_529), .B(n_540), .Y(n_575) );
OR2x2_ASAP7_75t_L g581 ( .A(n_529), .B(n_539), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_SL g598 ( .A(n_539), .Y(n_598) );
OR2x2_ASAP7_75t_L g726 ( .A(n_539), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_566), .B(n_569), .C(n_578), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI31xp33_ASAP7_75t_L g651 ( .A1(n_549), .A2(n_652), .A3(n_654), .B(n_655), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_550), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_551), .B(n_582), .Y(n_588) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_552), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g608 ( .A(n_552), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g613 ( .A(n_552), .B(n_583), .Y(n_613) );
AND2x2_ASAP7_75t_L g623 ( .A(n_552), .B(n_582), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_552), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g643 ( .A(n_552), .B(n_600), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_552), .B(n_620), .Y(n_648) );
OR2x2_ASAP7_75t_L g667 ( .A(n_552), .B(n_554), .Y(n_667) );
OR2x2_ASAP7_75t_L g669 ( .A(n_552), .B(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_552), .Y(n_716) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g616 ( .A(n_554), .B(n_583), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_554), .B(n_600), .Y(n_639) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx2_ASAP7_75t_L g585 ( .A(n_556), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g676 ( .A(n_568), .B(n_600), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g678 ( .A1(n_568), .A2(n_582), .A3(n_620), .B1(n_679), .B2(n_680), .C1(n_681), .C2(n_684), .Y(n_678) );
INVx1_ASAP7_75t_L g686 ( .A(n_568), .Y(n_686) );
NAND2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx1_ASAP7_75t_SL g680 ( .A(n_570), .Y(n_680) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
OR2x2_ASAP7_75t_L g632 ( .A(n_571), .B(n_577), .Y(n_632) );
INVx1_ASAP7_75t_L g663 ( .A(n_571), .Y(n_663) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI32xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .A3(n_584), .B1(n_586), .B2(n_588), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_581), .A2(n_596), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g633 ( .A(n_582), .Y(n_633) );
AND2x4_ASAP7_75t_L g630 ( .A(n_583), .B(n_600), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_583), .B(n_666), .Y(n_665) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_584), .A2(n_611), .A3(n_630), .B1(n_663), .B2(n_696), .C1(n_698), .C2(n_699), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_584), .A2(n_661), .B1(n_725), .B2(n_726), .C(n_728), .Y(n_724) );
AND2x2_ASAP7_75t_L g612 ( .A(n_585), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g592 ( .A(n_587), .Y(n_592) );
OR2x2_ASAP7_75t_L g664 ( .A(n_587), .B(n_649), .Y(n_664) );
OAI31xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .A3(n_594), .B(n_599), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_590), .A2(n_623), .B1(n_624), .B2(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g635 ( .A(n_592), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_594), .A2(n_635), .B1(n_688), .B2(n_691), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g677 ( .A(n_597), .B(n_646), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_597), .B(n_636), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_598), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g711 ( .A(n_598), .B(n_649), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_599), .A2(n_694), .B1(n_707), .B2(n_710), .Y(n_706) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx2_ASAP7_75t_L g615 ( .A(n_600), .Y(n_615) );
AND2x2_ASAP7_75t_L g698 ( .A(n_600), .B(n_620), .Y(n_698) );
OR2x2_ASAP7_75t_L g700 ( .A(n_600), .B(n_667), .Y(n_700) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_600), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_601), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_601), .B(n_646), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_607), .B(n_610), .C(n_622), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_614), .B2(n_617), .C(n_618), .Y(n_610) );
INVxp67_ASAP7_75t_L g722 ( .A(n_613), .Y(n_722) );
INVx1_ASAP7_75t_L g689 ( .A(n_614), .Y(n_689) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g653 ( .A(n_615), .B(n_620), .Y(n_653) );
INVx1_ASAP7_75t_L g670 ( .A(n_616), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_616), .B(n_643), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g685 ( .A(n_620), .Y(n_685) );
AND2x2_ASAP7_75t_L g691 ( .A(n_620), .B(n_646), .Y(n_691) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_SL g679 ( .A(n_627), .Y(n_679) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_630), .B(n_666), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_637), .C(n_640), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g727 ( .A(n_636), .Y(n_727) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g645 ( .A(n_639), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_643), .B(n_702), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B(n_649), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g692 ( .A1(n_647), .A2(n_693), .B(n_695), .C(n_701), .Y(n_692) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g704 ( .A(n_649), .Y(n_704) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI222xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B1(n_664), .B2(n_665), .C1(n_668), .C2(n_669), .Y(n_658) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g734 ( .A(n_665), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_666), .B(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_666), .A2(n_713), .B1(n_715), .B2(n_718), .Y(n_712) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
NOR4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_692), .C(n_705), .D(n_724), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_674), .B(n_704), .Y(n_714) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g681 ( .A(n_679), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_682), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_712), .C(n_719), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx2_ASAP7_75t_L g721 ( .A(n_717), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_731), .B(n_734), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g741 ( .A(n_735), .Y(n_741) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
XOR2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule