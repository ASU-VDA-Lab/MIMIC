module fake_jpeg_22464_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_7),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_41),
.CON(n_76),
.SN(n_76)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_19),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

CKINVDCx9p33_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_16),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_32),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_72),
.Y(n_106)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_64),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_18),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_17),
.B(n_21),
.C(n_22),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_78),
.A2(n_104),
.B(n_24),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_17),
.B1(n_21),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_81),
.A2(n_83),
.B1(n_25),
.B2(n_26),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_77),
.B1(n_58),
.B2(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_96),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_97),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_103),
.B1(n_108),
.B2(n_24),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_17),
.B1(n_47),
.B2(n_23),
.Y(n_103)
);

NAND2x1_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_35),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_63),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_35),
.B1(n_20),
.B2(n_30),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_16),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_31),
.B(n_26),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_31),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_35),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_122),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_51),
.B1(n_67),
.B2(n_22),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_118),
.A2(n_125),
.B1(n_143),
.B2(n_99),
.Y(n_169)
);

MAJx3_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_31),
.C(n_25),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_92),
.C(n_109),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_120),
.A2(n_89),
.B(n_23),
.Y(n_175)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_65),
.B(n_26),
.C(n_23),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_124),
.B(n_112),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_34),
.B(n_29),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_135),
.B1(n_99),
.B2(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_102),
.B1(n_89),
.B2(n_100),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_133),
.Y(n_179)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_92),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_158),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_106),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_138),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_103),
.B(n_109),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_175),
.B(n_180),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_166),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_103),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_165),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_85),
.B1(n_90),
.B2(n_114),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_170),
.B1(n_176),
.B2(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_168),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

AO21x1_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_34),
.B(n_9),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_110),
.C(n_102),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_173),
.C(n_127),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_103),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_123),
.B1(n_134),
.B2(n_136),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_82),
.B1(n_90),
.B2(n_52),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_82),
.B1(n_52),
.B2(n_101),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_34),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_145),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_120),
.A2(n_98),
.B(n_97),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_183),
.B(n_190),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_171),
.C(n_148),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_149),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_194),
.B(n_201),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_125),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_124),
.B1(n_133),
.B2(n_141),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_172),
.B1(n_153),
.B2(n_162),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_157),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_25),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_152),
.B(n_25),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_203),
.A2(n_204),
.B(n_208),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_145),
.B1(n_84),
.B2(n_80),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_212),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_213),
.B(n_175),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_34),
.B(n_1),
.C(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_220),
.C(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_150),
.C(n_148),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_227),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_172),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_224),
.A2(n_231),
.B(n_2),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_146),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_151),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_199),
.B1(n_204),
.B2(n_210),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_158),
.A3(n_165),
.B1(n_156),
.B2(n_152),
.C1(n_153),
.C2(n_162),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_239),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_156),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_200),
.C(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_182),
.B(n_179),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_245),
.A2(n_237),
.B1(n_264),
.B2(n_219),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_193),
.B1(n_187),
.B2(n_213),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_195),
.C(n_200),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_250),
.C(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_206),
.C(n_202),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_256),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_155),
.B(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_186),
.C(n_155),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_260),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_203),
.C(n_178),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_183),
.B1(n_208),
.B2(n_155),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_203),
.C(n_184),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_220),
.C(n_238),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_SL g262 ( 
.A1(n_218),
.A2(n_188),
.A3(n_214),
.B1(n_211),
.B2(n_11),
.C1(n_13),
.C2(n_7),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_262),
.B(n_13),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_9),
.Y(n_263)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_10),
.B(n_14),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_233),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_272),
.C(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_250),
.B(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_12),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_215),
.C(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_223),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_275),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_285),
.B1(n_261),
.B2(n_239),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_222),
.C(n_232),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_266),
.C(n_3),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_265),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_245),
.A2(n_232),
.B1(n_240),
.B2(n_226),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_248),
.CI(n_249),
.CON(n_287),
.SN(n_287)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_253),
.B1(n_243),
.B2(n_251),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_293),
.B1(n_268),
.B2(n_267),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_244),
.B1(n_251),
.B2(n_256),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_254),
.B(n_258),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_300),
.B(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_255),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_297),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_298),
.C(n_267),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_14),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_2),
.C(n_3),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_302),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_277),
.B(n_281),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_307),
.B(n_314),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_279),
.C(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_311),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_270),
.B(n_272),
.C(n_271),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_305),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_295),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_276),
.B(n_12),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_289),
.C(n_309),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_319),
.B(n_321),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_296),
.B(n_298),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_289),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_3),
.C(n_4),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_324),
.B(n_307),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_12),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_303),
.C(n_307),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_315),
.CI(n_306),
.CON(n_327),
.SN(n_327)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_329),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_316),
.B1(n_318),
.B2(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_331),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_325),
.A2(n_307),
.B1(n_4),
.B2(n_5),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_6),
.B(n_3),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_13),
.B(n_4),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_334),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_337),
.B(n_338),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_326),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_336),
.C(n_5),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_5),
.C(n_6),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_5),
.Y(n_342)
);


endmodule