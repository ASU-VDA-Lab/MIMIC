module fake_jpeg_27933_n_106 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_10),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_12),
.B1(n_15),
.B2(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_23),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_27),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_15),
.B1(n_17),
.B2(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_51),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_60),
.B1(n_38),
.B2(n_13),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_29),
.B(n_26),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_61),
.B1(n_62),
.B2(n_16),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_20),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_25),
.B1(n_33),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_19),
.B1(n_17),
.B2(n_33),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_13),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_69),
.B1(n_61),
.B2(n_57),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_80),
.B1(n_68),
.B2(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_48),
.B1(n_65),
.B2(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_49),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_65),
.B1(n_72),
.B2(n_53),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_59),
.C(n_55),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_81),
.C(n_84),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_60),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_82),
.C(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_14),
.Y(n_93)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.C(n_94),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_38),
.C(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_3),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_4),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_86),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_90),
.C(n_86),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_7),
.C(n_9),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_11),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_9),
.C(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);


endmodule