module real_jpeg_29386_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_37),
.B1(n_56),
.B2(n_58),
.Y(n_160)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_4),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_29),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_31),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_61),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_4),
.B(n_61),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_76),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_4),
.A2(n_123),
.B1(n_140),
.B2(n_206),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_4),
.A2(n_32),
.B(n_221),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_5),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_113),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_113),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_5),
.A2(n_56),
.B1(n_58),
.B2(n_113),
.Y(n_206)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_7),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_98),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_98),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_98),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_96),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_96),
.Y(n_200)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_279)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_12),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_103),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_12),
.A2(n_56),
.B1(n_58),
.B2(n_103),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_103),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_13),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_106),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_106),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_14),
.A2(n_27),
.B1(n_56),
.B2(n_58),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_14),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_269)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_17),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_17),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_22),
.B(n_43),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_24),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_35),
.B(n_110),
.C(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_28),
.A2(n_31),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_28),
.A2(n_31),
.B1(n_148),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_28),
.A2(n_31),
.B1(n_167),
.B2(n_260),
.Y(n_259)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_31),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_68),
.B(n_70),
.C(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_71),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g229 ( 
.A1(n_32),
.A2(n_62),
.A3(n_68),
.B1(n_222),
.B2(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_33),
.B(n_110),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_84),
.B(n_335),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_77),
.C(n_79),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_44),
.A2(n_45),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_64),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_46),
.B(n_319),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_48),
.A2(n_81),
.B1(n_83),
.B2(n_287),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_52),
.A2(n_310),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_52),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_52),
.A2(n_64),
.B1(n_313),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_63),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_53),
.A2(n_59),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_53),
.A2(n_59),
.B1(n_138),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_53),
.A2(n_59),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_53),
.A2(n_59),
.B1(n_181),
.B2(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_53),
.B(n_110),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_53),
.A2(n_59),
.B1(n_102),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_53),
.A2(n_59),
.B1(n_63),
.B2(n_269),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_54),
.A2(n_58),
.A3(n_61),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_55),
.B(n_56),
.Y(n_185)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_56),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_61),
.B(n_74),
.Y(n_230)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_65),
.A2(n_66),
.B1(n_76),
.B2(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_76),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_66),
.A2(n_76),
.B1(n_151),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_66),
.A2(n_76),
.B1(n_169),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_73),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_73),
.B1(n_94),
.B2(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_67),
.A2(n_73),
.B1(n_97),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_67),
.A2(n_73),
.B1(n_129),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_67),
.A2(n_73),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_77),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_81),
.A2(n_83),
.B1(n_112),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_81),
.A2(n_83),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_328),
.B(n_334),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_304),
.A3(n_323),
.B1(n_326),
.B2(n_327),
.C(n_339),
.Y(n_85)
);

AOI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_256),
.A3(n_293),
.B1(n_298),
.B2(n_303),
.C(n_340),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_153),
.C(n_171),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_133),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_89),
.B(n_133),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_114),
.C(n_125),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_90),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_108),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_100),
.C(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_104),
.A2(n_107),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_104),
.A2(n_107),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_110),
.B(n_123),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_114),
.A2(n_125),
.B1(n_126),
.B2(n_254),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_114),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_117),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_118),
.A2(n_122),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_140),
.B1(n_142),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_123),
.A2(n_140),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_123),
.A2(n_140),
.B1(n_200),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_123),
.A2(n_140),
.B1(n_195),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_123),
.A2(n_140),
.B(n_160),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_132),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_127),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_130),
.B(n_132),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_143),
.C(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_139),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_149),
.C(n_152),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_154),
.A2(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_155),
.B(n_156),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_170),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_163),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_158),
.B(n_163),
.C(n_170),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_159),
.B(n_161),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_250),
.B(n_255),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_236),
.B(n_249),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_215),
.B(n_235),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_196),
.B(n_214),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_186),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_194),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B(n_213),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_202),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_208),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_216),
.B(n_217),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_228),
.B1(n_233),
.B2(n_234),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_227),
.C(n_234),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_231),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_245),
.C(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_273),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_273),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.C(n_272),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_264),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_258),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.CI(n_263),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_261),
.C(n_263),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_270),
.B2(n_271),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_271),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_285),
.B(n_288),
.Y(n_315)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_291),
.B2(n_292),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_282),
.C(n_292),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B(n_281),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_280),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_279),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_306),
.C(n_315),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_281),
.B(n_306),
.CI(n_315),
.CON(n_325),
.SN(n_325)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_282)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_299),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_296),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_316),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_316),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_314),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_310),
.C(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_321),
.C(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_325),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);


endmodule