module fake_jpeg_10238_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_24),
.C(n_32),
.Y(n_65)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_52),
.B1(n_42),
.B2(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_21),
.B1(n_19),
.B2(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_33),
.B(n_31),
.C(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_42),
.B1(n_37),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_24),
.B1(n_18),
.B2(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_17),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_17),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_72),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_80),
.B1(n_82),
.B2(n_63),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_34),
.B1(n_24),
.B2(n_18),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_27),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_47),
.B1(n_55),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_46),
.B1(n_62),
.B2(n_53),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_0),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_67),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_83),
.C(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_91),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_62),
.B1(n_49),
.B2(n_44),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_49),
.B1(n_63),
.B2(n_60),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_119),
.B1(n_73),
.B2(n_82),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_25),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g115 ( 
.A(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_79),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_43),
.B1(n_39),
.B2(n_22),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_79),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_89),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_27),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_98),
.B(n_96),
.Y(n_154)
);

AO21x2_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_73),
.B(n_70),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_98),
.B1(n_103),
.B2(n_76),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_81),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_143),
.B1(n_96),
.B2(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_117),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_136),
.B(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_22),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_139),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_43),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_95),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_22),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_142),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_23),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_30),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_0),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_1),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_114),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_150),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_161),
.C(n_164),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_163),
.B(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_168),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_171),
.B1(n_74),
.B2(n_112),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_142),
.B1(n_135),
.B2(n_144),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_162),
.B1(n_166),
.B2(n_155),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_100),
.B1(n_97),
.B2(n_103),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_123),
.B(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_173),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_100),
.B1(n_119),
.B2(n_93),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_115),
.B1(n_114),
.B2(n_30),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_22),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_107),
.B(n_112),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_131),
.B(n_127),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_124),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_193),
.C(n_162),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_196),
.B1(n_181),
.B2(n_179),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_130),
.B(n_146),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_187),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_194),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_166),
.B1(n_147),
.B2(n_22),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_R g191 ( 
.A(n_154),
.B(n_146),
.C(n_125),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_167),
.C(n_152),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_151),
.C(n_163),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_125),
.C(n_139),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_22),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_210),
.C(n_211),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_209),
.Y(n_226)
);

OAI221xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_191),
.B1(n_218),
.B2(n_195),
.C(n_200),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_156),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_149),
.C(n_173),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_193),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_186),
.B1(n_180),
.B2(n_194),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_215),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_147),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_217),
.C(n_210),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_107),
.C(n_17),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_223),
.B1(n_225),
.B2(n_228),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_228),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_190),
.B(n_184),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_207),
.B1(n_216),
.B2(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_232),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_203),
.A2(n_184),
.B(n_197),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_217),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_205),
.C(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_177),
.C(n_17),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_178),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_226),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_235),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_245),
.C(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_247),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_239),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_230),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_236),
.B(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_256),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_258),
.C(n_255),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_233),
.B1(n_234),
.B2(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_7),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_246),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_5),
.B(n_6),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_254),
.B(n_257),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_240),
.B(n_5),
.Y(n_256)
);

AOI321xp33_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_12),
.C(n_13),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_237),
.B1(n_8),
.B2(n_9),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_266),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_258),
.A2(n_7),
.B(n_8),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_265),
.B(n_13),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_11),
.C(n_12),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_260),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

OA21x2_ASAP7_75t_SL g275 ( 
.A1(n_273),
.A2(n_268),
.B(n_15),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_274),
.C(n_14),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_16),
.C(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_16),
.Y(n_279)
);


endmodule