module fake_jpeg_25918_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_0),
.CON(n_38),
.SN(n_38)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_17),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_24),
.B(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_24),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_59),
.B1(n_74),
.B2(n_78),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_27),
.B1(n_23),
.B2(n_18),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_45),
.B1(n_48),
.B2(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_25),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_19),
.C(n_32),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_24),
.C(n_32),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_63),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_72),
.Y(n_93)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_17),
.B1(n_22),
.B2(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_34),
.B1(n_20),
.B2(n_49),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_17),
.B1(n_22),
.B2(n_36),
.Y(n_81)
);

OAI22x1_ASAP7_75t_L g146 ( 
.A1(n_81),
.A2(n_104),
.B1(n_35),
.B2(n_34),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_82),
.B(n_102),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_47),
.B1(n_39),
.B2(n_22),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_115),
.B1(n_36),
.B2(n_37),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_85),
.B(n_106),
.Y(n_131)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_49),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_111),
.Y(n_152)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_99),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_41),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_31),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_36),
.B1(n_38),
.B2(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_117),
.Y(n_135)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_109),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_76),
.B1(n_66),
.B2(n_20),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_21),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_58),
.A2(n_39),
.B1(n_70),
.B2(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_52),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_71),
.B1(n_60),
.B2(n_20),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_120),
.A2(n_149),
.B1(n_109),
.B2(n_86),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_122),
.B(n_136),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_36),
.B1(n_37),
.B2(n_25),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_20),
.B1(n_34),
.B2(n_49),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_124),
.A2(n_108),
.B1(n_114),
.B2(n_94),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_21),
.B1(n_25),
.B2(n_31),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_151),
.B1(n_103),
.B2(n_100),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_86),
.B1(n_90),
.B2(n_87),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_9),
.B(n_16),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_120),
.B(n_131),
.C(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_89),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_41),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_31),
.B1(n_32),
.B2(n_41),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_153),
.B(n_166),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_161),
.B1(n_175),
.B2(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_88),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_96),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_163),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_113),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_88),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

AO21x2_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_142),
.B(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_182),
.B1(n_128),
.B2(n_124),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_134),
.B1(n_127),
.B2(n_148),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_85),
.B(n_94),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_177),
.B(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_178),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_172),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_85),
.B(n_2),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_92),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_92),
.A3(n_89),
.B1(n_103),
.B2(n_100),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_133),
.A2(n_79),
.B1(n_31),
.B2(n_8),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_181),
.B1(n_133),
.B2(n_143),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_133),
.A2(n_79),
.B1(n_31),
.B2(n_7),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_32),
.B1(n_15),
.B2(n_10),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_1),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_185),
.B(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_199),
.B1(n_206),
.B2(n_161),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_177),
.B(n_131),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_156),
.B1(n_184),
.B2(n_164),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_210),
.B(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_185),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_122),
.B1(n_147),
.B2(n_134),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_141),
.B1(n_125),
.B2(n_139),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_141),
.B1(n_125),
.B2(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_211),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_145),
.C(n_15),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_10),
.C(n_9),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_217),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_155),
.A2(n_1),
.B(n_2),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_1),
.B(n_2),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_10),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_166),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_7),
.C(n_2),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_220),
.Y(n_264)
);

XOR2x2_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_188),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_190),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_227),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_237),
.B(n_244),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_161),
.B1(n_175),
.B2(n_164),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_228),
.Y(n_266)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_195),
.B1(n_206),
.B2(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_208),
.B1(n_187),
.B2(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_189),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_153),
.B1(n_170),
.B2(n_182),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_209),
.A2(n_162),
.B1(n_173),
.B2(n_167),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_173),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_1),
.B(n_3),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_250),
.B1(n_252),
.B2(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_188),
.C(n_198),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_261),
.C(n_265),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_217),
.B(n_214),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_187),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_257),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_259),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_213),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_221),
.A2(n_193),
.B1(n_215),
.B2(n_192),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_193),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_200),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_243),
.C(n_240),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_277),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_233),
.C(n_235),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_261),
.C(n_249),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_224),
.C(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_279),
.C(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_224),
.C(n_220),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_254),
.B(n_227),
.CI(n_222),
.CON(n_280),
.SN(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_285),
.B1(n_266),
.B2(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_232),
.C(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_236),
.C(n_238),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_246),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_231),
.B1(n_260),
.B2(n_227),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_293),
.B1(n_298),
.B2(n_192),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_273),
.B(n_268),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_246),
.B1(n_229),
.B2(n_219),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_3),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_269),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_267),
.B1(n_244),
.B2(n_237),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_251),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_223),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_255),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_186),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_275),
.C(n_270),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_308),
.C(n_291),
.Y(n_317)
);

XNOR2x1_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_279),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_309),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_276),
.B(n_280),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_310),
.B(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_268),
.C(n_223),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_287),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_317),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_297),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_316),
.B(n_304),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_288),
.B(n_292),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_291),
.C(n_295),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_312),
.C(n_308),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_324),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_296),
.B1(n_309),
.B2(n_299),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_325),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_304),
.B(n_186),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_317),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_326),
.A2(n_314),
.B(n_5),
.C(n_6),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_4),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_327),
.A2(n_329),
.B(n_323),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_323),
.C(n_321),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_314),
.C(n_5),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

HAxp5_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_5),
.CON(n_336),
.SN(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_264),
.Y(n_337)
);


endmodule