module fake_jpeg_8226_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_50),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_52),
.B1(n_54),
.B2(n_60),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_59),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_25),
.C(n_27),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_19),
.B1(n_17),
.B2(n_16),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_19),
.B1(n_17),
.B2(n_30),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_17),
.B1(n_19),
.B2(n_16),
.Y(n_105)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_75),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_83),
.Y(n_131)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_68),
.B1(n_67),
.B2(n_42),
.Y(n_121)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_21),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_92),
.B(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_90),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_23),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_40),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx11_ASAP7_75t_SL g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_18),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_62),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_101),
.B1(n_105),
.B2(n_17),
.Y(n_113)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_98),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_51),
.B(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_40),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_43),
.B(n_28),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_29),
.B(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_23),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_28),
.B(n_29),
.C(n_32),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_102),
.B1(n_32),
.B2(n_74),
.Y(n_141)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_128),
.Y(n_137)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_136),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_28),
.B(n_29),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_125),
.B(n_126),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_42),
.B1(n_41),
.B2(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_81),
.B1(n_103),
.B2(n_41),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_123),
.B1(n_80),
.B2(n_86),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_94),
.B1(n_74),
.B2(n_72),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_0),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_106),
.Y(n_152)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_72),
.C(n_78),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_143),
.C(n_130),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_78),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_139),
.A2(n_158),
.B(n_44),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_147),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_80),
.B1(n_122),
.B2(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_114),
.B1(n_109),
.B2(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_160),
.B1(n_165),
.B2(n_109),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_83),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_152),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_101),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_80),
.B(n_105),
.Y(n_158)
);

AO21x2_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_75),
.B(n_67),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_114),
.B(n_100),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_82),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_23),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_169),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_117),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_126),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_40),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_171),
.A2(n_174),
.B(n_195),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_133),
.B1(n_125),
.B2(n_130),
.C(n_118),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_180),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_132),
.B(n_42),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_178),
.C(n_183),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_41),
.C(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_185),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_37),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_40),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_193),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_159),
.A3(n_151),
.B1(n_139),
.B2(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_200),
.B(n_159),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_197),
.B1(n_159),
.B2(n_169),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_196),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_18),
.B(n_114),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_40),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_140),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_134),
.B1(n_38),
.B2(n_37),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_139),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_210),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_228),
.B1(n_218),
.B2(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_194),
.B(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_186),
.B(n_178),
.C(n_174),
.D(n_193),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_38),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_218),
.B(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_220),
.A2(n_172),
.B1(n_175),
.B2(n_170),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_223),
.B(n_224),
.C(n_225),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_168),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_160),
.B1(n_200),
.B2(n_201),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_183),
.B1(n_184),
.B2(n_177),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_234),
.A2(n_251),
.B1(n_203),
.B2(n_206),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_247),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_226),
.C(n_229),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_242),
.C(n_244),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_246),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_168),
.C(n_156),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_37),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_157),
.C(n_37),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_37),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_215),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_249),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_38),
.C(n_163),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_176),
.B1(n_134),
.B2(n_129),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_176),
.B1(n_129),
.B2(n_93),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_38),
.C(n_44),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_217),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_216),
.B(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_266),
.B(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_224),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_44),
.B1(n_9),
.B2(n_3),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_217),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_223),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_270),
.B(n_241),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_225),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_221),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_235),
.C(n_247),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_275),
.B(n_267),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_242),
.C(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_284),
.C(n_286),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_262),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_241),
.B(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_280),
.B(n_10),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_10),
.B(n_14),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_38),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_290),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_256),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_276),
.B1(n_275),
.B2(n_279),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_294),
.Y(n_300)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_257),
.C(n_44),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_11),
.B(n_4),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_10),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_1),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_306),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_283),
.B1(n_272),
.B2(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.C(n_293),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_9),
.B(n_15),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_12),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_289),
.B(n_293),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_311),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_315),
.B(n_301),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

AO221x1_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_316),
.B1(n_309),
.B2(n_305),
.C(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_297),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_11),
.C(n_4),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_320),
.A3(n_6),
.B1(n_7),
.B2(n_13),
.C1(n_15),
.C2(n_2),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_12),
.B(n_4),
.Y(n_321)
);

AOI321xp33_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.A3(n_13),
.B1(n_2),
.B2(n_318),
.C(n_44),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_13),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_2),
.Y(n_325)
);


endmodule