module fake_jpeg_12903_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_18),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_21),
.B1(n_15),
.B2(n_12),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_53),
.Y(n_62)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_29),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_58),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_33),
.A3(n_26),
.B1(n_19),
.B2(n_16),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_43),
.B(n_13),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_59),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_13),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_30),
.B1(n_20),
.B2(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_40),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_47),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_78),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_71),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_70),
.B(n_62),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_58),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_88),
.B(n_69),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_66),
.B1(n_70),
.B2(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_66),
.B(n_67),
.C(n_70),
.D(n_72),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_73),
.B(n_69),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_78),
.C(n_76),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_96),
.B(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_0),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_91),
.B1(n_84),
.B2(n_31),
.Y(n_98)
);

AO221x1_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_69),
.B1(n_52),
.B2(n_2),
.C(n_1),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_14),
.C(n_32),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_94),
.C(n_14),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_91),
.B(n_1),
.C(n_0),
.Y(n_100)
);

OAI33xp33_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_0),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.B3(n_9),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

OAI31xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_100),
.A3(n_8),
.B(n_10),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_101),
.B(n_5),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_106),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_108),
.Y(n_111)
);


endmodule