module fake_jpeg_11488_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_57),
.Y(n_69)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_50),
.B1(n_47),
.B2(n_58),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_74),
.B(n_2),
.C(n_4),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_50),
.B1(n_47),
.B2(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_82),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_48),
.B(n_2),
.C(n_3),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_0),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_22),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_25),
.C(n_39),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_5),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_5),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_6),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_93),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_36),
.B1(n_38),
.B2(n_97),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_10),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_11),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_13),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_41),
.B1(n_17),
.B2(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_15),
.B1(n_26),
.B2(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_112),
.A3(n_117),
.B1(n_98),
.B2(n_99),
.C1(n_103),
.C2(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_111),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_96),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_115),
.C(n_116),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_110),
.B1(n_121),
.B2(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_126),
.Y(n_133)
);


endmodule