module fake_jpeg_673_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_53),
.Y(n_82)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_59),
.B1(n_51),
.B2(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_83),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_19),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_61),
.B1(n_54),
.B2(n_49),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_61),
.B(n_54),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_50),
.B1(n_57),
.B2(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_46),
.C(n_47),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_93),
.C(n_6),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_97),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_62),
.C(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_57),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_58),
.A3(n_54),
.B1(n_52),
.B2(n_25),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_0),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_101),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_4),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_2),
.B(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_2),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_115),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_28),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_93),
.C(n_13),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_5),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_41),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_12),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_26),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_115),
.B1(n_112),
.B2(n_113),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_89),
.B1(n_100),
.B2(n_85),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_132),
.B(n_40),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_135),
.B1(n_37),
.B2(n_38),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_43),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_42),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_138),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_103),
.B(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_30),
.C(n_31),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_125),
.C(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_36),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_128),
.B1(n_122),
.B2(n_130),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_145),
.B(n_120),
.Y(n_160)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_156),
.B(n_146),
.CI(n_143),
.CON(n_159),
.SN(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_156),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_158),
.C(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_140),
.C(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_144),
.B(n_147),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_157),
.B(n_153),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_152),
.C(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_144),
.Y(n_169)
);


endmodule