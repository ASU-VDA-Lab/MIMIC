module fake_jpeg_16150_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_11),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_0),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.Y(n_73)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_25),
.B1(n_46),
.B2(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_25),
.B1(n_60),
.B2(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_85),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_48),
.B1(n_52),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_116),
.B1(n_74),
.B2(n_89),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_122),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_62),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_29),
.B(n_58),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_115),
.B(n_28),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_111),
.Y(n_149)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_54),
.Y(n_111)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_121),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_119),
.B1(n_82),
.B2(n_96),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_48),
.B1(n_64),
.B2(n_46),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_65),
.Y(n_136)
);

CKINVDCx12_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_40),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_141),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_77),
.B1(n_32),
.B2(n_92),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_133),
.B1(n_155),
.B2(n_96),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_135),
.A2(n_156),
.B1(n_109),
.B2(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_139),
.Y(n_175)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_125),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_50),
.C(n_49),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_47),
.C(n_49),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_41),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_157),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_100),
.A2(n_33),
.B1(n_40),
.B2(n_24),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_165),
.B1(n_156),
.B2(n_136),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_162),
.Y(n_181)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_33),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_100),
.C(n_47),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_173),
.C(n_144),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_118),
.C(n_66),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_147),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_165),
.C(n_153),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_164),
.B(n_179),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_185),
.B(n_198),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_157),
.B(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_133),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_194),
.B1(n_196),
.B2(n_101),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_195),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_133),
.B1(n_131),
.B2(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_139),
.B1(n_147),
.B2(n_149),
.Y(n_196)
);

MAJx3_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_149),
.C(n_141),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_112),
.B(n_132),
.C(n_125),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_145),
.B(n_137),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_158),
.A2(n_117),
.B1(n_150),
.B2(n_140),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_199),
.A2(n_178),
.B1(n_159),
.B2(n_170),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_172),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_207),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_206),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_150),
.Y(n_207)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_219),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_152),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_152),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_33),
.B1(n_125),
.B2(n_117),
.Y(n_216)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_180),
.C(n_189),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_177),
.B1(n_172),
.B2(n_140),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_220),
.B1(n_222),
.B2(n_225),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_176),
.B1(n_174),
.B2(n_142),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_194),
.A2(n_174),
.B1(n_132),
.B2(n_134),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_148),
.B(n_134),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_201),
.B(n_200),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_226),
.B(n_228),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_197),
.A2(n_162),
.B1(n_143),
.B2(n_97),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_189),
.C(n_199),
.Y(n_226)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_215),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_19),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_248),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_224),
.B(n_216),
.Y(n_261)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_183),
.B1(n_195),
.B2(n_187),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_239),
.B1(n_252),
.B2(n_1),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_166),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_246),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_209),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_23),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_249),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_21),
.B1(n_31),
.B2(n_41),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_212),
.A2(n_151),
.B1(n_97),
.B2(n_34),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_254),
.A2(n_203),
.B1(n_223),
.B2(n_227),
.Y(n_257)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_226),
.B1(n_222),
.B2(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_217),
.C(n_225),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_272),
.C(n_273),
.Y(n_285)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_261),
.B(n_237),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_224),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_266),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

AOI22x1_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_42),
.B1(n_39),
.B2(n_26),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_275),
.B1(n_277),
.B2(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_113),
.C(n_22),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_113),
.C(n_22),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_113),
.C(n_22),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_240),
.C(n_236),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_34),
.B1(n_39),
.B2(n_42),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_251),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_286),
.C(n_292),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_255),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_251),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_290),
.Y(n_308)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.Y(n_298)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_254),
.C(n_244),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_232),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_235),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_271),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_244),
.B1(n_250),
.B2(n_263),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_301),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_284),
.B1(n_292),
.B2(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_250),
.B1(n_263),
.B2(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_274),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_312),
.B(n_287),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_261),
.C(n_267),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_282),
.C(n_26),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_268),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_35),
.Y(n_319)
);

NAND2x1_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_267),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_311),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_4),
.B(n_5),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_5),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_315),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_35),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_42),
.C(n_39),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_319),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_26),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_308),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_310),
.B1(n_298),
.B2(n_297),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_35),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_327),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_306),
.B1(n_307),
.B2(n_304),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_330),
.B(n_333),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_321),
.A2(n_312),
.B(n_7),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_331),
.A2(n_336),
.B(n_10),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_332),
.B(n_317),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_23),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_323),
.C(n_23),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_9),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_324),
.A2(n_8),
.B(n_9),
.Y(n_336)
);

NAND2xp67_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_323),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_337),
.B(n_341),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_344),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_343),
.C(n_334),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_23),
.C(n_22),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_345),
.A2(n_338),
.B(n_12),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_338),
.A2(n_326),
.B(n_330),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_346),
.A2(n_349),
.B(n_14),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_347),
.B(n_348),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_10),
.B(n_13),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_354),
.B(n_350),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_43),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_355),
.A2(n_352),
.B(n_16),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_14),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_357),
.A2(n_14),
.B(n_16),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_18),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_43),
.C(n_356),
.Y(n_360)
);


endmodule