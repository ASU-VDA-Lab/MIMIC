module real_jpeg_18716_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_521),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_0),
.B(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_1),
.B(n_46),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_1),
.B(n_277),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_1),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_1),
.B(n_426),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_1),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_1),
.B(n_490),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_1),
.B(n_496),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_2),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_2),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_2),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_2),
.B(n_141),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g151 ( 
.A(n_2),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_3),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g467 ( 
.A(n_3),
.Y(n_467)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_4),
.Y(n_338)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_4),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_5),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_5),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_5),
.B(n_45),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_5),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_5),
.B(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_5),
.A2(n_12),
.B1(n_298),
.B2(n_302),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_6),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_6),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_6),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_7),
.Y(n_522)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_8),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_8),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_9),
.Y(n_341)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_9),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_10),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_10),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_10),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_10),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_10),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_10),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_10),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_10),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_11),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_11),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_11),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_11),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_11),
.B(n_421),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_11),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_11),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_11),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_12),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_12),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_12),
.B(n_69),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_12),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_12),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_12),
.B(n_482),
.Y(n_481)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_13),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_13),
.Y(n_279)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_14),
.B(n_69),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_14),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_14),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_14),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_14),
.B(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

BUFx4f_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_16),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_16),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_17),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_164),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_163),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_143),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_23),
.B(n_143),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.C(n_104),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_24),
.B(n_80),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_27),
.B(n_42),
.C(n_54),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.C(n_38),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_29),
.B1(n_38),
.B2(n_53),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_28),
.A2(n_29),
.B1(n_94),
.B2(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_28),
.A2(n_29),
.B1(n_286),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_94),
.C(n_99),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_29),
.B(n_286),
.C(n_287),
.Y(n_285)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_31),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_33),
.B(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_36),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_38),
.B(n_117),
.C(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_38),
.A2(n_53),
.B1(n_116),
.B2(n_117),
.Y(n_307)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_48),
.A2(n_52),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_48),
.B(n_53),
.C(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_48),
.A2(n_52),
.B1(n_219),
.B2(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_49),
.Y(n_270)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_52),
.B(n_123),
.C(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_56),
.B(n_72),
.C(n_78),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.C(n_68),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_57),
.A2(n_58),
.B1(n_68),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_62),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_63),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_65),
.Y(n_184)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_67),
.Y(n_199)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_68),
.B(n_192),
.C(n_195),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_68),
.B(n_195),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_72),
.B(n_191),
.C(n_197),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_72),
.A2(n_73),
.B1(n_197),
.B2(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_130),
.C(n_139),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_73),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_76),
.Y(n_259)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.C(n_93),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_81),
.B(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_83),
.B(n_93),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_91),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_89),
.A2(n_123),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_94),
.A2(n_95),
.B1(n_132),
.B2(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_132),
.C(n_135),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_95),
.B(n_239),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_SL g397 ( 
.A(n_95),
.B(n_295),
.Y(n_397)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_97),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_98),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_124),
.C(n_129),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_121),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_106),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_108),
.B(n_121),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_116),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_117),
.B(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_120),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_130),
.A2(n_131),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_182),
.C(n_185),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_132),
.A2(n_133),
.B1(n_185),
.B2(n_186),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_132),
.B(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_133),
.B(n_405),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_134),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_161),
.B2(n_162),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_150),
.B(n_232),
.C(n_242),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_150),
.A2(n_151),
.B1(n_242),
.B2(n_243),
.Y(n_361)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_245),
.B(n_518),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_203),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21x1_ASAP7_75t_SL g518 ( 
.A1(n_168),
.A2(n_519),
.B(n_520),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_169),
.B(n_171),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_174),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_190),
.C(n_200),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_178),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_188),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_179),
.B(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_181),
.B(n_188),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_183),
.B(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_183),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_185),
.A2(n_186),
.B1(n_282),
.B2(n_283),
.Y(n_333)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_186),
.B(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_200),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_217),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_194),
.Y(n_288)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_204),
.B(n_206),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_213),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_207),
.B(n_211),
.Y(n_382)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_213),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_226),
.C(n_230),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_214),
.A2(n_215),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_223),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_216),
.B(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_218),
.B(n_224),
.Y(n_368)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_226),
.A2(n_227),
.B1(n_230),
.B2(n_231),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_232),
.A2(n_233),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_234),
.A2(n_239),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_237),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_239),
.Y(n_295)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_512),
.Y(n_245)
);

NAND4xp25_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_369),
.C(n_383),
.D(n_388),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_346),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_322),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_249),
.B(n_322),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_289),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_250),
.B(n_290),
.C(n_305),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_260),
.B1(n_261),
.B2(n_264),
.Y(n_257)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_258),
.A2(n_261),
.B(n_265),
.C(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_260),
.B(n_264),
.Y(n_363)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_263),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_267),
.B(n_350),
.C(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_280),
.C(n_285),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_268),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_272),
.C(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_284),
.Y(n_505)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_287),
.B(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_305),
.Y(n_289)
);

XOR2x2_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_356),
.C(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_309),
.B(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_SL g483 ( 
.A(n_300),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_315),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_308),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.C(n_320),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_316),
.B(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_317),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.C(n_329),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_323),
.B(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_325),
.A2(n_326),
.B1(n_329),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.C(n_334),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_330),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_334),
.Y(n_393)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.C(n_342),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_335),
.B(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21x1_ASAP7_75t_SL g513 ( 
.A1(n_346),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_347),
.B(n_348),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_353),
.C(n_367),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_366),
.B2(n_367),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_362),
.B1(n_364),
.B2(n_365),
.Y(n_358)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_359),
.Y(n_364)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_362),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_377),
.C(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

A2O1A1O1Ixp25_ASAP7_75t_L g512 ( 
.A1(n_369),
.A2(n_383),
.B(n_513),
.C(n_516),
.D(n_517),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_381),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_370),
.B(n_381),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_375),
.C(n_379),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_372),
.B1(n_379),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_373),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_379),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_384),
.B(n_385),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_413),
.B(n_511),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_410),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_390),
.B(n_410),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.C(n_396),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_391),
.A2(n_392),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_394),
.B(n_396),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.C(n_404),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_397),
.A2(n_398),
.B1(n_399),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_404),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_409),
.Y(n_480)
);

AOI21x1_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_439),
.B(n_510),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_436),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_415),
.B(n_436),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.C(n_434),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_434),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.C(n_431),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_444),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_431),
.Y(n_444)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_458),
.B(n_509),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_456),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_441),
.B(n_456),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.C(n_454),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_442),
.A2(n_443),
.B1(n_469),
.B2(n_471),
.Y(n_468)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_445),
.A2(n_454),
.B1(n_455),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_451),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_446),
.A2(n_447),
.B1(n_451),
.B2(n_452),
.Y(n_461)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_472),
.B(n_508),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_468),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_460),
.B(n_468),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.C(n_466),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_485),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_466),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_469),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_487),
.B(n_507),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_484),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_474),
.B(n_484),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_481),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_481),
.Y(n_493)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_494),
.B(n_506),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_493),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_489),
.B(n_493),
.Y(n_506)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_502),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);


endmodule