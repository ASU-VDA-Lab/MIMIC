module fake_jpeg_25532_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_36),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_19),
.B1(n_14),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_29),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_19),
.B(n_14),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_1),
.B(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_3),
.B1(n_4),
.B2(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_39),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_63),
.Y(n_75)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_45),
.C(n_49),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.C(n_76),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_48),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_57),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_45),
.C(n_40),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_87),
.B(n_54),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_64),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_86),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_59),
.B1(n_51),
.B2(n_48),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_60),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_44),
.B1(n_41),
.B2(n_15),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_76),
.C(n_72),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_93),
.C(n_54),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_71),
.C(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_15),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_82),
.B1(n_93),
.B2(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_54),
.B1(n_4),
.B2(n_3),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_89),
.B(n_80),
.C(n_13),
.D(n_77),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_5),
.Y(n_117)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_13),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_98),
.C(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_114),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_117),
.C(n_109),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_4),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_9),
.B(n_11),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_122),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_12),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_115),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_126),
.A2(n_104),
.B(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_128),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_123),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.C(n_12),
.Y(n_131)
);


endmodule