module real_aes_17460_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_0), .A2(n_4), .B1(n_782), .B2(n_783), .Y(n_781) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_0), .A2(n_212), .B1(n_595), .B2(n_823), .Y(n_822) );
OAI22xp33_ASAP7_75t_SL g374 ( .A1(n_1), .A2(n_118), .B1(n_375), .B2(n_378), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_1), .A2(n_23), .B1(n_412), .B2(n_413), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_2), .A2(n_24), .B1(n_368), .B2(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_2), .A2(n_122), .B1(n_391), .B2(n_412), .Y(n_470) );
INVx1_ASAP7_75t_L g598 ( .A(n_3), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_4), .A2(n_216), .B1(n_823), .B2(n_827), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_5), .A2(n_1284), .B1(n_1285), .B2(n_1286), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1284 ( .A(n_5), .Y(n_1284) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_6), .A2(n_232), .B1(n_522), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_6), .A2(n_161), .B1(n_653), .B2(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_7), .Y(n_461) );
INVx1_ASAP7_75t_L g579 ( .A(n_8), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_9), .A2(n_213), .B1(n_522), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_9), .A2(n_195), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g1263 ( .A(n_10), .Y(n_1263) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_11), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_12), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g345 ( .A(n_12), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_13), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_14), .A2(n_205), .B1(n_518), .B2(n_522), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_14), .A2(n_54), .B1(n_546), .B2(n_549), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_15), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_16), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_17), .A2(n_188), .B1(n_467), .B2(n_679), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_17), .A2(n_188), .B1(n_753), .B2(n_755), .Y(n_752) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_18), .A2(n_191), .B1(n_363), .B2(n_370), .C1(n_487), .C2(n_489), .Y(n_486) );
OAI222xp33_ASAP7_75t_L g529 ( .A1(n_18), .A2(n_136), .B1(n_191), .B2(n_530), .C1(n_532), .C2(n_533), .Y(n_529) );
INVx1_ASAP7_75t_L g800 ( .A(n_19), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_19), .A2(n_37), .B1(n_472), .B2(n_532), .Y(n_812) );
INVx1_ASAP7_75t_L g807 ( .A(n_20), .Y(n_807) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_21), .B(n_1030), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_21), .B(n_102), .Y(n_1032) );
INVx2_ASAP7_75t_L g1036 ( .A(n_21), .Y(n_1036) );
OAI211xp5_ASAP7_75t_L g1289 ( .A1(n_22), .A2(n_724), .B(n_971), .C(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1298 ( .A(n_22), .Y(n_1298) );
OAI22xp33_ASAP7_75t_SL g367 ( .A1(n_23), .A2(n_215), .B1(n_368), .B2(n_371), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_24), .B(n_389), .Y(n_469) );
INVx1_ASAP7_75t_L g1232 ( .A(n_25), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_26), .A2(n_194), .B1(n_412), .B2(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_26), .A2(n_242), .B1(n_368), .B2(n_467), .Y(n_612) );
INVx1_ASAP7_75t_L g1306 ( .A(n_27), .Y(n_1306) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_28), .A2(n_146), .B1(n_378), .B2(n_466), .Y(n_1003) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_28), .A2(n_239), .B1(n_412), .B2(n_413), .Y(n_1005) );
INVx1_ASAP7_75t_L g504 ( .A(n_29), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_29), .A2(n_205), .B1(n_549), .B2(n_563), .Y(n_562) );
XOR2xp5_ASAP7_75t_L g255 ( .A(n_30), .B(n_256), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_31), .A2(n_162), .B1(n_1037), .B2(n_1041), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_32), .A2(n_156), .B1(n_1031), .B2(n_1037), .Y(n_1069) );
INVx1_ASAP7_75t_L g1236 ( .A(n_33), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_34), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_35), .A2(n_181), .B1(n_1027), .B2(n_1034), .Y(n_1084) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_36), .Y(n_442) );
INVx1_ASAP7_75t_L g803 ( .A(n_37), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_38), .A2(n_182), .B1(n_368), .B2(n_796), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_38), .A2(n_94), .B1(n_412), .B2(n_413), .Y(n_969) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_39), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_40), .Y(n_300) );
INVx1_ASAP7_75t_L g1292 ( .A(n_41), .Y(n_1292) );
OAI211xp5_ASAP7_75t_L g1296 ( .A1(n_41), .A2(n_451), .B(n_1272), .C(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g886 ( .A(n_42), .Y(n_886) );
INVx1_ASAP7_75t_L g1231 ( .A(n_43), .Y(n_1231) );
INVx1_ASAP7_75t_L g808 ( .A(n_44), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_45), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_46), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_47), .A2(n_187), .B1(n_1027), .B2(n_1037), .Y(n_1056) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_48), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_49), .A2(n_106), .B1(n_1027), .B2(n_1034), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g1068 ( .A1(n_50), .A2(n_98), .B1(n_1027), .B2(n_1034), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_51), .A2(n_138), .B1(n_532), .B2(n_892), .Y(n_891) );
INVxp67_ASAP7_75t_SL g903 ( .A(n_51), .Y(n_903) );
INVx1_ASAP7_75t_L g840 ( .A(n_52), .Y(n_840) );
INVx1_ASAP7_75t_L g273 ( .A(n_53), .Y(n_273) );
INVx1_ASAP7_75t_L g279 ( .A(n_53), .Y(n_279) );
INVx1_ASAP7_75t_L g508 ( .A(n_54), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_55), .Y(n_429) );
XOR2xp5_ASAP7_75t_L g565 ( .A(n_56), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g716 ( .A(n_57), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_58), .A2(n_76), .B1(n_782), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g821 ( .A(n_58), .Y(n_821) );
INVx1_ASAP7_75t_L g703 ( .A(n_59), .Y(n_703) );
XOR2x2_ASAP7_75t_L g882 ( .A(n_60), .B(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_61), .A2(n_180), .B1(n_639), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_61), .A2(n_186), .B1(n_662), .B2(n_666), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_62), .A2(n_77), .B1(n_522), .B2(n_659), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g926 ( .A1(n_62), .A2(n_220), .B1(n_827), .B2(n_927), .Y(n_926) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_63), .A2(n_349), .B(n_962), .C(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g973 ( .A(n_63), .Y(n_973) );
INVx2_ASAP7_75t_L g266 ( .A(n_64), .Y(n_266) );
INVx1_ASAP7_75t_L g571 ( .A(n_65), .Y(n_571) );
XNOR2x2_ASAP7_75t_L g692 ( .A(n_66), .B(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_66), .A2(n_88), .B1(n_1034), .B2(n_1041), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_67), .A2(n_200), .B1(n_682), .B2(n_748), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_67), .A2(n_200), .B1(n_764), .B2(n_765), .Y(n_763) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_68), .Y(n_889) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_68), .A2(n_138), .B1(n_684), .B2(n_688), .Y(n_904) );
INVx1_ASAP7_75t_L g1014 ( .A(n_69), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_70), .A2(n_133), .B1(n_1266), .B2(n_1267), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1275 ( .A1(n_70), .A2(n_133), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
INVx1_ASAP7_75t_L g1315 ( .A(n_71), .Y(n_1315) );
OAI222xp33_ASAP7_75t_L g628 ( .A1(n_72), .A2(n_104), .B1(n_211), .B2(n_393), .C1(n_629), .C2(n_630), .Y(n_628) );
OAI222xp33_ASAP7_75t_L g683 ( .A1(n_72), .A2(n_104), .B1(n_211), .B2(n_684), .C1(n_685), .C2(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g705 ( .A(n_73), .Y(n_705) );
INVx1_ASAP7_75t_L g794 ( .A(n_74), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_75), .A2(n_94), .B1(n_375), .B2(n_378), .Y(n_967) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_75), .A2(n_182), .B1(n_389), .B2(n_391), .Y(n_974) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_76), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_77), .A2(n_87), .B1(n_827), .B2(n_877), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_78), .A2(n_125), .B1(n_1258), .B2(n_1260), .Y(n_1257) );
OAI22xp33_ASAP7_75t_L g1269 ( .A1(n_78), .A2(n_125), .B1(n_481), .B2(n_1270), .Y(n_1269) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_79), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_80), .A2(n_246), .B1(n_645), .B2(n_647), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_80), .A2(n_128), .B1(n_673), .B2(n_674), .Y(n_672) );
XOR2xp5_ASAP7_75t_L g477 ( .A(n_81), .B(n_478), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_81), .A2(n_123), .B1(n_1027), .B2(n_1034), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_82), .A2(n_128), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_82), .A2(n_246), .B1(n_662), .B2(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g357 ( .A(n_83), .Y(n_357) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_83), .A2(n_393), .B(n_398), .C(n_408), .Y(n_392) );
INVx1_ASAP7_75t_L g845 ( .A(n_84), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_84), .A2(n_219), .B1(n_275), .B2(n_630), .C(n_851), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_85), .A2(n_145), .B1(n_458), .B2(n_466), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_85), .A2(n_145), .B1(n_389), .B2(n_391), .Y(n_849) );
INVx1_ASAP7_75t_L g801 ( .A(n_86), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_87), .A2(n_220), .B1(n_513), .B2(n_913), .Y(n_917) );
INVx1_ASAP7_75t_L g698 ( .A(n_89), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g737 ( .A1(n_90), .A2(n_738), .B(n_741), .C(n_746), .Y(n_737) );
INVx1_ASAP7_75t_L g762 ( .A(n_90), .Y(n_762) );
INVx1_ASAP7_75t_L g932 ( .A(n_91), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g1054 ( .A1(n_91), .A2(n_121), .B1(n_1027), .B2(n_1034), .Y(n_1054) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_92), .A2(n_242), .B1(n_389), .B2(n_413), .C(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g610 ( .A(n_92), .Y(n_610) );
AOI22xp5_ASAP7_75t_SL g1053 ( .A1(n_93), .A2(n_235), .B1(n_1037), .B2(n_1041), .Y(n_1053) );
OAI211xp5_ASAP7_75t_L g480 ( .A1(n_95), .A2(n_481), .B(n_482), .C(n_493), .Y(n_480) );
INVx1_ASAP7_75t_L g537 ( .A(n_95), .Y(n_537) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_96), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_96), .B(n_1014), .Y(n_1028) );
INVx1_ASAP7_75t_L g573 ( .A(n_97), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_99), .A2(n_195), .B1(n_484), .B2(n_859), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_99), .A2(n_213), .B1(n_867), .B2(n_869), .Y(n_866) );
INVx1_ASAP7_75t_L g1313 ( .A(n_100), .Y(n_1313) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_101), .A2(n_109), .B1(n_1031), .B2(n_1037), .Y(n_1065) );
INVx1_ASAP7_75t_L g1030 ( .A(n_102), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_102), .B(n_1036), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_103), .A2(n_243), .B1(n_1027), .B2(n_1031), .Y(n_1026) );
INVx1_ASAP7_75t_L g574 ( .A(n_105), .Y(n_574) );
INVx1_ASAP7_75t_L g894 ( .A(n_107), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g987 ( .A(n_108), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_110), .A2(n_203), .B1(n_600), .B2(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_110), .A2(n_203), .B1(n_371), .B2(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g265 ( .A(n_111), .Y(n_265) );
INVx1_ASAP7_75t_L g309 ( .A(n_111), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_112), .Y(n_938) );
INVx1_ASAP7_75t_L g1309 ( .A(n_113), .Y(n_1309) );
AOI22xp33_ASAP7_75t_SL g918 ( .A1(n_114), .A2(n_234), .B1(n_522), .B2(n_659), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_114), .A2(n_167), .B1(n_544), .B2(n_921), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_115), .A2(n_209), .B1(n_1027), .B2(n_1034), .Y(n_1042) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_116), .Y(n_941) );
INVx1_ASAP7_75t_L g1238 ( .A(n_117), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_118), .A2(n_215), .B1(n_389), .B2(n_391), .Y(n_388) );
OAI22xp33_ASAP7_75t_SL g465 ( .A1(n_119), .A2(n_122), .B1(n_466), .B2(n_467), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_119), .A2(n_126), .B1(n_403), .B2(n_404), .Y(n_474) );
INVx1_ASAP7_75t_L g621 ( .A(n_120), .Y(n_621) );
INVx1_ASAP7_75t_L g1264 ( .A(n_124), .Y(n_1264) );
OAI211xp5_ASAP7_75t_L g1271 ( .A1(n_124), .A2(n_451), .B(n_1272), .C(n_1273), .Y(n_1271) );
INVx1_ASAP7_75t_L g463 ( .A(n_126), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g1293 ( .A1(n_127), .A2(n_210), .B1(n_412), .B2(n_1294), .Y(n_1293) );
OAI22xp33_ASAP7_75t_L g1302 ( .A1(n_127), .A2(n_210), .B1(n_368), .B2(n_378), .Y(n_1302) );
XOR2xp5_ASAP7_75t_L g617 ( .A(n_129), .B(n_618), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_130), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_131), .A2(n_226), .B1(n_1037), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1241 ( .A(n_132), .Y(n_1241) );
INVx1_ASAP7_75t_L g1321 ( .A(n_134), .Y(n_1321) );
INVx1_ASAP7_75t_L g492 ( .A(n_135), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_135), .A2(n_199), .B1(n_389), .B2(n_391), .Y(n_534) );
INVx1_ASAP7_75t_L g483 ( .A(n_136), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_137), .Y(n_510) );
BUFx3_ASAP7_75t_L g271 ( .A(n_139), .Y(n_271) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_140), .A2(n_348), .B(n_349), .C(n_460), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g471 ( .A1(n_140), .A2(n_408), .B(n_472), .C(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g780 ( .A(n_141), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_142), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_143), .Y(n_991) );
INVx1_ASAP7_75t_L g700 ( .A(n_144), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g1009 ( .A1(n_146), .A2(n_244), .B1(n_389), .B2(n_391), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g988 ( .A(n_147), .Y(n_988) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_148), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_149), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_150), .Y(n_499) );
INVx1_ASAP7_75t_L g597 ( .A(n_151), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_152), .A2(n_186), .B1(n_639), .B2(n_642), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_152), .A2(n_180), .B1(n_659), .B2(n_660), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g980 ( .A(n_153), .Y(n_980) );
INVx1_ASAP7_75t_L g1318 ( .A(n_154), .Y(n_1318) );
INVx1_ASAP7_75t_L g712 ( .A(n_155), .Y(n_712) );
INVx1_ASAP7_75t_L g1322 ( .A(n_157), .Y(n_1322) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_158), .Y(n_282) );
INVx1_ASAP7_75t_L g797 ( .A(n_159), .Y(n_797) );
INVx1_ASAP7_75t_L g582 ( .A(n_160), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_161), .A2(n_222), .B1(n_804), .B2(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g497 ( .A(n_163), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_163), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_164), .A2(n_170), .B1(n_1031), .B2(n_1037), .Y(n_1083) );
AOI222xp33_ASAP7_75t_L g1223 ( .A1(n_164), .A2(n_1224), .B1(n_1278), .B2(n_1282), .C1(n_1332), .C2(n_1334), .Y(n_1223) );
XOR2xp5_ASAP7_75t_L g1225 ( .A(n_164), .B(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g887 ( .A(n_165), .Y(n_887) );
INVx1_ASAP7_75t_L g1235 ( .A(n_166), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_167), .A2(n_175), .B1(n_910), .B2(n_913), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g1288 ( .A1(n_168), .A2(n_177), .B1(n_389), .B2(n_765), .Y(n_1288) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_168), .A2(n_177), .B1(n_375), .B2(n_1301), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_169), .B(n_396), .Y(n_596) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_169), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_171), .Y(n_304) );
INVx1_ASAP7_75t_L g839 ( .A(n_172), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_173), .Y(n_984) );
OAI211xp5_ASAP7_75t_L g347 ( .A1(n_174), .A2(n_348), .B(n_349), .C(n_356), .Y(n_347) );
INVx1_ASAP7_75t_L g407 ( .A(n_174), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_175), .A2(n_234), .B1(n_544), .B2(n_921), .Y(n_920) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_176), .Y(n_940) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_178), .Y(n_321) );
INVx1_ASAP7_75t_L g844 ( .A(n_179), .Y(n_844) );
INVx1_ASAP7_75t_L g1001 ( .A(n_183), .Y(n_1001) );
OAI211xp5_ASAP7_75t_L g1006 ( .A1(n_183), .A2(n_732), .B(n_971), .C(n_1007), .Y(n_1006) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_184), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_185), .Y(n_937) );
INVx1_ASAP7_75t_L g1319 ( .A(n_189), .Y(n_1319) );
INVx1_ASAP7_75t_L g577 ( .A(n_190), .Y(n_577) );
INVx1_ASAP7_75t_L g745 ( .A(n_192), .Y(n_745) );
OAI211xp5_ASAP7_75t_L g756 ( .A1(n_192), .A2(n_408), .B(n_757), .C(n_758), .Y(n_756) );
OA22x2_ASAP7_75t_L g835 ( .A1(n_193), .A2(n_836), .B1(n_880), .B2(n_881), .Y(n_835) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_193), .Y(n_881) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_194), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_196), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_197), .Y(n_443) );
XOR2xp5_ASAP7_75t_L g421 ( .A(n_198), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g494 ( .A(n_199), .Y(n_494) );
BUFx3_ASAP7_75t_L g315 ( .A(n_201), .Y(n_315) );
INVx1_ASAP7_75t_L g377 ( .A(n_201), .Y(n_377) );
INVx1_ASAP7_75t_L g743 ( .A(n_202), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_204), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_206), .Y(n_431) );
INVx1_ASAP7_75t_L g570 ( .A(n_207), .Y(n_570) );
OAI211xp5_ASAP7_75t_L g998 ( .A1(n_208), .A2(n_349), .B(n_962), .C(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1008 ( .A(n_208), .Y(n_1008) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_212), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_214), .Y(n_946) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_216), .Y(n_786) );
INVx1_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
INVx2_ASAP7_75t_L g307 ( .A(n_217), .Y(n_307) );
INVx1_ASAP7_75t_L g557 ( .A(n_217), .Y(n_557) );
INVx1_ASAP7_75t_L g779 ( .A(n_218), .Y(n_779) );
OAI211xp5_ASAP7_75t_L g842 ( .A1(n_219), .A2(n_503), .B(n_805), .C(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g1291 ( .A(n_221), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_222), .A2(n_232), .B1(n_871), .B2(n_872), .Y(n_870) );
INVx1_ASAP7_75t_L g1243 ( .A(n_223), .Y(n_1243) );
OAI211xp5_ASAP7_75t_L g1261 ( .A1(n_224), .A2(n_629), .B(n_971), .C(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1274 ( .A(n_224), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_225), .A2(n_229), .B1(n_1034), .B2(n_1037), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_227), .Y(n_296) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_228), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g1239 ( .A(n_230), .Y(n_1239) );
INVx1_ASAP7_75t_L g581 ( .A(n_231), .Y(n_581) );
INVx1_ASAP7_75t_L g717 ( .A(n_233), .Y(n_717) );
INVx1_ASAP7_75t_L g896 ( .A(n_236), .Y(n_896) );
AOI21xp33_ASAP7_75t_L g512 ( .A1(n_237), .A2(n_513), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g542 ( .A(n_237), .Y(n_542) );
XNOR2xp5_ASAP7_75t_L g975 ( .A(n_238), .B(n_976), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g1002 ( .A1(n_239), .A2(n_244), .B1(n_368), .B2(n_796), .Y(n_1002) );
INVx1_ASAP7_75t_L g623 ( .A(n_240), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_241), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_245), .Y(n_490) );
INVx1_ASAP7_75t_L g710 ( .A(n_247), .Y(n_710) );
INVx1_ASAP7_75t_L g965 ( .A(n_248), .Y(n_965) );
OAI211xp5_ASAP7_75t_L g970 ( .A1(n_248), .A2(n_732), .B(n_971), .C(n_972), .Y(n_970) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_1011), .B(n_1019), .Y(n_249) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_772), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_613), .B1(n_770), .B2(n_771), .Y(n_251) );
INVx1_ASAP7_75t_L g770 ( .A(n_252), .Y(n_770) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
XNOR2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_476), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_421), .Y(n_254) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_346), .C(n_387), .Y(n_256) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_258), .B(n_311), .Y(n_257) );
OAI33xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_267), .A3(n_281), .B1(n_293), .B2(n_301), .B3(n_305), .Y(n_258) );
OAI33xp33_ASAP7_75t_L g424 ( .A1(n_259), .A2(n_305), .A3(n_425), .B1(n_430), .B2(n_436), .B3(n_441), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g935 ( .A1(n_259), .A2(n_305), .A3(n_936), .B1(n_939), .B2(n_942), .B3(n_947), .Y(n_935) );
OAI33xp33_ASAP7_75t_L g992 ( .A1(n_259), .A2(n_305), .A3(n_993), .B1(n_994), .B2(n_995), .B3(n_996), .Y(n_992) );
BUFx3_ASAP7_75t_L g1229 ( .A(n_259), .Y(n_1229) );
BUFx4f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g540 ( .A(n_260), .Y(n_540) );
BUFx4f_ASAP7_75t_L g719 ( .A(n_260), .Y(n_719) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
AND2x2_ASAP7_75t_SL g343 ( .A(n_261), .B(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_261), .Y(n_420) );
INVx1_ASAP7_75t_L g671 ( .A(n_261), .Y(n_671) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g386 ( .A(n_262), .Y(n_386) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp33_ASAP7_75t_SL g264 ( .A(n_265), .B(n_266), .Y(n_264) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_265), .Y(n_418) );
AND3x4_ASAP7_75t_L g636 ( .A(n_265), .B(n_396), .C(n_637), .Y(n_636) );
INVx3_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
BUFx3_ASAP7_75t_L g396 ( .A(n_266), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B1(n_274), .B2(n_275), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_268), .A2(n_302), .B1(n_317), .B2(n_323), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g301 ( .A1(n_269), .A2(n_302), .B1(n_303), .B2(n_304), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_269), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_269), .A2(n_303), .B1(n_442), .B2(n_443), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_269), .A2(n_530), .B1(n_570), .B2(n_571), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_269), .A2(n_275), .B1(n_581), .B2(n_582), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_269), .A2(n_427), .B1(n_937), .B2(n_938), .Y(n_936) );
BUFx4f_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x4_ASAP7_75t_L g389 ( .A(n_270), .B(n_390), .Y(n_389) );
OR2x4_ASAP7_75t_L g412 ( .A(n_270), .B(n_310), .Y(n_412) );
BUFx3_ASAP7_75t_L g723 ( .A(n_270), .Y(n_723) );
INVx2_ASAP7_75t_L g949 ( .A(n_270), .Y(n_949) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_271), .Y(n_280) );
INVx2_ASAP7_75t_L g287 ( .A(n_271), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_271), .B(n_279), .Y(n_291) );
AND2x4_ASAP7_75t_L g410 ( .A(n_271), .B(n_402), .Y(n_410) );
INVx1_ASAP7_75t_L g548 ( .A(n_272), .Y(n_548) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g286 ( .A(n_273), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_274), .A2(n_304), .B1(n_329), .B2(n_333), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_275), .A2(n_948), .B1(n_980), .B2(n_987), .Y(n_993) );
HB1xp67_ASAP7_75t_L g1242 ( .A(n_275), .Y(n_1242) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g428 ( .A(n_276), .Y(n_428) );
INVx4_ASAP7_75t_L g531 ( .A(n_276), .Y(n_531) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx3_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
BUFx2_ASAP7_75t_L g734 ( .A(n_277), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
BUFx2_ASAP7_75t_L g406 ( .A(n_278), .Y(n_406) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g402 ( .A(n_279), .Y(n_402) );
BUFx2_ASAP7_75t_L g397 ( .A(n_280), .Y(n_397) );
INVx2_ASAP7_75t_L g404 ( .A(n_280), .Y(n_404) );
AND2x4_ASAP7_75t_L g552 ( .A(n_280), .B(n_401), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_288), .B2(n_292), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_282), .A2(n_296), .B1(n_329), .B2(n_333), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g1237 ( .A1(n_283), .A2(n_578), .B1(n_1238), .B2(n_1239), .Y(n_1237) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g576 ( .A(n_284), .Y(n_576) );
INVx2_ASAP7_75t_SL g1317 ( .A(n_284), .Y(n_1317) );
BUFx8_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_285), .Y(n_295) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_285), .Y(n_415) );
INVx2_ASAP7_75t_L g560 ( .A(n_285), .Y(n_560) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x4_ASAP7_75t_L g547 ( .A(n_287), .B(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_288), .A2(n_943), .B1(n_944), .B2(n_946), .Y(n_942) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x6_ASAP7_75t_L g391 ( .A(n_290), .B(n_310), .Y(n_391) );
BUFx3_ASAP7_75t_L g729 ( .A(n_290), .Y(n_729) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g299 ( .A(n_291), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_292), .A2(n_300), .B1(n_323), .B2(n_339), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_296), .B1(n_297), .B2(n_300), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_SL g438 ( .A(n_295), .Y(n_438) );
INVx5_ASAP7_75t_L g727 ( .A(n_295), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_297), .A2(n_559), .B1(n_573), .B2(n_574), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_297), .A2(n_1317), .B1(n_1318), .B2(n_1319), .Y(n_1316) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_299), .Y(n_435) );
INVx2_ASAP7_75t_L g725 ( .A(n_303), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_303), .A2(n_948), .B1(n_950), .B2(n_951), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_303), .A2(n_948), .B1(n_982), .B2(n_988), .Y(n_996) );
OAI22xp33_ASAP7_75t_L g1320 ( .A1(n_303), .A2(n_1308), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
AND2x4_ASAP7_75t_L g313 ( .A(n_306), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g525 ( .A(n_306), .Y(n_525) );
OR2x6_ASAP7_75t_L g583 ( .A(n_306), .B(n_308), .Y(n_583) );
BUFx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g637 ( .A(n_307), .Y(n_637) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND3x1_ASAP7_75t_L g555 ( .A(n_309), .B(n_310), .C(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g390 ( .A(n_310), .Y(n_390) );
AND2x4_ASAP7_75t_L g409 ( .A(n_310), .B(n_410), .Y(n_409) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .A3(n_328), .B1(n_337), .B2(n_338), .B3(n_342), .Y(n_311) );
OAI33xp33_ASAP7_75t_L g584 ( .A1(n_312), .A2(n_342), .A3(n_585), .B1(n_586), .B2(n_587), .B3(n_590), .Y(n_584) );
OAI33xp33_ASAP7_75t_L g952 ( .A1(n_312), .A2(n_953), .A3(n_954), .B1(n_956), .B2(n_958), .B3(n_959), .Y(n_952) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g445 ( .A(n_313), .Y(n_445) );
INVx2_ASAP7_75t_L g696 ( .A(n_313), .Y(n_696) );
INVx4_ASAP7_75t_L g855 ( .A(n_313), .Y(n_855) );
AND2x4_ASAP7_75t_L g344 ( .A(n_315), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
BUFx2_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
AND2x4_ASAP7_75t_L g364 ( .A(n_315), .B(n_365), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_317), .A2(n_448), .B1(n_937), .B2(n_950), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_317), .A2(n_323), .B1(n_941), .B2(n_946), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_317), .A2(n_980), .B1(n_981), .B2(n_982), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_317), .A2(n_448), .B1(n_990), .B2(n_991), .Y(n_989) );
INVx4_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx3_ASAP7_75t_L g699 ( .A(n_318), .Y(n_699) );
BUFx6f_ASAP7_75t_L g1247 ( .A(n_318), .Y(n_1247) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
INVx3_ASAP7_75t_L g370 ( .A(n_319), .Y(n_370) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g327 ( .A(n_321), .Y(n_327) );
INVx2_ASAP7_75t_L g332 ( .A(n_321), .Y(n_332) );
NAND2x1_ASAP7_75t_L g336 ( .A(n_321), .B(n_322), .Y(n_336) );
AND2x2_ASAP7_75t_L g355 ( .A(n_321), .B(n_322), .Y(n_355) );
INVx1_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
AND2x2_ASAP7_75t_L g380 ( .A(n_321), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_322), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
INVx2_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
INVx1_ASAP7_75t_L g521 ( .A(n_322), .Y(n_521) );
AND2x2_ASAP7_75t_L g523 ( .A(n_322), .B(n_327), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_323), .A2(n_433), .B1(n_439), .B2(n_447), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_323), .A2(n_447), .B1(n_570), .B2(n_581), .Y(n_585) );
INVx4_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g449 ( .A(n_324), .Y(n_449) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_324), .Y(n_501) );
INVx2_ASAP7_75t_SL g981 ( .A(n_324), .Y(n_981) );
INVx1_ASAP7_75t_L g1249 ( .A(n_324), .Y(n_1249) );
INVx8_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g373 ( .A(n_325), .B(n_359), .Y(n_373) );
OR2x2_ASAP7_75t_L g458 ( .A(n_325), .B(n_351), .Y(n_458) );
BUFx2_ASAP7_75t_L g1327 ( .A(n_325), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_329), .A2(n_431), .B1(n_437), .B2(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g588 ( .A(n_330), .Y(n_588) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g453 ( .A(n_331), .Y(n_453) );
INVx2_ASAP7_75t_L g507 ( .A(n_331), .Y(n_507) );
BUFx2_ASAP7_75t_L g709 ( .A(n_331), .Y(n_709) );
BUFx2_ASAP7_75t_L g957 ( .A(n_331), .Y(n_957) );
AND2x2_ASAP7_75t_L g520 ( .A(n_332), .B(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_333), .A2(n_940), .B1(n_943), .B2(n_955), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_333), .A2(n_955), .B1(n_1235), .B2(n_1238), .Y(n_1250) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g454 ( .A(n_334), .Y(n_454) );
INVx1_ASAP7_75t_L g503 ( .A(n_334), .Y(n_503) );
INVx1_ASAP7_75t_L g962 ( .A(n_334), .Y(n_962) );
INVx4_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx4f_ASAP7_75t_L g348 ( .A(n_335), .Y(n_348) );
BUFx4f_ASAP7_75t_L g451 ( .A(n_335), .Y(n_451) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_335), .Y(n_511) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_335), .Y(n_589) );
BUFx4f_ASAP7_75t_L g740 ( .A(n_335), .Y(n_740) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g687 ( .A(n_336), .Y(n_687) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x6_ASAP7_75t_L g375 ( .A(n_341), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g466 ( .A(n_341), .B(n_376), .Y(n_466) );
BUFx4f_ASAP7_75t_L g498 ( .A(n_341), .Y(n_498) );
OR2x6_ASAP7_75t_L g679 ( .A(n_341), .B(n_369), .Y(n_679) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_342), .A2(n_445), .A3(n_446), .B1(n_450), .B2(n_452), .B3(n_455), .Y(n_444) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI33xp33_ASAP7_75t_L g853 ( .A1(n_343), .A2(n_854), .A3(n_856), .B1(n_858), .B2(n_861), .B3(n_862), .Y(n_853) );
INVx2_ASAP7_75t_L g959 ( .A(n_343), .Y(n_959) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_344), .A2(n_503), .B1(n_504), .B2(n_505), .C(n_508), .Y(n_502) );
AND2x4_ASAP7_75t_L g669 ( .A(n_344), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_344), .B(n_670), .Y(n_791) );
INVx1_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
AND2x4_ASAP7_75t_L g516 ( .A(n_345), .B(n_352), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_367), .A3(n_374), .B(n_382), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_348), .A2(n_453), .B1(n_573), .B2(n_577), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g603 ( .A(n_349), .B(n_604), .C(n_606), .Y(n_603) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g805 ( .A(n_350), .Y(n_805) );
AOI211xp5_ASAP7_75t_L g901 ( .A1(n_350), .A2(n_902), .B(n_903), .C(n_904), .Y(n_901) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
AND2x2_ASAP7_75t_L g488 ( .A(n_351), .B(n_360), .Y(n_488) );
AND2x2_ASAP7_75t_L g689 ( .A(n_351), .B(n_485), .Y(n_689) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_L g369 ( .A(n_352), .Y(n_369) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g667 ( .A(n_354), .Y(n_667) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_355), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_361), .B2(n_362), .Y(n_356) );
AOI222xp33_ASAP7_75t_L g604 ( .A1(n_358), .A2(n_464), .B1(n_484), .B2(n_597), .C1(n_598), .C2(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_358), .A2(n_1291), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x4_ASAP7_75t_L g462 ( .A(n_359), .B(n_360), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_359), .A2(n_483), .B(n_484), .C(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g491 ( .A(n_359), .Y(n_491) );
AND2x2_ASAP7_75t_L g608 ( .A(n_359), .B(n_609), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g398 ( .A1(n_361), .A2(n_399), .A3(n_403), .B1(n_405), .B2(n_407), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_362), .A2(n_488), .B1(n_800), .B2(n_801), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_362), .A2(n_488), .B1(n_844), .B2(n_845), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_362), .A2(n_488), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_362), .A2(n_742), .B1(n_1263), .B2(n_1274), .Y(n_1273) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g464 ( .A(n_364), .Y(n_464) );
INVx2_ASAP7_75t_L g688 ( .A(n_364), .Y(n_688) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g900 ( .A(n_368), .Y(n_900) );
OR2x6_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_369), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
BUFx3_ASAP7_75t_L g447 ( .A(n_370), .Y(n_447) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_370), .Y(n_591) );
BUFx3_ASAP7_75t_L g715 ( .A(n_370), .Y(n_715) );
INVx2_ASAP7_75t_SL g1326 ( .A(n_370), .Y(n_1326) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_372), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g749 ( .A(n_373), .Y(n_749) );
BUFx2_ASAP7_75t_L g796 ( .A(n_373), .Y(n_796) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_375), .Y(n_682) );
HB1xp67_ASAP7_75t_L g1276 ( .A(n_375), .Y(n_1276) );
AND2x4_ASAP7_75t_L g379 ( .A(n_376), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
CKINVDCx16_ASAP7_75t_R g378 ( .A(n_379), .Y(n_378) );
INVx4_ASAP7_75t_L g467 ( .A(n_379), .Y(n_467) );
INVx3_ASAP7_75t_SL g481 ( .A(n_379), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_379), .A2(n_621), .B1(n_623), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_379), .A2(n_678), .B1(n_807), .B2(n_808), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_379), .A2(n_678), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_379), .A2(n_886), .B1(n_887), .B2(n_900), .Y(n_899) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_380), .Y(n_514) );
INVx2_ASAP7_75t_L g665 ( .A(n_380), .Y(n_665) );
BUFx3_ASAP7_75t_L g912 ( .A(n_380), .Y(n_912) );
OAI31xp33_ASAP7_75t_L g960 ( .A1(n_382), .A2(n_961), .A3(n_966), .B(n_967), .Y(n_960) );
OAI31xp33_ASAP7_75t_L g997 ( .A1(n_382), .A2(n_998), .A3(n_1002), .B(n_1003), .Y(n_997) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI31xp33_ASAP7_75t_L g456 ( .A1(n_383), .A2(n_457), .A3(n_459), .B(n_465), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_383), .A2(n_603), .B(n_612), .Y(n_602) );
INVx1_ASAP7_75t_L g690 ( .A(n_383), .Y(n_690) );
BUFx3_ASAP7_75t_L g750 ( .A(n_383), .Y(n_750) );
BUFx2_ASAP7_75t_SL g906 ( .A(n_383), .Y(n_906) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI21xp5_ASAP7_75t_SL g479 ( .A1(n_384), .A2(n_480), .B(n_495), .Y(n_479) );
INVx1_ASAP7_75t_L g1018 ( .A(n_384), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_384), .B(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI31xp33_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_392), .A3(n_411), .B(n_416), .Y(n_387) );
BUFx2_ASAP7_75t_L g627 ( .A(n_389), .Y(n_627) );
BUFx3_ASAP7_75t_L g764 ( .A(n_389), .Y(n_764) );
INVx2_ASAP7_75t_SL g895 ( .A(n_389), .Y(n_895) );
AND2x2_ASAP7_75t_L g414 ( .A(n_390), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g624 ( .A(n_390), .B(n_415), .Y(n_624) );
INVx2_ASAP7_75t_L g601 ( .A(n_391), .Y(n_601) );
INVx1_ASAP7_75t_L g766 ( .A(n_391), .Y(n_766) );
INVx1_ASAP7_75t_L g897 ( .A(n_391), .Y(n_897) );
BUFx3_ASAP7_75t_L g1267 ( .A(n_391), .Y(n_1267) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_394), .A2(n_631), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_394), .A2(n_631), .B1(n_1291), .B2(n_1292), .Y(n_1290) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
AND2x2_ASAP7_75t_L g405 ( .A(n_395), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g475 ( .A(n_395), .B(n_397), .Y(n_475) );
AND2x4_ASAP7_75t_L g631 ( .A(n_395), .B(n_406), .Y(n_631) );
AND2x2_ASAP7_75t_L g760 ( .A(n_395), .B(n_397), .Y(n_760) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g399 ( .A(n_396), .B(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_399), .A2(n_461), .B1(n_474), .B2(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g472 ( .A(n_405), .Y(n_472) );
INVxp67_ASAP7_75t_L g533 ( .A(n_405), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g594 ( .A1(n_405), .A2(n_475), .B1(n_595), .B2(n_596), .C1(n_597), .C2(n_598), .Y(n_594) );
INVx1_ASAP7_75t_L g892 ( .A(n_405), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_405), .A2(n_475), .B1(n_964), .B2(n_973), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_405), .A2(n_475), .B1(n_1000), .B2(n_1008), .Y(n_1007) );
CKINVDCx8_ASAP7_75t_R g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_409), .B(n_529), .C(n_534), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_409), .B(n_626), .C(n_628), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g810 ( .A1(n_409), .A2(n_801), .B(n_811), .C(n_812), .Y(n_810) );
NOR3xp33_ASAP7_75t_L g848 ( .A(n_409), .B(n_849), .C(n_850), .Y(n_848) );
AOI211xp5_ASAP7_75t_L g888 ( .A1(n_409), .A2(n_889), .B(n_890), .C(n_891), .Y(n_888) );
CKINVDCx8_ASAP7_75t_R g971 ( .A(n_409), .Y(n_971) );
BUFx2_ASAP7_75t_L g549 ( .A(n_410), .Y(n_549) );
BUFx2_ASAP7_75t_L g595 ( .A(n_410), .Y(n_595) );
INVx2_ASAP7_75t_L g643 ( .A(n_410), .Y(n_643) );
BUFx3_ASAP7_75t_L g827 ( .A(n_410), .Y(n_827) );
BUFx2_ASAP7_75t_L g878 ( .A(n_410), .Y(n_878) );
BUFx2_ASAP7_75t_L g890 ( .A(n_410), .Y(n_890) );
INVx1_ASAP7_75t_L g536 ( .A(n_412), .Y(n_536) );
INVx2_ASAP7_75t_SL g622 ( .A(n_412), .Y(n_622) );
INVx2_ASAP7_75t_SL g754 ( .A(n_412), .Y(n_754) );
INVx1_ASAP7_75t_L g1259 ( .A(n_412), .Y(n_1259) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_414), .A2(n_490), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g432 ( .A(n_415), .Y(n_432) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_415), .Y(n_544) );
INVx2_ASAP7_75t_L g820 ( .A(n_415), .Y(n_820) );
INVx1_ASAP7_75t_L g875 ( .A(n_415), .Y(n_875) );
OAI31xp33_ASAP7_75t_SL g468 ( .A1(n_416), .A2(n_469), .A3(n_470), .B(n_471), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_416), .A2(n_593), .B(n_599), .Y(n_592) );
OAI31xp33_ASAP7_75t_SL g968 ( .A1(n_416), .A2(n_969), .A3(n_970), .B(n_974), .Y(n_968) );
OAI31xp33_ASAP7_75t_SL g1004 ( .A1(n_416), .A2(n_1005), .A3(n_1006), .B(n_1009), .Y(n_1004) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_SL g538 ( .A(n_417), .B(n_419), .Y(n_538) );
AND2x4_ASAP7_75t_L g633 ( .A(n_417), .B(n_419), .Y(n_633) );
AND2x2_ASAP7_75t_L g817 ( .A(n_417), .B(n_419), .Y(n_817) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_456), .C(n_468), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g423 ( .A(n_424), .B(n_444), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_426), .A2(n_442), .B1(n_447), .B2(n_448), .Y(n_446) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g1233 ( .A(n_428), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_429), .A2(n_443), .B1(n_453), .B2(n_454), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g824 ( .A1(n_432), .A2(n_440), .B1(n_780), .B2(n_825), .C(n_826), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_432), .A2(n_434), .B1(n_940), .B2(n_941), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_432), .A2(n_434), .B1(n_984), .B2(n_990), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_434), .A2(n_559), .B1(n_1235), .B2(n_1236), .Y(n_1234) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g440 ( .A(n_435), .Y(n_440) );
CKINVDCx8_ASAP7_75t_R g561 ( .A(n_435), .Y(n_561) );
INVx3_ASAP7_75t_L g578 ( .A(n_435), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_438), .A2(n_705), .B1(n_717), .B2(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_438), .A2(n_578), .B1(n_985), .B2(n_991), .Y(n_995) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_445), .Y(n_657) );
OAI33xp33_ASAP7_75t_L g978 ( .A1(n_445), .A2(n_959), .A3(n_979), .B1(n_983), .B2(n_986), .B3(n_989), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_448), .A2(n_574), .B1(n_579), .B2(n_591), .Y(n_590) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_451), .A2(n_588), .B1(n_779), .B2(n_780), .C(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g611 ( .A(n_458), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g684 ( .A(n_462), .Y(n_684) );
BUFx3_ASAP7_75t_L g742 ( .A(n_462), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_464), .A2(n_488), .B1(n_1000), .B2(n_1001), .Y(n_999) );
INVx1_ASAP7_75t_L g532 ( .A(n_475), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_475), .B(n_844), .Y(n_851) );
XOR2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_565), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_524), .B(n_526), .Y(n_478) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_485), .Y(n_804) );
BUFx3_ASAP7_75t_L g913 ( .A(n_485), .Y(n_913) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_502), .B(n_509), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
OAI221xp5_ASAP7_75t_L g558 ( .A1(n_499), .A2(n_510), .B1(n_559), .B2(n_561), .C(n_562), .Y(n_558) );
INVx5_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx6_ASAP7_75t_L g701 ( .A(n_501), .Y(n_701) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g704 ( .A(n_507), .Y(n_704) );
INVx2_ASAP7_75t_L g955 ( .A(n_507), .Y(n_955) );
OAI211xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_511), .B(n_512), .C(n_517), .Y(n_509) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g860 ( .A(n_514), .Y(n_860) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g659 ( .A(n_519), .Y(n_659) );
INVx2_ASAP7_75t_SL g673 ( .A(n_519), .Y(n_673) );
INVx2_ASAP7_75t_L g782 ( .A(n_519), .Y(n_782) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_520), .Y(n_609) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_522), .Y(n_660) );
BUFx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g675 ( .A(n_523), .Y(n_675) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_523), .Y(n_790) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_538), .B(n_539), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_528), .B(n_535), .Y(n_527) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g629 ( .A(n_531), .Y(n_629) );
INVx2_ASAP7_75t_L g757 ( .A(n_531), .Y(n_757) );
BUFx2_ASAP7_75t_L g767 ( .A(n_538), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_538), .A2(n_884), .B1(n_898), .B2(n_906), .C(n_907), .Y(n_883) );
OAI31xp33_ASAP7_75t_L g1256 ( .A1(n_538), .A2(n_1257), .A3(n_1261), .B(n_1265), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B1(n_553), .B2(n_558), .Y(n_539) );
OAI33xp33_ASAP7_75t_L g568 ( .A1(n_540), .A2(n_569), .A3(n_572), .B1(n_575), .B2(n_580), .B3(n_583), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_540), .A2(n_819), .B1(n_824), .B2(n_828), .Y(n_818) );
OAI33xp33_ASAP7_75t_L g1304 ( .A1(n_540), .A2(n_583), .A3(n_1305), .B1(n_1312), .B2(n_1316), .B3(n_1320), .Y(n_1304) );
OAI211xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_545), .C(n_550), .Y(n_541) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g641 ( .A(n_546), .Y(n_641) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx8_ASAP7_75t_L g564 ( .A(n_547), .Y(n_564) );
BUFx3_ASAP7_75t_L g868 ( .A(n_547), .Y(n_868) );
BUFx2_ASAP7_75t_L g650 ( .A(n_549), .Y(n_650) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx5_ASAP7_75t_L g648 ( .A(n_552), .Y(n_648) );
BUFx12f_ASAP7_75t_L g921 ( .A(n_552), .Y(n_921) );
INVx1_ASAP7_75t_L g654 ( .A(n_553), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g730 ( .A(n_554), .Y(n_730) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g830 ( .A(n_555), .Y(n_830) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g646 ( .A(n_560), .Y(n_646) );
INVx1_ASAP7_75t_L g652 ( .A(n_560), .Y(n_652) );
INVx3_ASAP7_75t_L g945 ( .A(n_560), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_561), .A2(n_703), .B1(n_716), .B2(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g823 ( .A(n_564), .Y(n_823) );
INVx8_ASAP7_75t_L g877 ( .A(n_564), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_592), .C(n_602), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_584), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_571), .A2(n_582), .B1(n_588), .B2(n_589), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_578), .A2(n_1313), .B1(n_1314), .B2(n_1315), .Y(n_1312) );
INVx1_ASAP7_75t_L g879 ( .A(n_583), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_589), .A2(n_707), .B1(n_785), .B2(n_786), .C(n_787), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_589), .A2(n_955), .B1(n_987), .B2(n_988), .Y(n_986) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_589), .Y(n_1252) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_601), .A2(n_794), .B1(n_797), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_610), .B2(n_611), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_608), .A2(n_794), .B1(n_795), .B2(n_797), .C(n_798), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_608), .A2(n_749), .B1(n_894), .B2(n_896), .Y(n_905) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_609), .Y(n_857) );
INVx3_ASAP7_75t_L g864 ( .A(n_609), .Y(n_864) );
INVx1_ASAP7_75t_L g771 ( .A(n_613), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_691), .B1(n_692), .B2(n_768), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g769 ( .A(n_617), .Y(n_769) );
NAND4xp25_ASAP7_75t_SL g618 ( .A(n_619), .B(n_634), .C(n_655), .D(n_676), .Y(n_618) );
AO21x1_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_625), .B(n_632), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_622), .A2(n_624), .B1(n_839), .B2(n_840), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_622), .A2(n_624), .B1(n_886), .B2(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g755 ( .A(n_624), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_624), .A2(n_754), .B1(n_807), .B2(n_808), .Y(n_813) );
INVx1_ASAP7_75t_L g1260 ( .A(n_624), .Y(n_1260) );
INVx2_ASAP7_75t_L g1294 ( .A(n_624), .Y(n_1294) );
INVx1_ASAP7_75t_L g815 ( .A(n_627), .Y(n_815) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_631), .Y(n_761) );
CKINVDCx14_ASAP7_75t_R g632 ( .A(n_633), .Y(n_632) );
AOI33xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .A3(n_644), .B1(n_649), .B2(n_651), .B3(n_654), .Y(n_634) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI33xp33_ASAP7_75t_L g865 ( .A1(n_636), .A2(n_866), .A3(n_870), .B1(n_873), .B2(n_876), .B3(n_879), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_636), .B(n_920), .C(n_922), .Y(n_919) );
BUFx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g811 ( .A(n_643), .Y(n_811) );
INVx1_ASAP7_75t_L g869 ( .A(n_643), .Y(n_869) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g653 ( .A(n_648), .Y(n_653) );
INVx2_ASAP7_75t_R g872 ( .A(n_648), .Y(n_872) );
AOI33xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .A3(n_661), .B1(n_668), .B2(n_669), .B3(n_672), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_657), .A2(n_778), .B1(n_784), .B2(n_791), .Y(n_777) );
OAI33xp33_ASAP7_75t_L g1244 ( .A1(n_657), .A2(n_1245), .A3(n_1250), .B1(n_1251), .B2(n_1253), .B3(n_1255), .Y(n_1244) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g902 ( .A(n_667), .Y(n_902) );
INVx2_ASAP7_75t_L g713 ( .A(n_669), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_669), .B(n_917), .C(n_918), .Y(n_916) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx3_ASAP7_75t_L g783 ( .A(n_675), .Y(n_783) );
AO21x1_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B(n_690), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_678), .B(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1270 ( .A(n_678), .Y(n_1270) );
AND2x4_ASAP7_75t_SL g1279 ( .A(n_678), .B(n_1280), .Y(n_1279) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .C(n_689), .Y(n_680) );
INVx5_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_687), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
BUFx2_ASAP7_75t_SL g711 ( .A(n_687), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_687), .A2(n_938), .B1(n_951), .B2(n_957), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_687), .A2(n_955), .B1(n_984), .B2(n_985), .Y(n_983) );
BUFx3_ASAP7_75t_L g1329 ( .A(n_687), .Y(n_1329) );
INVx2_ASAP7_75t_L g744 ( .A(n_688), .Y(n_744) );
INVx2_ASAP7_75t_L g1299 ( .A(n_688), .Y(n_1299) );
INVx1_ASAP7_75t_L g746 ( .A(n_689), .Y(n_746) );
INVx3_ASAP7_75t_L g1272 ( .A(n_689), .Y(n_1272) );
AOI21xp33_ASAP7_75t_L g792 ( .A1(n_690), .A2(n_793), .B(n_806), .Y(n_792) );
AO21x1_ASAP7_75t_L g837 ( .A1(n_690), .A2(n_838), .B(n_841), .Y(n_837) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_735), .C(n_751), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_718), .Y(n_694) );
OAI33xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .A3(n_702), .B1(n_706), .B2(n_713), .B3(n_714), .Y(n_695) );
OAI22xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_698), .A2(n_710), .B1(n_721), .B2(n_724), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_700), .A2(n_712), .B1(n_721), .B2(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_701), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
OAI22xp33_ASAP7_75t_SL g1251 ( .A1(n_704), .A2(n_1232), .B1(n_1243), .B2(n_1252), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx4_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI33xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .A3(n_726), .B1(n_728), .B2(n_730), .B3(n_731), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_729), .A2(n_779), .B1(n_820), .B2(n_821), .C(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g1311 ( .A(n_734), .Y(n_1311) );
OAI31xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .A3(n_747), .B(n_750), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_743), .A2(n_759), .B1(n_761), .B2(n_762), .Y(n_758) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_SL g1301 ( .A(n_749), .Y(n_1301) );
OAI31xp33_ASAP7_75t_SL g1268 ( .A1(n_750), .A2(n_1269), .A3(n_1271), .B(n_1275), .Y(n_1268) );
OAI31xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_756), .A3(n_763), .B(n_767), .Y(n_751) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
BUFx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_831), .B2(n_832), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NOR4xp25_ASAP7_75t_L g776 ( .A(n_777), .B(n_792), .C(n_809), .D(n_818), .Y(n_776) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g1254 ( .A(n_791), .Y(n_1254) );
INVx1_ASAP7_75t_L g1277 ( .A(n_795), .Y(n_1277) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .C(n_805), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AOI31xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_813), .A3(n_814), .B(n_816), .Y(n_809) );
AO21x1_ASAP7_75t_L g847 ( .A1(n_816), .A2(n_848), .B(n_852), .Y(n_847) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI31xp33_ASAP7_75t_L g1287 ( .A1(n_817), .A2(n_1288), .A3(n_1289), .B(n_1293), .Y(n_1287) );
INVx1_ASAP7_75t_L g871 ( .A(n_820), .Y(n_871) );
OAI33xp33_ASAP7_75t_L g1228 ( .A1(n_828), .A2(n_1229), .A3(n_1230), .B1(n_1234), .B2(n_1237), .B3(n_1240), .Y(n_1228) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
BUFx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
BUFx2_ASAP7_75t_L g925 ( .A(n_830), .Y(n_925) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_929), .B2(n_1010), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_882), .Y(n_834) );
INVx1_ASAP7_75t_L g880 ( .A(n_836), .Y(n_880) );
NAND4xp75_ASAP7_75t_L g836 ( .A(n_837), .B(n_847), .C(n_853), .D(n_865), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_846), .Y(n_841) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_854), .Y(n_915) );
INVx2_ASAP7_75t_SL g854 ( .A(n_855), .Y(n_854) );
OAI33xp33_ASAP7_75t_L g1323 ( .A1(n_855), .A2(n_959), .A3(n_1324), .B1(n_1328), .B2(n_1330), .B3(n_1331), .Y(n_1323) );
INVx2_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
BUFx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g928 ( .A(n_868), .Y(n_928) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_888), .C(n_893), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_896), .B2(n_897), .Y(n_893) );
INVx2_ASAP7_75t_L g1266 ( .A(n_895), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_901), .C(n_905), .Y(n_898) );
OAI31xp33_ASAP7_75t_L g1295 ( .A1(n_906), .A2(n_1296), .A3(n_1300), .B(n_1302), .Y(n_1295) );
NAND4xp25_ASAP7_75t_L g907 ( .A(n_908), .B(n_916), .C(n_919), .D(n_923), .Y(n_907) );
NAND3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_914), .C(n_915), .Y(n_908) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .C(n_926), .Y(n_923) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
BUFx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g1010 ( .A(n_930), .Y(n_1010) );
XNOR2x1_ASAP7_75t_L g930 ( .A(n_931), .B(n_975), .Y(n_930) );
XNOR2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .Y(n_931) );
AND3x1_ASAP7_75t_L g933 ( .A(n_934), .B(n_960), .C(n_968), .Y(n_933) );
NOR2xp33_ASAP7_75t_SL g934 ( .A(n_935), .B(n_952), .Y(n_934) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx2_ASAP7_75t_L g1314 ( .A(n_945), .Y(n_1314) );
OAI22xp33_ASAP7_75t_L g1230 ( .A1(n_948), .A2(n_1231), .B1(n_1232), .B2(n_1233), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_948), .A2(n_1241), .B1(n_1242), .B2(n_1243), .Y(n_1240) );
INVx2_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
INVx3_ASAP7_75t_L g1308 ( .A(n_949), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_957), .A2(n_1313), .B1(n_1318), .B2(n_1329), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_957), .A2(n_1309), .B1(n_1322), .B2(n_1329), .Y(n_1330) );
AND3x1_ASAP7_75t_L g976 ( .A(n_977), .B(n_997), .C(n_1004), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_992), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_981), .A2(n_1315), .B1(n_1319), .B2(n_1325), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1017), .Y(n_1011) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1012), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1015), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1013), .B(n_1016), .Y(n_1333) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1013), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1016), .B(n_1335), .Y(n_1337) );
OAI21xp33_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1219), .B(n_1223), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1174), .Y(n_1020) );
NAND3xp33_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1113), .C(n_1143), .Y(n_1021) );
AOI211xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1043), .B(n_1076), .C(n_1093), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1023), .B(n_1117), .Y(n_1116) );
AOI322xp5_ASAP7_75t_L g1125 ( .A1(n_1023), .A2(n_1051), .A3(n_1074), .B1(n_1078), .B2(n_1121), .C1(n_1126), .C2(n_1129), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1039), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1024), .B(n_1155), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1024), .B(n_1156), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1024), .B(n_1067), .Y(n_1211) );
INVx3_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1025), .B(n_1081), .Y(n_1080) );
INVx3_ASAP7_75t_L g1092 ( .A(n_1025), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1025), .B(n_1039), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1025), .B(n_1142), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1025), .B(n_1117), .Y(n_1160) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1025), .B(n_1122), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1025), .B(n_1101), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1025), .B(n_1039), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1025), .B(n_1215), .Y(n_1214) );
AND2x4_ASAP7_75t_SL g1025 ( .A(n_1026), .B(n_1033), .Y(n_1025) );
AND2x6_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1028), .B(n_1032), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_1028), .B(n_1035), .Y(n_1034) );
AND2x6_ASAP7_75t_L g1037 ( .A(n_1028), .B(n_1038), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1028), .B(n_1032), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1028), .B(n_1032), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1030), .B(n_1036), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1222 ( .A(n_1031), .Y(n_1222) );
OAI21xp5_ASAP7_75t_L g1334 ( .A1(n_1032), .A2(n_1335), .B(n_1336), .Y(n_1334) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_1039), .B(n_1073), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1039), .B(n_1064), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1156 ( .A(n_1039), .B(n_1064), .Y(n_1156) );
OAI221xp5_ASAP7_75t_SL g1180 ( .A1(n_1039), .A2(n_1044), .B1(n_1181), .B2(n_1182), .C(n_1183), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1042), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1079 ( .A(n_1040), .B(n_1042), .Y(n_1079) );
A2O1A1Ixp33_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1058), .B(n_1062), .C(n_1070), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1044), .B(n_1086), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1044), .B(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1045), .B(n_1074), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1051), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_1046), .B(n_1059), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1046), .B(n_1096), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1046), .B(n_1127), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1046), .B(n_1151), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1046), .B(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1046), .B(n_1088), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_1047), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1047), .B(n_1051), .Y(n_1075) );
NOR2xp33_ASAP7_75t_L g1098 ( .A(n_1047), .B(n_1067), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1047), .B(n_1055), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1047), .B(n_1088), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1047), .B(n_1067), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1047), .B(n_1151), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1050), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1048), .B(n_1050), .Y(n_1133) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1051), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1051), .B(n_1197), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1055), .Y(n_1051) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1052), .Y(n_1061) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1052), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1055), .B(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1055), .Y(n_1097) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1055), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_1055), .B(n_1061), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1199 ( .A(n_1058), .B(n_1200), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1059), .B(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1060), .B(n_1107), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1061), .B(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1061), .Y(n_1151) );
INVxp33_ASAP7_75t_SL g1149 ( .A(n_1062), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1067), .Y(n_1062) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1063), .Y(n_1108) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1063), .Y(n_1177) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1064), .Y(n_1073) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1064), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1066), .Y(n_1064) );
INVx3_ASAP7_75t_L g1074 ( .A(n_1067), .Y(n_1074) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1067), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_1067), .B(n_1073), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1067), .B(n_1158), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1069), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1075), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1147 ( .A(n_1072), .B(n_1148), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1074), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1073), .B(n_1079), .Y(n_1078) );
NAND3xp33_ASAP7_75t_L g1102 ( .A(n_1074), .B(n_1081), .C(n_1087), .Y(n_1102) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1074), .Y(n_1107) );
NOR2xp33_ASAP7_75t_L g1129 ( .A(n_1074), .B(n_1130), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1074), .B(n_1164), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1074), .B(n_1150), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1075), .B(n_1090), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1075), .B(n_1118), .Y(n_1124) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1075), .Y(n_1161) );
OAI21xp5_ASAP7_75t_L g1207 ( .A1(n_1075), .A2(n_1208), .B(n_1209), .Y(n_1207) );
OAI21xp33_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1087), .B(n_1089), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1080), .C(n_1085), .Y(n_1077) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1078), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_1079), .A2(n_1147), .B1(n_1149), .B2(n_1150), .Y(n_1146) );
OAI211xp5_ASAP7_75t_L g1165 ( .A1(n_1079), .A2(n_1166), .B(n_1168), .C(n_1172), .Y(n_1165) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1079), .Y(n_1215) );
OAI21xp33_ASAP7_75t_L g1175 ( .A1(n_1080), .A2(n_1176), .B(n_1180), .Y(n_1175) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1082), .Y(n_1091) );
OAI31xp33_ASAP7_75t_SL g1143 ( .A1(n_1082), .A2(n_1144), .A3(n_1153), .B(n_1165), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1085), .B(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NAND2xp5_ASAP7_75t_SL g1167 ( .A(n_1086), .B(n_1127), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1086), .B(n_1155), .Y(n_1206) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1090), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1092), .Y(n_1090) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1091), .Y(n_1110) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1092), .Y(n_1152) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1099), .B1(n_1100), .B2(n_1102), .C(n_1103), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1098), .Y(n_1095) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1096), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1096), .B(n_1133), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1098), .B(n_1127), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1098), .B(n_1112), .Y(n_1181) );
INVx2_ASAP7_75t_SL g1142 ( .A(n_1099), .Y(n_1142) );
OAI322xp33_ASAP7_75t_L g1131 ( .A1(n_1100), .A2(n_1132), .A3(n_1134), .B1(n_1135), .B2(n_1136), .C1(n_1138), .C2(n_1140), .Y(n_1131) );
CKINVDCx14_ASAP7_75t_R g1100 ( .A(n_1101), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1101), .B(n_1107), .Y(n_1170) );
NAND4xp25_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1106), .C(n_1109), .D(n_1111), .Y(n_1103) );
OAI21xp5_ASAP7_75t_L g1162 ( .A1(n_1104), .A2(n_1163), .B(n_1164), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1104), .B(n_1179), .Y(n_1201) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1107), .B(n_1123), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1107), .B(n_1142), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1107), .B(n_1217), .Y(n_1216) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_1109), .A2(n_1114), .B1(n_1116), .B2(n_1119), .C(n_1131), .Y(n_1113) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_1111), .A2(n_1121), .B1(n_1127), .B2(n_1142), .C(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI21xp33_ASAP7_75t_L g1120 ( .A1(n_1116), .A2(n_1121), .B(n_1123), .Y(n_1120) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1117), .Y(n_1182) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
NAND3xp33_ASAP7_75t_SL g1119 ( .A(n_1120), .B(n_1124), .C(n_1125), .Y(n_1119) );
CKINVDCx14_ASAP7_75t_R g1121 ( .A(n_1122), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1126), .B(n_1173), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1127), .B(n_1133), .Y(n_1139) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1130), .Y(n_1171) );
OAI21xp33_ASAP7_75t_L g1204 ( .A1(n_1130), .A2(n_1205), .B(n_1207), .Y(n_1204) );
OAI321xp33_ASAP7_75t_L g1153 ( .A1(n_1133), .A2(n_1154), .A3(n_1157), .B1(n_1159), .B2(n_1161), .C(n_1162), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_1133), .B(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
AOI21xp33_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1146), .B(n_1152), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1148), .B(n_1158), .Y(n_1157) );
AOI211xp5_ASAP7_75t_L g1202 ( .A1(n_1155), .A2(n_1203), .B(n_1204), .C(n_1212), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1155), .B(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_1159), .A2(n_1213), .B1(n_1216), .B2(n_1218), .Y(n_1212) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1164), .Y(n_1187) );
OAI21xp5_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1170), .B(n_1171), .Y(n_1168) );
NAND4xp25_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1185), .C(n_1198), .D(n_1202), .Y(n_1174) );
NOR2xp33_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1182), .B(n_1196), .Y(n_1195) );
AOI211xp5_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1188), .B(n_1189), .C(n_1194), .Y(n_1185) );
AOI21xp33_ASAP7_75t_SL g1189 ( .A1(n_1190), .A2(n_1192), .B(n_1193), .Y(n_1189) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1190), .Y(n_1203) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1193), .B(n_1195), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1201), .Y(n_1198) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
CKINVDCx20_ASAP7_75t_R g1219 ( .A(n_1220), .Y(n_1219) );
CKINVDCx20_ASAP7_75t_R g1220 ( .A(n_1221), .Y(n_1220) );
INVx4_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
NAND3xp33_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1256), .C(n_1268), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1244), .Y(n_1227) );
OAI22xp33_ASAP7_75t_L g1245 ( .A1(n_1231), .A2(n_1241), .B1(n_1246), .B2(n_1248), .Y(n_1245) );
OAI22xp33_ASAP7_75t_L g1255 ( .A1(n_1236), .A2(n_1239), .B1(n_1246), .B2(n_1248), .Y(n_1255) );
INVx2_ASAP7_75t_SL g1246 ( .A(n_1247), .Y(n_1246) );
BUFx3_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
NAND3xp33_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1295), .C(n_1303), .Y(n_1286) );
NOR2xp33_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1323), .Y(n_1303) );
OAI22xp33_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B1(n_1309), .B2(n_1310), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1306), .A2(n_1321), .B1(n_1325), .B2(n_1327), .Y(n_1324) );
BUFx4f_ASAP7_75t_SL g1307 ( .A(n_1308), .Y(n_1307) );
INVxp67_ASAP7_75t_SL g1310 ( .A(n_1311), .Y(n_1310) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
HB1xp67_ASAP7_75t_SL g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
endmodule