module fake_jpeg_9534_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_35),
.B1(n_17),
.B2(n_39),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_17),
.B(n_28),
.C(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_30),
.Y(n_55)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_16),
.B1(n_28),
.B2(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_15),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_18),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_51),
.B(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_71),
.Y(n_102)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_74),
.B1(n_34),
.B2(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_27),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_85),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_88),
.B(n_63),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_31),
.B(n_44),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_56),
.C(n_31),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_58),
.C(n_56),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_97),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_34),
.B1(n_49),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_98),
.B1(n_99),
.B2(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_73),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_34),
.B1(n_49),
.B2(n_32),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_53),
.B1(n_60),
.B2(n_44),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_32),
.B1(n_40),
.B2(n_53),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_40),
.B1(n_19),
.B2(n_31),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_65),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_100),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_48),
.B1(n_26),
.B2(n_23),
.C(n_25),
.Y(n_141)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_74),
.B1(n_76),
.B2(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_61),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_72),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_58),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_123),
.B(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_82),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_96),
.C(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_68),
.B1(n_71),
.B2(n_56),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_33),
.B(n_37),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_97),
.C(n_101),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_141),
.C(n_103),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_93),
.C(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_130),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_107),
.B(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_140),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_101),
.B1(n_23),
.B2(n_25),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_118),
.B(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_137),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_158),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_113),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_156),
.B(n_80),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_138),
.B1(n_131),
.B2(n_139),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_127),
.B1(n_134),
.B2(n_118),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_120),
.B1(n_119),
.B2(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_164),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_158),
.A2(n_138),
.B1(n_86),
.B2(n_126),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_150),
.B1(n_86),
.B2(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_130),
.C(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_170),
.C(n_171),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_1),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_37),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_80),
.C(n_33),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_33),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_174),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_146),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_154),
.B(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_178),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_179),
.B1(n_167),
.B2(n_2),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_144),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_170),
.C(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_168),
.C(n_163),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_37),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.C(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_183),
.B(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_14),
.C(n_13),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_13),
.C(n_11),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_11),
.C(n_2),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_1),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

OAI321xp33_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_194),
.A3(n_3),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_188),
.B(n_5),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.C(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_192),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

AOI21x1_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_201),
.B(n_202),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_192),
.B(n_8),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);


endmodule