module fake_netlist_6_3956_n_1774 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1774);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1774;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_66),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_71),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_58),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_46),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_27),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_28),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_60),
.Y(n_170)
);

INVxp33_ASAP7_75t_SL g171 ( 
.A(n_76),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_75),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_14),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_62),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_38),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_23),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_52),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_34),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_102),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_32),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_17),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_28),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_100),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_103),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_26),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_132),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_59),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_31),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_51),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_54),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_46),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_114),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_10),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_34),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_32),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_33),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_63),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_31),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_19),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_94),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_18),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_84),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_98),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_6),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_5),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_107),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_7),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_51),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_9),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_130),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_68),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_140),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_136),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_48),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_138),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_52),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_24),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_21),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_2),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_99),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_57),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_88),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_125),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_87),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_27),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_92),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_93),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_85),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_50),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_22),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_11),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_144),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_20),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_142),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_137),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_105),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_55),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_97),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_53),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_141),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_91),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_108),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_21),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_65),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_8),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_129),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_154),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_22),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_29),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_20),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_80),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_14),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_19),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_29),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_50),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_155),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_124),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_64),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_23),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_49),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_24),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_95),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_157),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_158),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_173),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_173),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_173),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_0),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_173),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_164),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_215),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_215),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_170),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_215),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_228),
.B(n_1),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_168),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_215),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_215),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_185),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_180),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_277),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_292),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_228),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_160),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_160),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_191),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_191),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_252),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_195),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_195),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_172),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_205),
.B(n_3),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_221),
.B(n_3),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_5),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_205),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_209),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_209),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_304),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_175),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_180),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_235),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_237),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_161),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_237),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_177),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_167),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_211),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_181),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_184),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_239),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_167),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_189),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_235),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_194),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_217),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_196),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_197),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_182),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_217),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_234),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_167),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_171),
.B(n_7),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_199),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_231),
.B(n_10),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_200),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_286),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

BUFx8_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_182),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_L g393 ( 
.A(n_325),
.B(n_230),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_188),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g397 ( 
.A(n_315),
.B(n_188),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_315),
.B(n_231),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_366),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_186),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_316),
.B(n_192),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_348),
.B(n_299),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_335),
.A2(n_248),
.B1(n_290),
.B2(n_261),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_360),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_316),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_159),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_317),
.B(n_192),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_326),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_319),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_321),
.B(n_246),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_321),
.B(n_246),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g420 ( 
.A1(n_322),
.A2(n_243),
.B(n_234),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_324),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_201),
.Y(n_424)
);

AND2x2_ASAP7_75t_SL g425 ( 
.A(n_378),
.B(n_262),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_336),
.B(n_186),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_336),
.B(n_216),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_327),
.B(n_216),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_328),
.B(n_203),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_329),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_329),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_331),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_339),
.B(n_208),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_331),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_338),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_318),
.B(n_159),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_339),
.B(n_262),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_341),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_342),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_387),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_340),
.B1(n_343),
.B2(n_347),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_359),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_447),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_425),
.A2(n_441),
.B1(n_386),
.B2(n_393),
.Y(n_455)
);

AOI21x1_ASAP7_75t_L g456 ( 
.A1(n_401),
.A2(n_165),
.B(n_162),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_394),
.B(n_344),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_447),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_403),
.A2(n_340),
.B1(n_298),
.B2(n_302),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_425),
.B(n_311),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_386),
.B(n_254),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_347),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_386),
.A2(n_330),
.B1(n_333),
.B2(n_353),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_387),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_162),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

OR2x6_ASAP7_75t_L g475 ( 
.A(n_400),
.B(n_165),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_386),
.B(n_213),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_384),
.B(n_167),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_394),
.B(n_345),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_403),
.A2(n_179),
.B1(n_309),
.B2(n_308),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_404),
.B(n_334),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_411),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_390),
.B(n_166),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_425),
.B(n_312),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_441),
.A2(n_241),
.B1(n_163),
.B2(n_169),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_390),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_399),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_425),
.A2(n_220),
.B1(n_243),
.B2(n_245),
.Y(n_494)
);

BUFx6f_ASAP7_75t_SL g495 ( 
.A(n_390),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_313),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_404),
.A2(n_382),
.B1(n_245),
.B2(n_256),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_411),
.B(n_320),
.Y(n_499)
);

INVx4_ASAP7_75t_SL g500 ( 
.A(n_388),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_384),
.B(n_167),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_384),
.B(n_167),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_384),
.B(n_167),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_424),
.B(n_323),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_412),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_412),
.B(n_346),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_390),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_420),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_388),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_414),
.B(n_354),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_431),
.B(n_361),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_390),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_420),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_444),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_399),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_384),
.B(n_167),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_414),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_396),
.A2(n_233),
.B1(n_174),
.B2(n_176),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_388),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_426),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_390),
.B(n_166),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_435),
.B(n_364),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_395),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_386),
.B(n_365),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_396),
.A2(n_236),
.B1(n_178),
.B2(n_183),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_395),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_395),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_395),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_388),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_444),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_386),
.B(n_372),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_426),
.B(n_373),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_388),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_443),
.B(n_167),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_443),
.B(n_263),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_428),
.B(n_398),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_385),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_426),
.B(n_345),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_435),
.B(n_379),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_385),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_431),
.A2(n_198),
.B1(n_259),
.B2(n_257),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_393),
.A2(n_220),
.B1(n_256),
.B2(n_258),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_388),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_388),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_385),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_406),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_427),
.B(n_381),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_443),
.B(n_263),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_413),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_413),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_443),
.B(n_285),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_406),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_413),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_427),
.A2(n_258),
.B1(n_268),
.B2(n_307),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_413),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_413),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_406),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_427),
.A2(n_268),
.B1(n_301),
.B2(n_307),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_415),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_443),
.B(n_285),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_405),
.B(n_213),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_398),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_413),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_413),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_398),
.B(n_291),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_398),
.B(n_291),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_405),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_415),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_417),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_417),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_434),
.B(n_350),
.Y(n_593)
);

AND2x2_ASAP7_75t_SL g594 ( 
.A(n_398),
.B(n_230),
.Y(n_594)
);

INVxp33_ASAP7_75t_SL g595 ( 
.A(n_416),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_452),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_455),
.B(n_210),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_461),
.A2(n_368),
.B1(n_370),
.B2(n_275),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_497),
.B(n_401),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_533),
.B(n_230),
.Y(n_602)
);

OAI221xp5_ASAP7_75t_L g603 ( 
.A1(n_494),
.A2(n_301),
.B1(n_190),
.B2(n_281),
.C(n_193),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_508),
.B(n_401),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_547),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

BUFx6f_ASAP7_75t_SL g607 ( 
.A(n_547),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_537),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_536),
.B(n_401),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_537),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_555),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

NOR3xp33_ASAP7_75t_L g613 ( 
.A(n_459),
.B(n_479),
.C(n_499),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_488),
.A2(n_250),
.B1(n_218),
.B2(n_278),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_533),
.A2(n_284),
.B1(n_238),
.B2(n_255),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_558),
.B(n_401),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_481),
.A2(n_271),
.B1(n_219),
.B2(n_287),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_554),
.B(n_230),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_509),
.B(n_187),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_509),
.B(n_202),
.Y(n_621)
);

INVx8_ASAP7_75t_L g622 ( 
.A(n_473),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_448),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_542),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_554),
.B(n_401),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_542),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_554),
.B(n_230),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_554),
.B(n_555),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_448),
.B(n_416),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_464),
.A2(n_249),
.B1(n_193),
.B2(n_212),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_520),
.B(n_457),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_464),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_594),
.B(n_409),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_550),
.B(n_204),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_557),
.A2(n_190),
.B(n_212),
.C(n_310),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_457),
.B(n_409),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_513),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_513),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_594),
.B(n_513),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_543),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_521),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_568),
.B(n_519),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_521),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_594),
.B(n_409),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_521),
.B(n_409),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_478),
.B(n_409),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_478),
.B(n_409),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_454),
.A2(n_419),
.B(n_418),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_547),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_543),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_495),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_481),
.B(n_206),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_559),
.B(n_418),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_559),
.B(n_418),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_557),
.B(n_418),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_527),
.B(n_383),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_559),
.B(n_418),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_544),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_454),
.B(n_418),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_458),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_473),
.A2(n_475),
.B1(n_464),
.B2(n_538),
.Y(n_663)
);

AND2x6_ASAP7_75t_SL g664 ( 
.A(n_464),
.B(n_350),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_584),
.B(n_442),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_544),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_458),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_474),
.B(n_442),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_584),
.B(n_442),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_207),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_544),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_584),
.B(n_442),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_473),
.A2(n_240),
.B1(n_297),
.B2(n_267),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_474),
.B(n_442),
.Y(n_674)
);

INVx8_ASAP7_75t_L g675 ( 
.A(n_473),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_464),
.B(n_214),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_549),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_486),
.B(n_524),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_549),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_473),
.B(n_224),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_547),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_487),
.B(n_442),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_486),
.B(n_445),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_530),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_445),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_549),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_487),
.B(n_280),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_493),
.B(n_434),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_583),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_450),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_475),
.B(n_225),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_595),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_489),
.B(n_289),
.C(n_229),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_593),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_551),
.A2(n_419),
.B(n_397),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_541),
.B(n_445),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_593),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_489),
.B(n_434),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_502),
.A2(n_281),
.B1(n_223),
.B2(n_226),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_475),
.A2(n_283),
.B1(n_306),
.B2(n_397),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_541),
.B(n_445),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_502),
.B(n_222),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_498),
.B(n_383),
.C(n_227),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_546),
.B(n_446),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_482),
.B(n_351),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_475),
.A2(n_247),
.B1(n_222),
.B2(n_310),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_475),
.B(n_251),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_515),
.A2(n_244),
.B1(n_303),
.B2(n_270),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_546),
.B(n_446),
.Y(n_709)
);

NAND2x1_ASAP7_75t_L g710 ( 
.A(n_467),
.B(n_415),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_482),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_515),
.B(n_223),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_527),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_516),
.A2(n_244),
.B1(n_303),
.B2(n_270),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_516),
.B(n_446),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_522),
.B(n_433),
.Y(n_716)
);

BUFx12f_ASAP7_75t_SL g717 ( 
.A(n_482),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_482),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_556),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_450),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_450),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_522),
.B(n_433),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_460),
.Y(n_723)
);

INVx4_ASAP7_75t_SL g724 ( 
.A(n_495),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_535),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_523),
.B(n_446),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_523),
.B(n_433),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_498),
.A2(n_226),
.B1(n_242),
.B2(n_247),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_535),
.B(n_421),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_535),
.B(n_421),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_476),
.B(n_433),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_527),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_527),
.B(n_561),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_535),
.B(n_556),
.Y(n_734)
);

BUFx5_ASAP7_75t_L g735 ( 
.A(n_560),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_548),
.A2(n_242),
.B1(n_249),
.B2(n_253),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_528),
.B(n_272),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_525),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_576),
.B(n_351),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_532),
.B(n_589),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_460),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_476),
.B(n_433),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_580),
.B(n_352),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_540),
.B(n_273),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_530),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_566),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_566),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_567),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_567),
.B(n_421),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_574),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_460),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_574),
.B(n_422),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_579),
.B(n_422),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_462),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_579),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_463),
.B(n_433),
.Y(n_756)
);

NOR2xp67_ASAP7_75t_L g757 ( 
.A(n_587),
.B(n_588),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_581),
.B(n_422),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_451),
.A2(n_266),
.B(n_253),
.C(n_260),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_589),
.B(n_383),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_463),
.B(n_433),
.Y(n_761)
);

NAND2x1p5_ASAP7_75t_L g762 ( 
.A(n_449),
.B(n_260),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_552),
.A2(n_266),
.B(n_264),
.C(n_357),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_759),
.A2(n_587),
.B(n_588),
.C(n_573),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_632),
.B(n_581),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_623),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_606),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_601),
.A2(n_468),
.B(n_467),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_597),
.B(n_465),
.C(n_264),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_643),
.B(n_583),
.Y(n_770)
);

AOI33xp33_ASAP7_75t_L g771 ( 
.A1(n_728),
.A2(n_371),
.A3(n_376),
.B1(n_375),
.B2(n_352),
.B3(n_357),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_735),
.B(n_551),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_740),
.B(n_480),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_600),
.B(n_363),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_609),
.B(n_590),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_613),
.A2(n_495),
.B1(n_590),
.B2(n_480),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_760),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_652),
.B(n_449),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_682),
.A2(n_562),
.B(n_564),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_692),
.B(n_495),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_643),
.A2(n_490),
.B1(n_483),
.B2(n_471),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_617),
.B(n_449),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_604),
.A2(n_468),
.B(n_467),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_735),
.B(n_551),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_596),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_694),
.B(n_449),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_630),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_757),
.A2(n_468),
.B(n_467),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_600),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_653),
.B(n_563),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_697),
.B(n_453),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_689),
.B(n_453),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_611),
.B(n_615),
.Y(n_793)
);

BUFx12f_ASAP7_75t_L g794 ( 
.A(n_664),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_738),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_633),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_628),
.A2(n_468),
.B(n_530),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_699),
.B(n_453),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_719),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_733),
.B(n_453),
.Y(n_800)
);

O2A1O1Ixp5_ASAP7_75t_L g801 ( 
.A1(n_731),
.A2(n_456),
.B(n_569),
.C(n_553),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_699),
.B(n_471),
.Y(n_802)
);

AOI21xp33_ASAP7_75t_L g803 ( 
.A1(n_635),
.A2(n_274),
.B(n_305),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_759),
.A2(n_569),
.B(n_573),
.C(n_553),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_708),
.B(n_471),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_708),
.B(n_471),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_738),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_733),
.A2(n_517),
.B1(n_565),
.B2(n_490),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_735),
.B(n_562),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_714),
.B(n_483),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_653),
.B(n_483),
.Y(n_811)
);

BUFx2_ASAP7_75t_SL g812 ( 
.A(n_607),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_682),
.A2(n_530),
.B(n_562),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_714),
.B(n_530),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_607),
.B(n_213),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_663),
.A2(n_517),
.B1(n_545),
.B2(n_490),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_637),
.B(n_483),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_620),
.B(n_490),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_646),
.A2(n_530),
.B(n_564),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_596),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_716),
.A2(n_564),
.B(n_582),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_746),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_646),
.A2(n_517),
.B(n_545),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_747),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_SL g825 ( 
.A1(n_640),
.A2(n_552),
.B(n_582),
.C(n_507),
.Y(n_825)
);

O2A1O1Ixp5_ASAP7_75t_L g826 ( 
.A1(n_731),
.A2(n_456),
.B(n_517),
.C(n_545),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_716),
.A2(n_565),
.B(n_545),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_603),
.A2(n_505),
.B(n_477),
.C(n_506),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_620),
.B(n_565),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_748),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_715),
.A2(n_565),
.B(n_491),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_621),
.B(n_232),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_750),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_647),
.B(n_462),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_726),
.A2(n_491),
.B(n_506),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_737),
.B(n_276),
.C(n_282),
.Y(n_836)
);

BUFx4f_ASAP7_75t_L g837 ( 
.A(n_657),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_665),
.A2(n_491),
.B(n_526),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_665),
.A2(n_491),
.B(n_526),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_648),
.B(n_462),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_687),
.A2(n_598),
.B(n_756),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_656),
.B(n_466),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_669),
.A2(n_491),
.B(n_505),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_669),
.A2(n_491),
.B(n_507),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_722),
.A2(n_503),
.B(n_466),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_755),
.B(n_466),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_705),
.B(n_469),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_596),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_662),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_737),
.B(n_744),
.C(n_676),
.Y(n_850)
);

OAI321xp33_ASAP7_75t_L g851 ( 
.A1(n_728),
.A2(n_376),
.A3(n_375),
.B1(n_371),
.B2(n_363),
.C(n_477),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_672),
.A2(n_491),
.B(n_577),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_735),
.B(n_500),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_605),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_672),
.A2(n_577),
.B(n_571),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_705),
.B(n_735),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_667),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_599),
.B(n_438),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_625),
.A2(n_577),
.B(n_571),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_735),
.B(n_469),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_629),
.A2(n_592),
.B1(n_591),
.B2(n_570),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_734),
.A2(n_571),
.B(n_572),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_640),
.A2(n_718),
.B1(n_711),
.B2(n_612),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_638),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_596),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_SL g866 ( 
.A1(n_634),
.A2(n_572),
.B(n_585),
.C(n_586),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_621),
.B(n_469),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_739),
.A2(n_232),
.B1(n_279),
.B2(n_288),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_654),
.A2(n_572),
.B(n_585),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_612),
.B(n_470),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_711),
.B(n_500),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_654),
.A2(n_586),
.B(n_585),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_655),
.A2(n_658),
.B(n_645),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_698),
.B(n_470),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_633),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_718),
.B(n_470),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_655),
.A2(n_586),
.B(n_591),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_688),
.B(n_279),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_722),
.A2(n_484),
.B(n_472),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_639),
.A2(n_592),
.B1(n_591),
.B2(n_578),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_658),
.A2(n_592),
.B(n_591),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_634),
.A2(n_592),
.B(n_578),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_642),
.B(n_500),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_608),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_739),
.A2(n_743),
.B1(n_744),
.B2(n_702),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_717),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_644),
.B(n_472),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_729),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_645),
.A2(n_578),
.B(n_575),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_SL g890 ( 
.A(n_670),
.B(n_294),
.C(n_300),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_712),
.B(n_472),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_727),
.A2(n_578),
.B(n_575),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_650),
.B(n_279),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_678),
.B(n_635),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_684),
.B(n_500),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_743),
.B(n_484),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_670),
.B(n_295),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_680),
.A2(n_575),
.B(n_570),
.C(n_534),
.Y(n_898)
);

NAND2x1_ASAP7_75t_L g899 ( 
.A(n_684),
.B(n_570),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_636),
.A2(n_496),
.B(n_484),
.C(n_534),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_693),
.B(n_296),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_680),
.A2(n_575),
.B1(n_570),
.B2(n_534),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_691),
.B(n_707),
.Y(n_903)
);

BUFx8_ASAP7_75t_L g904 ( 
.A(n_681),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_730),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_691),
.B(n_531),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_727),
.A2(n_531),
.B(n_529),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_707),
.B(n_531),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_610),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_602),
.B(n_529),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_602),
.B(n_529),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_636),
.A2(n_518),
.B(n_514),
.C(n_511),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_763),
.A2(n_518),
.B(n_514),
.C(n_511),
.Y(n_913)
);

NOR2x1_ASAP7_75t_L g914 ( 
.A(n_652),
.B(n_430),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_710),
.A2(n_518),
.B(n_514),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_668),
.B(n_674),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_676),
.A2(n_511),
.B1(n_510),
.B2(n_504),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_724),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_661),
.A2(n_510),
.B(n_504),
.Y(n_919)
);

BUFx2_ASAP7_75t_SL g920 ( 
.A(n_713),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_732),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_687),
.A2(n_504),
.B(n_503),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_614),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_684),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_684),
.A2(n_510),
.B(n_503),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_736),
.A2(n_501),
.B1(n_485),
.B2(n_496),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_725),
.B(n_500),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_619),
.A2(n_501),
.B(n_496),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_631),
.B(n_627),
.C(n_619),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_749),
.B(n_501),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_627),
.A2(n_485),
.B(n_423),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_703),
.B(n_232),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_756),
.B(n_761),
.C(n_618),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_622),
.B(n_440),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_700),
.A2(n_485),
.B1(n_430),
.B2(n_423),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_724),
.B(n_440),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_683),
.A2(n_423),
.B(n_430),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_761),
.A2(n_440),
.B(n_439),
.C(n_438),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_742),
.A2(n_437),
.B(n_436),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_706),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_752),
.B(n_437),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_673),
.A2(n_439),
.B(n_438),
.C(n_437),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_742),
.A2(n_437),
.B(n_436),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_753),
.B(n_436),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_622),
.B(n_74),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_758),
.B(n_436),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_690),
.B(n_432),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_745),
.A2(n_432),
.B(n_429),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_814),
.A2(n_916),
.B(n_782),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_799),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_785),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_888),
.B(n_685),
.Y(n_952)
);

AND2x2_ASAP7_75t_SL g953 ( 
.A(n_850),
.B(n_622),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_780),
.B(n_724),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_849),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_785),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_905),
.B(n_696),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_897),
.A2(n_675),
.B(n_649),
.C(n_616),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_793),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_894),
.B(n_701),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_885),
.A2(n_675),
.B1(n_762),
.B2(n_704),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_918),
.B(n_745),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_770),
.B(n_675),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_897),
.B(n_709),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_765),
.B(n_790),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_770),
.B(n_725),
.Y(n_966)
);

OAI21xp33_ASAP7_75t_SL g967 ( 
.A1(n_885),
.A2(n_677),
.B(n_624),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_822),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_903),
.B(n_666),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_800),
.B(n_671),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_SL g971 ( 
.A1(n_923),
.A2(n_762),
.B1(n_439),
.B2(n_679),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_795),
.Y(n_972)
);

BUFx8_ASAP7_75t_SL g973 ( 
.A(n_766),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_787),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_800),
.B(n_754),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_850),
.B(n_837),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_775),
.A2(n_695),
.B(n_626),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_836),
.A2(n_659),
.B1(n_641),
.B2(n_651),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_824),
.B(n_686),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_777),
.B(n_660),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_830),
.B(n_751),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_841),
.A2(n_741),
.B(n_723),
.C(n_721),
.Y(n_982)
);

BUFx4_ASAP7_75t_SL g983 ( 
.A(n_886),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_773),
.B(n_720),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_873),
.A2(n_432),
.B(n_433),
.C(n_429),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_836),
.B(n_432),
.C(n_429),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_774),
.B(n_67),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_768),
.A2(n_429),
.B(n_417),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_796),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_832),
.B(n_11),
.Y(n_990)
);

OR2x4_ASAP7_75t_L g991 ( 
.A(n_890),
.B(n_429),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_868),
.A2(n_429),
.B(n_417),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_L g993 ( 
.A(n_803),
.B(n_13),
.C(n_18),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_796),
.B(n_13),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_837),
.B(n_417),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_875),
.B(n_30),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_807),
.B(n_30),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_774),
.B(n_78),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_SL g999 ( 
.A1(n_898),
.A2(n_72),
.B(n_151),
.C(n_148),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_776),
.A2(n_429),
.B1(n_417),
.B2(n_36),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_904),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_915),
.A2(n_70),
.B(n_145),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_904),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_875),
.B(n_33),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_901),
.A2(n_429),
.B1(n_417),
.B2(n_61),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_932),
.B(n_35),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_940),
.B(n_35),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_833),
.B(n_417),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_789),
.B(n_921),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_783),
.A2(n_788),
.B(n_856),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_780),
.B(n_56),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_797),
.A2(n_79),
.B(n_122),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_811),
.B(n_123),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_811),
.B(n_818),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_918),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_901),
.B(n_121),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_818),
.B(n_119),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_884),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_789),
.B(n_111),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_896),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_868),
.B(n_36),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_769),
.A2(n_851),
.B1(n_893),
.B2(n_929),
.C(n_815),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_769),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_945),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_785),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_857),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_834),
.A2(n_110),
.B(n_109),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_785),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_848),
.B(n_101),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_812),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_820),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_SL g1032 ( 
.A(n_878),
.B(n_39),
.C(n_40),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_933),
.A2(n_829),
.B(n_764),
.C(n_858),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_933),
.A2(n_908),
.B(n_906),
.C(n_864),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_829),
.B(n_41),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_794),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_942),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_945),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_767),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_854),
.B(n_42),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_862),
.A2(n_81),
.B(n_89),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_828),
.A2(n_44),
.B(n_45),
.C(n_47),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_786),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_791),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_792),
.B(n_45),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_792),
.B(n_867),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_847),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_883),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1048)
);

OAI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_934),
.A2(n_863),
.B1(n_874),
.B2(n_848),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_920),
.B(n_865),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_772),
.A2(n_784),
.B(n_809),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_820),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_865),
.B(n_820),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_909),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_840),
.B(n_842),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_924),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_817),
.A2(n_860),
.B(n_825),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_930),
.B(n_941),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_887),
.B(n_846),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_820),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_871),
.B(n_772),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_936),
.B(n_914),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_871),
.B(n_784),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_936),
.A2(n_808),
.B1(n_816),
.B2(n_902),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_924),
.B(n_876),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_944),
.B(n_946),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_798),
.B(n_802),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_938),
.A2(n_866),
.B(n_804),
.C(n_880),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_801),
.A2(n_826),
.B(n_821),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_859),
.A2(n_872),
.B(n_855),
.C(n_869),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_924),
.B(n_781),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_924),
.B(n_910),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_771),
.B(n_917),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_870),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_805),
.A2(n_810),
.B(n_806),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_809),
.A2(n_844),
.B(n_843),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_838),
.A2(n_839),
.B(n_835),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_882),
.B(n_889),
.Y(n_1078)
);

AOI22x1_ASAP7_75t_L g1079 ( 
.A1(n_881),
.A2(n_877),
.B1(n_823),
.B2(n_819),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_911),
.B(n_827),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_779),
.B(n_947),
.Y(n_1081)
);

BUFx4f_ASAP7_75t_L g1082 ( 
.A(n_778),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_891),
.A2(n_853),
.B(n_813),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_919),
.B(n_937),
.Y(n_1084)
);

OR2x6_ASAP7_75t_SL g1085 ( 
.A(n_926),
.B(n_778),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_861),
.B(n_935),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_852),
.B(n_927),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_883),
.A2(n_912),
.B(n_900),
.C(n_913),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_845),
.Y(n_1089)
);

AND2x2_ASAP7_75t_SL g1090 ( 
.A(n_927),
.B(n_853),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_879),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_988),
.A2(n_922),
.B(n_943),
.Y(n_1092)
);

AO21x2_ASAP7_75t_L g1093 ( 
.A1(n_1069),
.A2(n_1033),
.B(n_1077),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1010),
.A2(n_939),
.B(n_907),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1015),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_SL g1096 ( 
.A(n_1022),
.B(n_931),
.C(n_892),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_949),
.A2(n_831),
.B(n_928),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_985),
.A2(n_1070),
.A3(n_1057),
.B(n_1014),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_963),
.A2(n_895),
.B1(n_899),
.B2(n_925),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_990),
.B(n_948),
.C(n_895),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_984),
.B(n_980),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1014),
.A2(n_964),
.B(n_1055),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1009),
.B(n_1062),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1076),
.A2(n_1083),
.B(n_1079),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_982),
.A2(n_977),
.B(n_1051),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_989),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_958),
.A2(n_965),
.B(n_966),
.C(n_1013),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_1015),
.B(n_986),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_974),
.B(n_959),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1007),
.B(n_1006),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1075),
.A2(n_976),
.B(n_1017),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1055),
.A2(n_1058),
.B(n_1066),
.Y(n_1112)
);

BUFx2_ASAP7_75t_R g1113 ( 
.A(n_973),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_993),
.A2(n_1021),
.B1(n_1000),
.B2(n_1032),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1069),
.A2(n_1017),
.B(n_1013),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_960),
.B(n_1020),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1034),
.A2(n_967),
.B(n_1035),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1086),
.A2(n_1046),
.B(n_1064),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1058),
.A2(n_1066),
.B(n_1078),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1042),
.A2(n_1016),
.B(n_1019),
.C(n_1045),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_960),
.A2(n_957),
.B1(n_952),
.B2(n_961),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1078),
.A2(n_1084),
.B(n_969),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_1024),
.B(n_1038),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_972),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_950),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_952),
.A2(n_957),
.B1(n_961),
.B2(n_955),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1000),
.A2(n_994),
.B1(n_996),
.B2(n_1004),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1030),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_983),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_SL g1130 ( 
.A1(n_1037),
.A2(n_1088),
.B(n_1023),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1080),
.A2(n_1067),
.B(n_1063),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1002),
.A2(n_1087),
.B(n_1041),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1068),
.A2(n_1081),
.B(n_1071),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1029),
.A2(n_992),
.B(n_970),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_975),
.A2(n_1049),
.B(n_1080),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1047),
.B(n_1074),
.Y(n_1137)
);

BUFx10_ASAP7_75t_L g1138 ( 
.A(n_1009),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1015),
.Y(n_1139)
);

AOI221x1_ASAP7_75t_L g1140 ( 
.A1(n_1012),
.A2(n_975),
.B1(n_971),
.B2(n_1027),
.C(n_1061),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1060),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_987),
.B(n_998),
.Y(n_1142)
);

AOI221x1_ASAP7_75t_L g1143 ( 
.A1(n_1089),
.A2(n_1091),
.B1(n_1073),
.B2(n_1044),
.C(n_1043),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_987),
.B(n_998),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1059),
.A2(n_1082),
.B1(n_968),
.B2(n_1026),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1039),
.Y(n_1146)
);

INVx3_ASAP7_75t_SL g1147 ( 
.A(n_1040),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1056),
.A2(n_995),
.B(n_953),
.Y(n_1148)
);

CKINVDCx11_ASAP7_75t_R g1149 ( 
.A(n_1036),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1008),
.A2(n_1053),
.A3(n_981),
.B(n_979),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_978),
.A2(n_962),
.B(n_956),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1005),
.A2(n_1050),
.B(n_1048),
.C(n_1054),
.Y(n_1152)
);

CKINVDCx11_ASAP7_75t_R g1153 ( 
.A(n_1085),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_1025),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1018),
.A2(n_1062),
.B(n_1090),
.C(n_1029),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1056),
.A2(n_999),
.B(n_951),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1067),
.B(n_1065),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1056),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_954),
.A2(n_991),
.B(n_1011),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1025),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1067),
.A2(n_962),
.B(n_1028),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_997),
.B(n_1028),
.C(n_1031),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_991),
.A2(n_1031),
.B(n_1025),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1052),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1067),
.A2(n_988),
.B(n_1010),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1067),
.A2(n_850),
.B1(n_613),
.B2(n_770),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1072),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_990),
.A2(n_850),
.B(n_770),
.C(n_897),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_950),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_965),
.B(n_597),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_965),
.B(n_597),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_990),
.A2(n_850),
.B(n_770),
.C(n_897),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_974),
.Y(n_1173)
);

AOI221x1_ASAP7_75t_L g1174 ( 
.A1(n_1000),
.A2(n_850),
.B1(n_836),
.B2(n_1042),
.C(n_897),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_963),
.A2(n_885),
.B1(n_770),
.B2(n_903),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1022),
.A2(n_850),
.B1(n_613),
.B2(n_770),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_1036),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1009),
.B(n_980),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_949),
.A2(n_814),
.B(n_1033),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_990),
.B(n_850),
.C(n_897),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1033),
.A2(n_841),
.A3(n_985),
.B(n_1070),
.Y(n_1181)
);

INVxp67_ASAP7_75t_SL g1182 ( 
.A(n_989),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_965),
.B(n_597),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_1033),
.A2(n_958),
.B(n_1022),
.C(n_1042),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1075),
.A2(n_949),
.B(n_1057),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1025),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_1025),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_990),
.A2(n_850),
.B1(n_770),
.B2(n_613),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_950),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1069),
.A2(n_1033),
.B(n_1057),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_950),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_949),
.A2(n_814),
.B(n_1033),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_974),
.B(n_597),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_990),
.B(n_850),
.C(n_897),
.Y(n_1194)
);

OAI22x1_ASAP7_75t_L g1195 ( 
.A1(n_1021),
.A2(n_770),
.B1(n_480),
.B2(n_990),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_990),
.A2(n_850),
.B(n_770),
.C(n_897),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_949),
.A2(n_814),
.B(n_1033),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_988),
.A2(n_1010),
.B(n_1076),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_949),
.A2(n_814),
.B(n_1033),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_1033),
.A2(n_958),
.B(n_1022),
.C(n_1042),
.Y(n_1200)
);

NOR2xp67_ASAP7_75t_L g1201 ( 
.A(n_1015),
.B(n_986),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_990),
.A2(n_850),
.B1(n_770),
.B2(n_613),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1015),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_SL g1204 ( 
.A(n_972),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_L g1205 ( 
.A(n_1015),
.B(n_986),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_990),
.A2(n_770),
.B(n_850),
.C(n_597),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1033),
.A2(n_841),
.A3(n_985),
.B(n_1070),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1025),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_989),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1025),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_988),
.A2(n_1010),
.B(n_1076),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_990),
.A2(n_850),
.B(n_770),
.C(n_897),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_SL g1213 ( 
.A1(n_1033),
.A2(n_958),
.B(n_1022),
.C(n_1042),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_974),
.B(n_597),
.Y(n_1214)
);

O2A1O1Ixp5_ASAP7_75t_SL g1215 ( 
.A1(n_976),
.A2(n_403),
.B(n_1000),
.C(n_1016),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1033),
.A2(n_841),
.A3(n_985),
.B(n_1070),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_1033),
.A2(n_958),
.B(n_1022),
.C(n_1042),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_950),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_965),
.B(n_597),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_990),
.A2(n_850),
.B1(n_770),
.B2(n_613),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_990),
.A2(n_770),
.B(n_850),
.C(n_597),
.Y(n_1221)
);

BUFx8_ASAP7_75t_L g1222 ( 
.A(n_1036),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_988),
.A2(n_1010),
.B(n_1076),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_990),
.A2(n_770),
.B(n_850),
.C(n_597),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_973),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1033),
.A2(n_841),
.A3(n_985),
.B(n_1070),
.Y(n_1226)
);

AO32x2_ASAP7_75t_L g1227 ( 
.A1(n_1000),
.A2(n_631),
.A3(n_971),
.B1(n_961),
.B2(n_498),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_950),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1069),
.A2(n_1033),
.B(n_1077),
.Y(n_1229)
);

AO22x2_ASAP7_75t_L g1230 ( 
.A1(n_1000),
.A2(n_850),
.B1(n_1021),
.B2(n_613),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1173),
.Y(n_1231)
);

BUFx4f_ASAP7_75t_L g1232 ( 
.A(n_1124),
.Y(n_1232)
);

CKINVDCx9p33_ASAP7_75t_R g1233 ( 
.A(n_1109),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1187),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1194),
.A2(n_1180),
.B1(n_1212),
.B2(n_1196),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1178),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1127),
.A2(n_1194),
.B1(n_1176),
.B2(n_1230),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1149),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1168),
.A2(n_1172),
.B(n_1188),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1127),
.A2(n_1230),
.B1(n_1202),
.B2(n_1188),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1202),
.A2(n_1220),
.B1(n_1142),
.B2(n_1166),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1220),
.A2(n_1110),
.B1(n_1195),
.B2(n_1144),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1114),
.A2(n_1174),
.B1(n_1219),
.B2(n_1183),
.Y(n_1243)
);

CKINVDCx12_ASAP7_75t_R g1244 ( 
.A(n_1123),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1178),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1142),
.A2(n_1171),
.B1(n_1170),
.B2(n_1193),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1187),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1101),
.B(n_1116),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1177),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1175),
.A2(n_1118),
.B1(n_1130),
.B2(n_1142),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1187),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1114),
.A2(n_1153),
.B1(n_1117),
.B2(n_1121),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1125),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1102),
.A2(n_1126),
.B1(n_1112),
.B2(n_1199),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1204),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1103),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1189),
.Y(n_1257)
);

INVx6_ASAP7_75t_L g1258 ( 
.A(n_1210),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1214),
.A2(n_1206),
.B1(n_1221),
.B2(n_1224),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1190),
.A2(n_1227),
.B1(n_1197),
.B2(n_1179),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1147),
.A2(n_1145),
.B1(n_1162),
.B2(n_1103),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1191),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1218),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1128),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1119),
.Y(n_1265)
);

INVx6_ASAP7_75t_L g1266 ( 
.A(n_1210),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1141),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1138),
.B(n_1123),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1228),
.Y(n_1269)
);

BUFx2_ASAP7_75t_SL g1270 ( 
.A(n_1129),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1122),
.Y(n_1271)
);

BUFx2_ASAP7_75t_SL g1272 ( 
.A(n_1210),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1137),
.B(n_1106),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1190),
.A2(n_1227),
.B1(n_1192),
.B2(n_1209),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1093),
.A2(n_1229),
.B1(n_1115),
.B2(n_1096),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1164),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1146),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

CKINVDCx14_ASAP7_75t_R g1279 ( 
.A(n_1225),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1138),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1160),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1158),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

BUFx12f_ASAP7_75t_L g1284 ( 
.A(n_1222),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1162),
.A2(n_1131),
.B1(n_1167),
.B2(n_1229),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1154),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1227),
.A2(n_1093),
.B1(n_1135),
.B2(n_1200),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1115),
.A2(n_1136),
.B1(n_1133),
.B2(n_1100),
.Y(n_1288)
);

INVx6_ASAP7_75t_L g1289 ( 
.A(n_1164),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1157),
.A2(n_1159),
.B1(n_1213),
.B2(n_1184),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1095),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1158),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1113),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1107),
.B(n_1155),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1160),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1217),
.A2(n_1222),
.B1(n_1134),
.B2(n_1215),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1143),
.A2(n_1140),
.B1(n_1205),
.B2(n_1201),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_1108),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1152),
.A2(n_1148),
.B(n_1111),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1139),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1161),
.A2(n_1201),
.B1(n_1205),
.B2(n_1108),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1120),
.B(n_1150),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1186),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1208),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1099),
.A2(n_1163),
.B1(n_1151),
.B2(n_1156),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_1203),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1150),
.B(n_1181),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1150),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1098),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_SL g1310 ( 
.A(n_1181),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1104),
.A2(n_1165),
.B1(n_1223),
.B2(n_1211),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1198),
.A2(n_1092),
.B1(n_1226),
.B2(n_1181),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1207),
.B(n_1226),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1207),
.B(n_1226),
.Y(n_1314)
);

BUFx4f_ASAP7_75t_SL g1315 ( 
.A(n_1207),
.Y(n_1315)
);

BUFx2_ASAP7_75t_SL g1316 ( 
.A(n_1097),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1098),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1098),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1216),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1216),
.B(n_1185),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1105),
.A2(n_1202),
.B1(n_1220),
.B2(n_1188),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1132),
.B(n_1094),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1169),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1187),
.Y(n_1324)
);

INVx8_ASAP7_75t_L g1325 ( 
.A(n_1187),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1194),
.A2(n_850),
.B1(n_1180),
.B2(n_1127),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1187),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1169),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1158),
.Y(n_1329)
);

INVx3_ASAP7_75t_SL g1330 ( 
.A(n_1204),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1194),
.A2(n_850),
.B1(n_1180),
.B2(n_1127),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1187),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1093),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1169),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1128),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1095),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1187),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1127),
.A2(n_850),
.B1(n_1194),
.B2(n_1180),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1101),
.B(n_1170),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1188),
.A2(n_1220),
.B1(n_1202),
.B2(n_1114),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1169),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1169),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_1193),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1178),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1128),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1169),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1095),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1169),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1194),
.A2(n_1180),
.B1(n_770),
.B2(n_1172),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1127),
.A2(n_850),
.B1(n_1194),
.B2(n_1180),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1127),
.A2(n_850),
.B1(n_1194),
.B2(n_1180),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1101),
.B(n_1110),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1101),
.B(n_1170),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1308),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1278),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1318),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1313),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1302),
.A2(n_1309),
.A3(n_1317),
.B(n_1235),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1314),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1325),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1340),
.A2(n_1259),
.B1(n_1252),
.B2(n_1331),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1307),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1319),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1322),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1322),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1349),
.A2(n_1333),
.B(n_1294),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1238),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1310),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1333),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1310),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1265),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1247),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1315),
.Y(n_1373)
);

NOR2xp67_ASAP7_75t_SL g1374 ( 
.A(n_1282),
.B(n_1329),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1315),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_1273),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1298),
.Y(n_1377)
);

BUFx12f_ASAP7_75t_L g1378 ( 
.A(n_1284),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1286),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1267),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1287),
.B(n_1338),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1339),
.B(n_1353),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1255),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1271),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1285),
.B(n_1268),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1244),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1271),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1253),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1257),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1291),
.B(n_1300),
.Y(n_1392)
);

AOI211xp5_ASAP7_75t_L g1393 ( 
.A1(n_1340),
.A2(n_1243),
.B(n_1241),
.C(n_1246),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1330),
.Y(n_1394)
);

INVx8_ASAP7_75t_L g1395 ( 
.A(n_1325),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1262),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1263),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1269),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1248),
.B(n_1243),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1352),
.B(n_1326),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1275),
.A2(n_1288),
.B(n_1299),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1277),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1287),
.B(n_1338),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1274),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1254),
.A2(n_1297),
.B(n_1320),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1283),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1274),
.Y(n_1407)
);

CKINVDCx8_ASAP7_75t_R g1408 ( 
.A(n_1270),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1275),
.A2(n_1288),
.B(n_1254),
.Y(n_1409)
);

CKINVDCx9p33_ASAP7_75t_R g1410 ( 
.A(n_1233),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1321),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1316),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1297),
.A2(n_1321),
.B(n_1260),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1312),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1336),
.B(n_1347),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1417)
);

AOI32xp33_ASAP7_75t_L g1418 ( 
.A1(n_1237),
.A2(n_1252),
.A3(n_1250),
.B1(n_1296),
.B2(n_1260),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1312),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1348),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1237),
.B(n_1242),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1323),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1346),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1282),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1328),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1334),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1341),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1250),
.B(n_1342),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1233),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1305),
.A2(n_1301),
.B(n_1290),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1343),
.A2(n_1344),
.B1(n_1236),
.B2(n_1245),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1231),
.B(n_1261),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1290),
.B(n_1296),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1256),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1311),
.A2(n_1304),
.B(n_1303),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1311),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1325),
.B(n_1272),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1306),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1329),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1343),
.B(n_1264),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1335),
.A2(n_1345),
.B(n_1292),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1330),
.B(n_1276),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1361),
.A2(n_1279),
.B1(n_1293),
.B2(n_1280),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1406),
.B(n_1289),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1396),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1376),
.B(n_1281),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1369),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1441),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1396),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1442),
.Y(n_1450)
);

OAI21xp33_ASAP7_75t_L g1451 ( 
.A1(n_1361),
.A2(n_1234),
.B(n_1251),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1393),
.A2(n_1232),
.B(n_1332),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1417),
.B(n_1292),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1387),
.B(n_1281),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1380),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1418),
.A2(n_1232),
.B(n_1234),
.C(n_1251),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1387),
.B(n_1281),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1394),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1413),
.A2(n_1327),
.B(n_1247),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1387),
.B(n_1295),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1405),
.A2(n_1266),
.B(n_1324),
.Y(n_1461)
);

AO32x2_ASAP7_75t_L g1462 ( 
.A1(n_1372),
.A2(n_1295),
.A3(n_1337),
.B1(n_1258),
.B2(n_1266),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1441),
.Y(n_1463)
);

OAI211xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1418),
.A2(n_1249),
.B(n_1337),
.C(n_1258),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1415),
.B(n_1234),
.C(n_1251),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1359),
.B(n_1258),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1415),
.A2(n_1266),
.B(n_1324),
.C(n_1337),
.Y(n_1467)
);

NOR2x1_ASAP7_75t_SL g1468 ( 
.A(n_1363),
.B(n_1324),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1428),
.B(n_1429),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1429),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1359),
.B(n_1355),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1399),
.B(n_1381),
.Y(n_1473)
);

AO32x2_ASAP7_75t_L g1474 ( 
.A1(n_1362),
.A2(n_1366),
.A3(n_1407),
.B1(n_1404),
.B2(n_1419),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1381),
.A2(n_1421),
.B(n_1403),
.C(n_1382),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1430),
.A2(n_1411),
.B(n_1421),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1382),
.A2(n_1403),
.B1(n_1440),
.B2(n_1432),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1386),
.A2(n_1389),
.B(n_1371),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1430),
.A2(n_1411),
.B(n_1366),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1362),
.B(n_1379),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1363),
.B(n_1425),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1433),
.A2(n_1383),
.B(n_1400),
.C(n_1363),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1441),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1433),
.A2(n_1434),
.B(n_1426),
.C(n_1389),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1412),
.A2(n_1371),
.B(n_1384),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1363),
.B(n_1408),
.Y(n_1487)
);

AO32x2_ASAP7_75t_L g1488 ( 
.A1(n_1404),
.A2(n_1407),
.A3(n_1419),
.B1(n_1414),
.B2(n_1358),
.Y(n_1488)
);

AOI211xp5_ASAP7_75t_L g1489 ( 
.A1(n_1388),
.A2(n_1436),
.B(n_1414),
.C(n_1438),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1408),
.A2(n_1431),
.B1(n_1377),
.B2(n_1384),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1438),
.B(n_1375),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1357),
.B(n_1391),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1436),
.A2(n_1435),
.B(n_1354),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1375),
.B(n_1368),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1390),
.B(n_1397),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1378),
.A2(n_1368),
.B1(n_1375),
.B2(n_1385),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1378),
.A2(n_1368),
.B1(n_1416),
.B2(n_1392),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1360),
.B(n_1395),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1445),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1493),
.B(n_1409),
.Y(n_1500)
);

AND2x2_ASAP7_75t_SL g1501 ( 
.A(n_1482),
.B(n_1401),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1448),
.B(n_1463),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1449),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1488),
.B(n_1484),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1473),
.B(n_1386),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1484),
.Y(n_1506)
);

AOI21xp33_ASAP7_75t_L g1507 ( 
.A1(n_1464),
.A2(n_1409),
.B(n_1401),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1488),
.B(n_1401),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1488),
.B(n_1401),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1471),
.B(n_1369),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1462),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1474),
.B(n_1356),
.Y(n_1512)
);

NAND4xp25_ASAP7_75t_L g1513 ( 
.A(n_1456),
.B(n_1422),
.C(n_1420),
.D(n_1423),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1480),
.B(n_1447),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1447),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1486),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1356),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1495),
.B(n_1358),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1358),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1474),
.B(n_1358),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1464),
.A2(n_1386),
.B1(n_1367),
.B2(n_1368),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1458),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1492),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1479),
.B(n_1358),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1492),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1473),
.B(n_1358),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_L g1527 ( 
.A(n_1478),
.B(n_1364),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1467),
.A2(n_1412),
.B(n_1424),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1476),
.B(n_1398),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1526),
.B(n_1476),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1526),
.B(n_1485),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1512),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1481),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1512),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1521),
.A2(n_1483),
.B1(n_1475),
.B2(n_1477),
.C(n_1452),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1515),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1516),
.A2(n_1490),
.B1(n_1489),
.B2(n_1451),
.C(n_1485),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1450),
.Y(n_1540)
);

OAI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1507),
.A2(n_1443),
.B(n_1452),
.C(n_1459),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1523),
.B(n_1491),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1455),
.Y(n_1543)
);

OAI222xp33_ASAP7_75t_L g1544 ( 
.A1(n_1521),
.A2(n_1490),
.B1(n_1487),
.B2(n_1497),
.C1(n_1496),
.C2(n_1469),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1522),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1500),
.A2(n_1365),
.B(n_1459),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1523),
.B(n_1491),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1499),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1499),
.Y(n_1549)
);

OAI211xp5_ASAP7_75t_L g1550 ( 
.A1(n_1507),
.A2(n_1461),
.B(n_1467),
.C(n_1465),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1513),
.A2(n_1453),
.B1(n_1461),
.B2(n_1470),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1529),
.B(n_1374),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1522),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1510),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1512),
.Y(n_1555)
);

AOI221xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1513),
.A2(n_1453),
.B1(n_1446),
.B2(n_1457),
.C(n_1454),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1499),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1503),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1503),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1502),
.B(n_1512),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1531),
.Y(n_1561)
);

OAI33xp33_ASAP7_75t_L g1562 ( 
.A1(n_1530),
.A2(n_1446),
.A3(n_1402),
.B1(n_1420),
.B2(n_1427),
.B3(n_1423),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1517),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1518),
.B(n_1466),
.Y(n_1564)
);

OAI31xp33_ASAP7_75t_L g1565 ( 
.A1(n_1516),
.A2(n_1460),
.A3(n_1410),
.B(n_1494),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1517),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1502),
.B(n_1472),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1548),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1560),
.B(n_1504),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1548),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1528),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1545),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1504),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1549),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1560),
.B(n_1504),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1560),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_L g1578 ( 
.A(n_1532),
.B(n_1528),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1532),
.B(n_1518),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1567),
.B(n_1504),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1557),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1561),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1534),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1533),
.B(n_1523),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1542),
.B(n_1525),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1567),
.B(n_1535),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1501),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1542),
.B(n_1525),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1536),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1537),
.A2(n_1509),
.B1(n_1508),
.B2(n_1519),
.C(n_1520),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1556),
.B(n_1505),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1558),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1559),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1550),
.B(n_1527),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1559),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1547),
.B(n_1506),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1501),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1538),
.Y(n_1599)
);

NOR3xp33_ASAP7_75t_SL g1600 ( 
.A(n_1544),
.B(n_1529),
.C(n_1530),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1571),
.B(n_1556),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1586),
.B(n_1540),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1568),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1594),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1586),
.B(n_1540),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1571),
.B(n_1551),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1600),
.A2(n_1537),
.B1(n_1551),
.B2(n_1539),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1591),
.B(n_1539),
.Y(n_1608)
);

AOI32xp33_ASAP7_75t_L g1609 ( 
.A1(n_1590),
.A2(n_1509),
.A3(n_1508),
.B1(n_1524),
.B2(n_1520),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1572),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1568),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1583),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1598),
.B(n_1567),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1598),
.B(n_1555),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1569),
.B(n_1555),
.Y(n_1617)
);

O2A1O1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1600),
.A2(n_1594),
.B(n_1541),
.C(n_1590),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1597),
.B(n_1564),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1569),
.B(n_1555),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1572),
.A2(n_1541),
.B1(n_1501),
.B2(n_1552),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_L g1623 ( 
.A1(n_1572),
.A2(n_1550),
.B1(n_1562),
.B2(n_1509),
.C1(n_1508),
.C2(n_1524),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1583),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1583),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1570),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1570),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1574),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1569),
.B(n_1563),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1574),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1573),
.B(n_1563),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1576),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1597),
.B(n_1564),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1576),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1578),
.B(n_1565),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1581),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1582),
.B(n_1545),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1573),
.B(n_1563),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1578),
.A2(n_1552),
.B(n_1565),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1581),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1573),
.B(n_1566),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1579),
.B(n_1554),
.Y(n_1642)
);

NOR3xp33_ASAP7_75t_SL g1643 ( 
.A(n_1607),
.B(n_1553),
.C(n_1595),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1604),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1620),
.B(n_1579),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1608),
.B(n_1610),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1603),
.Y(n_1648)
);

NAND3x1_ASAP7_75t_L g1649 ( 
.A(n_1639),
.B(n_1577),
.C(n_1575),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1618),
.B(n_1545),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1603),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1611),
.Y(n_1652)
);

INVxp33_ASAP7_75t_L g1653 ( 
.A(n_1637),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1602),
.B(n_1575),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1605),
.B(n_1614),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1606),
.A2(n_1552),
.B(n_1546),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1605),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1611),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1575),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1626),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1601),
.B(n_1582),
.Y(n_1661)
);

XNOR2xp5_ASAP7_75t_L g1662 ( 
.A(n_1622),
.B(n_1444),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1635),
.B(n_1580),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1585),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1612),
.Y(n_1665)
);

AND4x1_ASAP7_75t_L g1666 ( 
.A(n_1623),
.B(n_1498),
.C(n_1374),
.D(n_1587),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1580),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1612),
.A2(n_1577),
.B(n_1589),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1626),
.Y(n_1670)
);

OAI31xp33_ASAP7_75t_L g1671 ( 
.A1(n_1642),
.A2(n_1582),
.A3(n_1524),
.B(n_1587),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1627),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1627),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_L g1674 ( 
.A1(n_1609),
.A2(n_1524),
.B(n_1509),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1620),
.B(n_1585),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1616),
.B(n_1619),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1615),
.B(n_1577),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1664),
.A2(n_1609),
.B1(n_1628),
.B2(n_1640),
.C(n_1632),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1648),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

AO22x1_ASAP7_75t_L g1681 ( 
.A1(n_1650),
.A2(n_1612),
.B1(n_1628),
.B2(n_1640),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1651),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1650),
.B(n_1633),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1643),
.A2(n_1508),
.B(n_1520),
.C(n_1519),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1645),
.B(n_1633),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1651),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

NOR3xp33_ASAP7_75t_SL g1688 ( 
.A(n_1647),
.B(n_1636),
.C(n_1634),
.Y(n_1688)
);

OAI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1666),
.A2(n_1642),
.B(n_1632),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1588),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1652),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1658),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1655),
.B(n_1617),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1655),
.B(n_1663),
.Y(n_1695)
);

NAND2xp33_ASAP7_75t_L g1696 ( 
.A(n_1649),
.B(n_1395),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1660),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1674),
.A2(n_1520),
.B(n_1519),
.C(n_1527),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1660),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1644),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1670),
.Y(n_1702)
);

NOR2xp67_ASAP7_75t_SL g1703 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1678),
.A2(n_1674),
.B1(n_1653),
.B2(n_1673),
.C(n_1672),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1695),
.B(n_1644),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1693),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1679),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1695),
.B(n_1701),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1685),
.B(n_1662),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1681),
.A2(n_1662),
.B(n_1670),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1680),
.Y(n_1711)
);

O2A1O1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1689),
.A2(n_1666),
.B(n_1671),
.C(n_1673),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1700),
.B(n_1657),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1688),
.B(n_1657),
.Y(n_1714)
);

OAI31xp33_ASAP7_75t_L g1715 ( 
.A1(n_1684),
.A2(n_1649),
.A3(n_1676),
.B(n_1646),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1682),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1688),
.B(n_1654),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1684),
.A2(n_1654),
.B1(n_1659),
.B2(n_1646),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1690),
.B(n_1667),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1696),
.A2(n_1659),
.B1(n_1546),
.B2(n_1677),
.Y(n_1720)
);

OAI31xp33_ASAP7_75t_L g1721 ( 
.A1(n_1698),
.A2(n_1675),
.A3(n_1677),
.B(n_1667),
.Y(n_1721)
);

XNOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1708),
.B(n_1686),
.Y(n_1722)
);

AO21x1_ASAP7_75t_L g1723 ( 
.A1(n_1710),
.A2(n_1696),
.B(n_1691),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1715),
.A2(n_1698),
.B1(n_1699),
.B2(n_1702),
.C(n_1697),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1709),
.B(n_1687),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1705),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1713),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1707),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1717),
.Y(n_1730)
);

XOR2xp5_ASAP7_75t_L g1731 ( 
.A(n_1710),
.B(n_1468),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1711),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1714),
.B(n_1694),
.Y(n_1733)
);

AOI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1723),
.A2(n_1703),
.B(n_1722),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1728),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1728),
.B(n_1704),
.Y(n_1736)
);

NAND3xp33_ASAP7_75t_L g1737 ( 
.A(n_1724),
.B(n_1704),
.C(n_1712),
.Y(n_1737)
);

NAND4xp75_ASAP7_75t_L g1738 ( 
.A(n_1729),
.B(n_1721),
.C(n_1716),
.D(n_1720),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1729),
.Y(n_1739)
);

NAND4xp25_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_1718),
.C(n_1672),
.D(n_1668),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1730),
.B(n_1675),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1722),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1737),
.A2(n_1742),
.B(n_1736),
.C(n_1740),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1734),
.A2(n_1731),
.B1(n_1726),
.B2(n_1727),
.C(n_1733),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1742),
.A2(n_1732),
.B(n_1727),
.C(n_1665),
.Y(n_1745)
);

OAI211xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1741),
.A2(n_1665),
.B(n_1668),
.C(n_1612),
.Y(n_1746)
);

AOI211x1_ASAP7_75t_SL g1747 ( 
.A1(n_1738),
.A2(n_1625),
.B(n_1613),
.C(n_1624),
.Y(n_1747)
);

OAI211xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1743),
.A2(n_1735),
.B(n_1739),
.C(n_1665),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1744),
.B(n_1745),
.Y(n_1749)
);

NAND4xp25_ASAP7_75t_SL g1750 ( 
.A(n_1747),
.B(n_1634),
.C(n_1636),
.D(n_1630),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1746),
.A2(n_1630),
.B1(n_1613),
.B2(n_1625),
.C(n_1624),
.Y(n_1751)
);

AOI211x1_ASAP7_75t_SL g1752 ( 
.A1(n_1746),
.A2(n_1625),
.B(n_1624),
.C(n_1589),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1745),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1753),
.B(n_1617),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1750),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1748),
.B(n_1599),
.Y(n_1756)
);

XNOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1749),
.B(n_1437),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1752),
.B(n_1621),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1754),
.B(n_1751),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1755),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_L g1761 ( 
.A(n_1756),
.B(n_1669),
.C(n_1360),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1757),
.B1(n_1758),
.B2(n_1669),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1759),
.B1(n_1761),
.B2(n_1641),
.Y(n_1763)
);

XNOR2xp5_ASAP7_75t_L g1764 ( 
.A(n_1763),
.B(n_1437),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1638),
.B1(n_1631),
.B2(n_1629),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1765),
.Y(n_1766)
);

AOI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1599),
.B1(n_1592),
.B2(n_1596),
.C(n_1593),
.Y(n_1767)
);

INVxp67_ASAP7_75t_SL g1768 ( 
.A(n_1766),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1588),
.B(n_1595),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1767),
.B(n_1360),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1395),
.B(n_1631),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1769),
.Y(n_1772)
);

OAI221xp5_ASAP7_75t_R g1773 ( 
.A1(n_1772),
.A2(n_1395),
.B1(n_1629),
.B2(n_1621),
.C(n_1638),
.Y(n_1773)
);

AOI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1771),
.B(n_1424),
.C(n_1439),
.Y(n_1774)
);


endmodule