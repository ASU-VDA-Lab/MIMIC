module fake_jpeg_8114_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_62),
.B(n_53),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_68),
.B(n_75),
.C(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_0),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_64),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_2),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_79),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_63),
.B1(n_48),
.B2(n_65),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_17),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_60),
.B1(n_58),
.B2(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_88),
.B1(n_81),
.B2(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_94),
.B1(n_90),
.B2(n_91),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_92),
.B1(n_55),
.B2(n_52),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_76),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_19),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_21),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_24),
.B(n_26),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_27),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_28),
.B(n_30),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_105)
);

AOI321xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_37),
.A3(n_39),
.B1(n_40),
.B2(n_42),
.C(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_81),
.Y(n_107)
);


endmodule