module fake_jpeg_30024_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_52),
.Y(n_146)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_55),
.Y(n_144)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_88),
.Y(n_125)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_72),
.Y(n_112)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_21),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_43),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_10),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_10),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_92),
.B(n_103),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

CKINVDCx6p67_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_33),
.B(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_39),
.Y(n_128)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g109 ( 
.A(n_101),
.Y(n_109)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_102),
.B(n_51),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_42),
.B(n_8),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_53),
.B(n_18),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_110),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_131),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_41),
.B1(n_51),
.B2(n_44),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_124),
.A2(n_142),
.B1(n_68),
.B2(n_83),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_133),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_158),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_43),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_34),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_34),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_70),
.A2(n_41),
.B1(n_49),
.B2(n_42),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_74),
.A2(n_41),
.B1(n_28),
.B2(n_37),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_100),
.B1(n_101),
.B2(n_97),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_52),
.B(n_49),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_95),
.B(n_48),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_54),
.A2(n_28),
.B1(n_31),
.B2(n_37),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_81),
.B1(n_75),
.B2(n_66),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_76),
.B(n_48),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_35),
.Y(n_188)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_172),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_173),
.A2(n_164),
.B1(n_162),
.B2(n_153),
.Y(n_252)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_174),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_176),
.Y(n_264)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_179),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_180),
.B(n_182),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_107),
.B(n_63),
.C(n_59),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_189),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_115),
.Y(n_182)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

CKINVDCx6p67_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_186),
.B(n_188),
.Y(n_271)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_113),
.A2(n_94),
.B1(n_93),
.B2(n_91),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_198),
.B1(n_124),
.B2(n_150),
.Y(n_230)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_200),
.Y(n_232)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_129),
.A2(n_87),
.B1(n_60),
.B2(n_82),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_55),
.C(n_80),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_225),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_109),
.A2(n_85),
.B1(n_62),
.B2(n_61),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_201),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_32),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_207),
.Y(n_233)
);

CKINVDCx6p67_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_203),
.Y(n_250)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_32),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_217),
.Y(n_238)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_116),
.Y(n_210)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_159),
.A2(n_35),
.B(n_71),
.C(n_72),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_151),
.B(n_134),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_151),
.B1(n_162),
.B2(n_150),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_108),
.B(n_64),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_228),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_218),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_154),
.A2(n_51),
.B1(n_44),
.B2(n_37),
.Y(n_219)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_105),
.B(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_222),
.Y(n_239)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_112),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_226),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_154),
.A2(n_37),
.B1(n_31),
.B2(n_2),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_224),
.A2(n_164),
.B1(n_143),
.B2(n_167),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_149),
.B(n_31),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_31),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_112),
.B(n_11),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_130),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_230),
.B(n_234),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_241),
.A2(n_252),
.B1(n_257),
.B2(n_201),
.Y(n_306)
);

NOR2x1_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_147),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_242),
.B(n_251),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_169),
.B(n_171),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_183),
.A2(n_146),
.B(n_167),
.C(n_143),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_258),
.B(n_261),
.Y(n_297)
);

OR2x2_ASAP7_75t_SL g259 ( 
.A(n_170),
.B(n_155),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_226),
.C(n_225),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_19),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_179),
.B(n_19),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_265),
.Y(n_286)
);

AOI32xp33_ASAP7_75t_L g265 ( 
.A1(n_194),
.A2(n_165),
.A3(n_167),
.B1(n_130),
.B2(n_139),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_212),
.A2(n_153),
.B1(n_139),
.B2(n_19),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_199),
.B(n_0),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_170),
.B(n_0),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_284),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_173),
.B1(n_189),
.B2(n_190),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_283),
.A2(n_290),
.B1(n_303),
.B2(n_310),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_203),
.B1(n_175),
.B2(n_205),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_287),
.A2(n_318),
.B1(n_322),
.B2(n_243),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_181),
.B1(n_219),
.B2(n_190),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_288),
.B(n_311),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_289),
.B(n_266),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_234),
.A2(n_198),
.B1(n_184),
.B2(n_206),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_204),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g365 ( 
.A(n_292),
.B(n_273),
.CI(n_255),
.CON(n_365),
.SN(n_365)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_238),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_308),
.Y(n_346)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_174),
.C(n_218),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_301),
.C(n_305),
.Y(n_329)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_222),
.C(n_209),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_230),
.A2(n_198),
.B1(n_220),
.B2(n_203),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_304),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_268),
.C(n_245),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_306),
.A2(n_265),
.B(n_240),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_263),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_320),
.Y(n_335)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_245),
.A2(n_195),
.A3(n_192),
.B1(n_185),
.B2(n_176),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_235),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_312),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_268),
.A2(n_215),
.B1(n_197),
.B2(n_229),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_230),
.A2(n_224),
.B1(n_191),
.B2(n_193),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_313),
.B(n_319),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_185),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_316),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_242),
.A2(n_196),
.B1(n_3),
.B2(n_4),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_315),
.A2(n_255),
.B1(n_247),
.B2(n_256),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_233),
.B(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_239),
.B(n_217),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_321),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_253),
.A2(n_217),
.B1(n_19),
.B2(n_5),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_233),
.B(n_1),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_250),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_232),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_293),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_258),
.B(n_1),
.C(n_3),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_278),
.C(n_277),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_266),
.B(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_325),
.B(n_281),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_241),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_252),
.B1(n_250),
.B2(n_235),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_328),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_330),
.A2(n_321),
.B1(n_296),
.B2(n_285),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_363),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_339),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_305),
.B(n_230),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_282),
.A2(n_286),
.B(n_297),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_366),
.B(n_324),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_317),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_342),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_295),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_343),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_316),
.B(n_260),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_354),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_263),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_314),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_282),
.A2(n_272),
.B(n_247),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_350),
.A2(n_351),
.B(n_355),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_283),
.A2(n_254),
.B1(n_243),
.B2(n_231),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_282),
.A2(n_254),
.B1(n_243),
.B2(n_264),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_302),
.A2(n_272),
.B(n_264),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_302),
.A2(n_260),
.B1(n_231),
.B2(n_236),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_328),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_256),
.B1(n_267),
.B2(n_236),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_309),
.B1(n_299),
.B2(n_320),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_300),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_360),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_278),
.B1(n_277),
.B2(n_273),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_365),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_323),
.A2(n_244),
.B(n_6),
.Y(n_366)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_371),
.B(n_365),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_298),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_384),
.C(n_399),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_375),
.Y(n_427)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_362),
.Y(n_376)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_332),
.B(n_291),
.Y(n_378)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_378),
.B(n_401),
.C(n_377),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_336),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_382),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_344),
.A2(n_288),
.B1(n_301),
.B2(n_315),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_381),
.B1(n_383),
.B2(n_391),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_344),
.A2(n_308),
.B1(n_294),
.B2(n_292),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_327),
.B(n_292),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_350),
.A2(n_326),
.B(n_289),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_385),
.A2(n_355),
.B(n_349),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_319),
.B(n_313),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_386),
.A2(n_398),
.B(n_366),
.Y(n_412)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_346),
.A2(n_342),
.B1(n_354),
.B2(n_340),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_393),
.A2(n_395),
.B1(n_396),
.B2(n_400),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_346),
.A2(n_312),
.B1(n_304),
.B2(n_244),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_340),
.A2(n_5),
.B1(n_8),
.B2(n_11),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

AOI32xp33_ASAP7_75t_L g398 ( 
.A1(n_339),
.A2(n_8),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_329),
.B(n_12),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_330),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_L g401 ( 
.A1(n_332),
.A2(n_12),
.B(n_14),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_329),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_429),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_378),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_405),
.B(n_398),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_387),
.A2(n_357),
.B1(n_352),
.B2(n_345),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_406),
.A2(n_411),
.B1(n_425),
.B2(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_345),
.Y(n_408)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_368),
.B(n_384),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_426),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_387),
.A2(n_347),
.B1(n_363),
.B2(n_331),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_412),
.A2(n_421),
.B1(n_375),
.B2(n_394),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_353),
.Y(n_413)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_358),
.Y(n_419)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_419),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_SL g436 ( 
.A(n_420),
.B(n_373),
.C(n_377),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_361),
.B1(n_337),
.B2(n_335),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_388),
.B(n_348),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_428),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_358),
.Y(n_424)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_380),
.A2(n_364),
.B1(n_361),
.B2(n_337),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_368),
.B(n_334),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_356),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_430),
.B(n_396),
.Y(n_454)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_392),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_372),
.Y(n_445)
);

BUFx12_ASAP7_75t_L g433 ( 
.A(n_420),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_439),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_399),
.C(n_369),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_438),
.C(n_449),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_436),
.A2(n_427),
.B(n_413),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_418),
.A2(n_394),
.B(n_389),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_417),
.B(n_416),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_369),
.C(n_386),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_441),
.A2(n_448),
.B1(n_436),
.B2(n_456),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_443),
.B(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_406),
.A2(n_425),
.B1(n_394),
.B2(n_418),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_419),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_414),
.A2(n_367),
.B1(n_372),
.B2(n_373),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_385),
.C(n_367),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_402),
.B(n_400),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_451),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_408),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_456),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_343),
.Y(n_455)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_364),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_360),
.Y(n_457)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_411),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_465),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_470),
.B(n_455),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_478),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_410),
.C(n_427),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_440),
.C(n_450),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_430),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_445),
.Y(n_466)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_466),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_467),
.A2(n_474),
.B1(n_477),
.B2(n_437),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_404),
.Y(n_468)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_433),
.A2(n_424),
.B(n_414),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_453),
.A2(n_381),
.B1(n_417),
.B2(n_412),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_440),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_458),
.A2(n_407),
.B1(n_426),
.B2(n_422),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_364),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_407),
.Y(n_479)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_479),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_484),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_434),
.B1(n_439),
.B2(n_447),
.Y(n_482)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_482),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_463),
.B(n_444),
.Y(n_483)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_472),
.A2(n_433),
.B(n_457),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_475),
.A2(n_448),
.B(n_458),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_488),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_490),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_461),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_492),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_474),
.A2(n_446),
.B1(n_454),
.B2(n_338),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_467),
.A2(n_364),
.B1(n_338),
.B2(n_370),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_478),
.Y(n_509)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_497),
.A2(n_466),
.B1(n_480),
.B2(n_471),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_501),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_489),
.A2(n_480),
.B1(n_462),
.B2(n_477),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_500),
.A2(n_505),
.B1(n_507),
.B2(n_496),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_463),
.C(n_460),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_487),
.B(n_497),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_495),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_494),
.A2(n_493),
.B1(n_496),
.B2(n_488),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_494),
.A2(n_476),
.B1(n_468),
.B2(n_479),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_490),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_491),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_493),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_512),
.A2(n_518),
.B1(n_509),
.B2(n_504),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_516),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g524 ( 
.A1(n_515),
.A2(n_517),
.B(n_521),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_499),
.A2(n_506),
.B(n_511),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_510),
.A2(n_459),
.B1(n_465),
.B2(n_485),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_484),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_519),
.A2(n_520),
.B(n_464),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_502),
.B(n_481),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_508),
.A2(n_470),
.B1(n_397),
.B2(n_459),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_501),
.C(n_504),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_525),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_521),
.A2(n_508),
.B(n_505),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_517),
.B(n_515),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_526),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_530),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_527),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_514),
.C(n_500),
.Y(n_533)
);

AOI211xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_531),
.B(n_524),
.C(n_359),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_524),
.Y(n_535)
);

CKINVDCx14_ASAP7_75t_R g536 ( 
.A(n_535),
.Y(n_536)
);

AOI221xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_532),
.B1(n_359),
.B2(n_397),
.C(n_17),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_537),
.B(n_16),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_16),
.B(n_17),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_16),
.B(n_18),
.Y(n_540)
);


endmodule