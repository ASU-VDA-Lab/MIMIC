module fake_netlist_6_3944_n_178 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_178);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_178;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_85;
wire n_99;
wire n_66;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVxp33_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_R g50 ( 
.A(n_7),
.B(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_3),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_4),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_32),
.B(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_51),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_51),
.B(n_34),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_50),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_53),
.B(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_43),
.B1(n_47),
.B2(n_25),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_43),
.B(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_28),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_67),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_58),
.B1(n_72),
.B2(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_57),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_59),
.B(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx2_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_74),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_84),
.B(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_85),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_82),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_94),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_78),
.B(n_80),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_94),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_91),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_92),
.B(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_96),
.B1(n_105),
.B2(n_109),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_122),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_112),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_122),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_119),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_113),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_75),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_77),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_133),
.Y(n_142)
);

NOR4xp75_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_125),
.C(n_66),
.D(n_101),
.Y(n_143)
);

OAI211xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_64),
.B(n_132),
.C(n_60),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_128),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_63),
.C(n_129),
.Y(n_146)
);

OAI221xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_60),
.B1(n_66),
.B2(n_56),
.C(n_127),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_127),
.B(n_115),
.C(n_133),
.Y(n_148)
);

NOR3x1_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_101),
.C(n_56),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_87),
.C(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND4xp75_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_143),
.C(n_130),
.D(n_57),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_58),
.C(n_130),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_123),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_62),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_62),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_155),
.B1(n_152),
.B2(n_153),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_58),
.C(n_108),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_104),
.B1(n_108),
.B2(n_92),
.C(n_103),
.Y(n_169)
);

NAND5xp2_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_109),
.C(n_103),
.D(n_104),
.E(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_163),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_109),
.C(n_93),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_109),
.B1(n_103),
.B2(n_93),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_160),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_167),
.B1(n_161),
.B2(n_100),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_167),
.C(n_172),
.Y(n_177)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_175),
.B1(n_170),
.B2(n_174),
.C(n_173),
.Y(n_178)
);


endmodule