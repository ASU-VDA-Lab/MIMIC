module fake_jpeg_10220_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_48),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_47),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_8),
.B1(n_15),
.B2(n_13),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_41),
.B(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_24),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_18),
.B1(n_35),
.B2(n_19),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_66),
.B1(n_38),
.B2(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_70),
.Y(n_76)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_67),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_34),
.B(n_18),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_73),
.A2(n_83),
.B1(n_50),
.B2(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_81),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_87),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_25),
.B1(n_47),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_91),
.B1(n_26),
.B2(n_20),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_20),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_47),
.B1(n_53),
.B2(n_39),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_102),
.B1(n_100),
.B2(n_77),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_40),
.B1(n_66),
.B2(n_64),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx10_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_84),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_50),
.B1(n_35),
.B2(n_26),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_128),
.B1(n_21),
.B2(n_90),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_125),
.B1(n_120),
.B2(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_50),
.B1(n_26),
.B2(n_21),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_87),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_132),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_131),
.A2(n_136),
.B1(n_105),
.B2(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_99),
.B1(n_78),
.B2(n_80),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_133),
.A2(n_31),
.B1(n_23),
.B2(n_32),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_93),
.Y(n_137)
);

CKINVDCx12_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_139),
.B(n_31),
.C(n_23),
.Y(n_186)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_93),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_87),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_83),
.B1(n_94),
.B2(n_77),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_147),
.B1(n_119),
.B2(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_83),
.B1(n_74),
.B2(n_97),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_28),
.Y(n_149)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_155),
.Y(n_187)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_103),
.B(n_29),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_32),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_28),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_28),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_159),
.A2(n_162),
.B(n_163),
.Y(n_213)
);

AO21x2_ASAP7_75t_SL g160 ( 
.A1(n_135),
.A2(n_112),
.B(n_56),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_132),
.B(n_138),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_33),
.B(n_109),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_37),
.B(n_33),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_164),
.B(n_180),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_31),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_150),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_145),
.B1(n_136),
.B2(n_143),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_172),
.B1(n_176),
.B2(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_126),
.B1(n_110),
.B2(n_116),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_127),
.B1(n_104),
.B2(n_105),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_179),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_137),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_183),
.C(n_188),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_115),
.B1(n_114),
.B2(n_112),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_56),
.B1(n_29),
.B2(n_55),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_186),
.B1(n_158),
.B2(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_28),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_131),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_55),
.B(n_57),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_141),
.A2(n_55),
.B1(n_71),
.B2(n_95),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_152),
.B1(n_141),
.B2(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_57),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_199),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_155),
.B(n_151),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_205),
.B1(n_179),
.B2(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_200),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_153),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_32),
.Y(n_234)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_152),
.B1(n_71),
.B2(n_23),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_163),
.B1(n_184),
.B2(n_32),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_32),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_211),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_58),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_212),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_173),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_188),
.C(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_217),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_95),
.C(n_58),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_159),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_181),
.B1(n_189),
.B2(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_222),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_215),
.B(n_182),
.CI(n_180),
.CON(n_222),
.SN(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_227),
.A2(n_237),
.B1(n_239),
.B2(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_232),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_186),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_229),
.B(n_230),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_206),
.B(n_162),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_231),
.A2(n_200),
.B1(n_213),
.B2(n_10),
.Y(n_268)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_0),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_194),
.B(n_201),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_243),
.B(n_246),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_216),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_9),
.B(n_15),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_9),
.B(n_12),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_9),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_196),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_214),
.C(n_212),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_267),
.C(n_235),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_257),
.B(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_203),
.B(n_192),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_210),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_231),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_198),
.B(n_194),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_266),
.A2(n_268),
.B1(n_237),
.B2(n_239),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_214),
.C(n_191),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_225),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.C(n_278),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_225),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_226),
.C(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_226),
.C(n_222),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_222),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_248),
.A2(n_241),
.B1(n_227),
.B2(n_234),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_271),
.B1(n_282),
.B2(n_283),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_258),
.B(n_243),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_257),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_248),
.B1(n_254),
.B2(n_255),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_270),
.B1(n_280),
.B2(n_252),
.Y(n_305)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_300),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_250),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_278),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_253),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_8),
.B(n_12),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_249),
.B(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_263),
.B1(n_268),
.B2(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_276),
.B1(n_256),
.B2(n_259),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_11),
.B1(n_16),
.B2(n_6),
.Y(n_315)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_256),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_10),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_311),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_305),
.B1(n_307),
.B2(n_296),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_288),
.A2(n_274),
.B1(n_233),
.B2(n_246),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_297),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_229),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_313),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_233),
.B1(n_10),
.B2(n_11),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_11),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_307),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_321),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_295),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_299),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_324),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_292),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_294),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_315),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_16),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_330),
.C(n_7),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_308),
.C(n_312),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_320),
.A3(n_16),
.B1(n_6),
.B2(n_7),
.C1(n_4),
.C2(n_3),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_321),
.B(n_316),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_329),
.B(n_327),
.C(n_335),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_336),
.B(n_326),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_7),
.Y(n_343)
);


endmodule