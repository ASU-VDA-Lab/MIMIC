module real_jpeg_535_n_7 (n_5, n_4, n_39, n_0, n_40, n_43, n_1, n_41, n_2, n_38, n_6, n_42, n_3, n_7);

input n_5;
input n_4;
input n_39;
input n_0;
input n_40;
input n_43;
input n_1;
input n_41;
input n_2;
input n_38;
input n_6;
input n_42;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_13),
.C(n_29),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

FAx1_ASAP7_75t_SL g7 ( 
.A(n_3),
.B(n_8),
.CI(n_11),
.CON(n_7),
.SN(n_7)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_5),
.A2(n_20),
.B(n_23),
.Y(n_19)
);

AO22x1_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_14),
.B1(n_18),
.B2(n_28),
.Y(n_13)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_32),
.C(n_33),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_17),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.C(n_27),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_26),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_38),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_39),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_40),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_41),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_42),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_43),
.Y(n_35)
);


endmodule