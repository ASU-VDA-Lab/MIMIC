module fake_jpeg_1875_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_1),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_51),
.B1(n_56),
.B2(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_61),
.B1(n_57),
.B2(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_53),
.B1(n_50),
.B2(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_53),
.B1(n_49),
.B2(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_64),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_89),
.Y(n_101)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_16),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_86),
.B1(n_48),
.B2(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_41),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_61),
.B1(n_60),
.B2(n_43),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_46),
.B(n_52),
.C(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_68),
.B1(n_73),
.B2(n_59),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_104),
.B1(n_105),
.B2(n_8),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_100),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_9),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_1),
.C(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_2),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_22),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_6),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_121),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_88),
.C(n_24),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_118),
.C(n_29),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_117),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_8),
.B(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_34),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_25),
.C(n_38),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_11),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_13),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_131),
.B1(n_134),
.B2(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_14),
.B1(n_21),
.B2(n_27),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_39),
.C(n_111),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_138),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_145),
.B1(n_137),
.B2(n_127),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_112),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_126),
.B(n_132),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_144),
.A2(n_139),
.B1(n_119),
.B2(n_131),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_142),
.C(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_140),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_154),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_107),
.C(n_131),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_129),
.Y(n_162)
);


endmodule