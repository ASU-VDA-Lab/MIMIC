module fake_jpeg_10069_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_38),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.C(n_1),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_26),
.C(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_50),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_26),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_24),
.B1(n_22),
.B2(n_31),
.Y(n_93)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_21),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_34),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_68),
.B(n_38),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_34),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_21),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_37),
.B(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_32),
.B1(n_38),
.B2(n_37),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_86),
.B(n_95),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_74),
.B(n_58),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_25),
.B1(n_34),
.B2(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_55),
.B1(n_48),
.B2(n_53),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_44),
.A3(n_42),
.B1(n_28),
.B2(n_25),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_58),
.C(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_40),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_92),
.C(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_42),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_24),
.B1(n_18),
.B2(n_31),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_47),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_55),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_40),
.B1(n_25),
.B2(n_18),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_108),
.B(n_85),
.Y(n_144)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_106),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_86),
.Y(n_146)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_120),
.B1(n_82),
.B2(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_110),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_113),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_46),
.B1(n_60),
.B2(n_31),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_123),
.B(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_122),
.B1(n_126),
.B2(n_84),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_46),
.C(n_63),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_77),
.C(n_47),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_60),
.B1(n_70),
.B2(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_28),
.B1(n_20),
.B2(n_33),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_71),
.B(n_86),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_127),
.A2(n_143),
.B(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_133),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_85),
.C(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_134),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_15),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_20),
.B(n_30),
.C(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_113),
.B(n_116),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.C(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_152),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_106),
.B(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_170),
.B(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_164),
.C(n_165),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_115),
.B1(n_117),
.B2(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_175),
.B1(n_181),
.B2(n_153),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_108),
.C(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_129),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_144),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_103),
.C(n_123),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_103),
.A3(n_47),
.B1(n_28),
.B2(n_20),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_87),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_101),
.B1(n_78),
.B2(n_30),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_27),
.B(n_33),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_44),
.C(n_35),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_149),
.C(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_177),
.B1(n_138),
.B2(n_141),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_101),
.B1(n_78),
.B2(n_97),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2x1_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_44),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_97),
.B1(n_76),
.B2(n_124),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_173),
.B(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_152),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_206),
.B1(n_170),
.B2(n_156),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_180),
.A3(n_146),
.B1(n_150),
.B2(n_171),
.C1(n_178),
.C2(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_154),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_191),
.B1(n_199),
.B2(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_44),
.C(n_136),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_140),
.B1(n_138),
.B2(n_131),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_208),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_151),
.B1(n_139),
.B2(n_130),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_153),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_2),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_181),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_178),
.B1(n_162),
.B2(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_203),
.A2(n_205),
.B1(n_193),
.B2(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_134),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_166),
.A2(n_146),
.B1(n_133),
.B2(n_136),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_146),
.C(n_44),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_27),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_155),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_175),
.B1(n_165),
.B2(n_167),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_216),
.B1(n_218),
.B2(n_231),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_214),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_204),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_232),
.B1(n_186),
.B2(n_188),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_156),
.B(n_179),
.C(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_220),
.C(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_64),
.C(n_41),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_76),
.B1(n_118),
.B2(n_33),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_64),
.C(n_41),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_118),
.B1(n_67),
.B2(n_33),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_189),
.B1(n_194),
.B2(n_198),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_201),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_118),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_27),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_233),
.C(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_30),
.B1(n_20),
.B2(n_4),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_30),
.B1(n_27),
.B2(n_4),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_27),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_235),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_196),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_247),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_188),
.B1(n_189),
.B2(n_202),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_256),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_248),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_209),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_203),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_190),
.C(n_27),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_190),
.C(n_27),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_30),
.B1(n_16),
.B2(n_15),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_226),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_212),
.B1(n_217),
.B2(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_211),
.B(n_234),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_14),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_259),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_266),
.Y(n_278)
);

AO221x1_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_223),
.B1(n_212),
.B2(n_230),
.C(n_232),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_243),
.B(n_229),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_253),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_225),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_271),
.Y(n_280)
);

AO22x1_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_223),
.B1(n_227),
.B2(n_219),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_233),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_267),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_240),
.B(n_247),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_236),
.C(n_246),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_281),
.C(n_271),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_245),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_251),
.B1(n_244),
.B2(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_288),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_285),
.A2(n_290),
.B1(n_2),
.B2(n_3),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_16),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_267),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_275),
.B1(n_260),
.B2(n_268),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_303),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_275),
.B1(n_264),
.B2(n_258),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_271),
.B(n_270),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_12),
.B(n_13),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_278),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_285),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_5),
.C(n_6),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_6),
.C(n_7),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_311),
.B(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_277),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_7),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_306),
.B(n_312),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_13),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_305),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_14),
.C(n_8),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_299),
.B(n_297),
.C(n_291),
.D(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_317),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_316),
.B(n_318),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_302),
.B1(n_297),
.B2(n_9),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_8),
.C(n_9),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_7),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_324),
.A2(n_325),
.B(n_9),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_8),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_319),
.B(n_9),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_322),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_10),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_10),
.Y(n_332)
);


endmodule