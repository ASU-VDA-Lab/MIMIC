module fake_jpeg_17951_n_387 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_39),
.B(n_49),
.Y(n_80)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_13),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_62),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_52),
.B(n_60),
.Y(n_116)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_65),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_68),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_11),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_10),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_71),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_32),
.B1(n_34),
.B2(n_16),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_74),
.A2(n_76),
.B1(n_89),
.B2(n_94),
.Y(n_140)
);

BUFx2_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2x1_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_37),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_34),
.B1(n_24),
.B2(n_32),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_86),
.B(n_95),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_32),
.B1(n_20),
.B2(n_31),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_37),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g144 ( 
.A(n_91),
.B(n_37),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_33),
.B1(n_35),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_93),
.A2(n_112),
.B1(n_115),
.B2(n_37),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_24),
.B1(n_35),
.B2(n_38),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_38),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_97),
.B(n_7),
.Y(n_173)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_18),
.B(n_28),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_99),
.A2(n_2),
.B(n_4),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_48),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_20),
.B1(n_31),
.B2(n_30),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_56),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_123),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_40),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_118),
.Y(n_171)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_44),
.A2(n_23),
.B1(n_2),
.B2(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_57),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_124),
.A2(n_155),
.B(n_172),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_121),
.B1(n_106),
.B2(n_90),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_126),
.A2(n_169),
.B1(n_87),
.B2(n_113),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_1),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_127),
.A2(n_87),
.B1(n_8),
.B2(n_88),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_18),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_138),
.Y(n_183)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

BUFx2_ASAP7_75t_SL g130 ( 
.A(n_83),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_130),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_133),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_132),
.A2(n_160),
.B(n_163),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_77),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_136),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_84),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_137),
.B(n_142),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_28),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_SL g142 ( 
.A(n_75),
.B(n_45),
.C(n_9),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_173),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_28),
.B1(n_18),
.B2(n_37),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_28),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_156),
.Y(n_196)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_150),
.B(n_153),
.Y(n_201)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_45),
.Y(n_154)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_18),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_18),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_88),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_80),
.B(n_9),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_127),
.B1(n_156),
.B2(n_8),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_9),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_165),
.C(n_96),
.Y(n_186)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_78),
.B(n_5),
.C(n_6),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_110),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_120),
.C(n_115),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_186),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_111),
.B1(n_112),
.B2(n_85),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_187),
.B1(n_193),
.B2(n_204),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_194),
.A2(n_206),
.B(n_207),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_96),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_208),
.C(n_176),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_199),
.B(n_217),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_161),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_155),
.A2(n_147),
.B1(n_145),
.B2(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_151),
.B1(n_149),
.B2(n_164),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_127),
.A2(n_92),
.B1(n_105),
.B2(n_88),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_144),
.B(n_92),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_165),
.C(n_168),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_194),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_131),
.B(n_105),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_162),
.A2(n_103),
.B(n_159),
.C(n_124),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_162),
.A2(n_103),
.B1(n_134),
.B2(n_137),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_139),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_162),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_238),
.Y(n_261)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_141),
.B(n_129),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_222),
.A2(n_223),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_175),
.B(n_135),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_229),
.Y(n_276)
);

BUFx24_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_175),
.B(n_125),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_167),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_232),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_167),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_234),
.B(n_254),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_141),
.B1(n_171),
.B2(n_148),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_236),
.B1(n_246),
.B2(n_252),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_196),
.A2(n_171),
.B1(n_152),
.B2(n_143),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_182),
.C(n_219),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_198),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_239),
.B(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_195),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_243),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_247),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_218),
.A2(n_191),
.B1(n_187),
.B2(n_198),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_206),
.B(n_189),
.C(n_207),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_243),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_202),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_183),
.A2(n_208),
.B1(n_193),
.B2(n_204),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_189),
.A2(n_176),
.B1(n_197),
.B2(n_210),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_253),
.A2(n_255),
.B1(n_237),
.B2(n_222),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_189),
.A2(n_197),
.B1(n_210),
.B2(n_190),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_203),
.B(n_180),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_228),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

OAI22x1_ASAP7_75t_SL g259 ( 
.A1(n_249),
.A2(n_192),
.B1(n_177),
.B2(n_205),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_227),
.B1(n_266),
.B2(n_260),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_272),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_256),
.B(n_249),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_263),
.A2(n_277),
.B(n_267),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_185),
.B(n_188),
.Y(n_266)
);

AO22x2_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_273),
.B1(n_288),
.B2(n_270),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_225),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_225),
.C(n_241),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_256),
.C(n_252),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_220),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_287),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_297),
.C(n_298),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_272),
.A2(n_223),
.B1(n_246),
.B2(n_234),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_248),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_251),
.C(n_236),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_263),
.A2(n_223),
.B1(n_250),
.B2(n_227),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_304),
.B1(n_313),
.B2(n_314),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_309),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_267),
.A2(n_277),
.B(n_273),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_289),
.C(n_277),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_286),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_266),
.B1(n_285),
.B2(n_289),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_261),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_286),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_266),
.B1(n_281),
.B2(n_265),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_317),
.A2(n_327),
.B1(n_336),
.B2(n_292),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_334),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_316),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_298),
.C(n_293),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_314),
.A2(n_294),
.B1(n_299),
.B2(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_328),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_295),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_331),
.B(n_332),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_308),
.B(n_276),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_333),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_280),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_310),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_341),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_319),
.B(n_305),
.CI(n_309),
.CON(n_340),
.SN(n_340)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_319),
.B(n_314),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_342),
.B(n_345),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_312),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_344),
.C(n_347),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_291),
.C(n_293),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_330),
.A2(n_302),
.B1(n_294),
.B2(n_311),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_315),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_318),
.A2(n_283),
.B1(n_287),
.B2(n_275),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_353),
.B1(n_321),
.B2(n_325),
.Y(n_354)
);

AOI211xp5_ASAP7_75t_SL g353 ( 
.A1(n_322),
.A2(n_297),
.B(n_264),
.C(n_276),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_354),
.A2(n_351),
.B1(n_341),
.B2(n_324),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_348),
.A2(n_324),
.B(n_335),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_357),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_329),
.C(n_325),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_329),
.C(n_321),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_361),
.B(n_363),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_318),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_353),
.B(n_352),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_317),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_336),
.C(n_262),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_347),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_337),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_372),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_362),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_371),
.C(n_355),
.Y(n_377)
);

AO22x1_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_340),
.B1(n_346),
.B2(n_349),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_357),
.C(n_365),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_369),
.A2(n_364),
.B(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_376),
.Y(n_379)
);

AOI322xp5_ASAP7_75t_L g380 ( 
.A1(n_377),
.A2(n_366),
.A3(n_371),
.B1(n_355),
.B2(n_359),
.C1(n_372),
.C2(n_358),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_374),
.B(n_375),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_382),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_350),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_383),
.B(n_379),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_384),
.A2(n_346),
.B1(n_375),
.B2(n_290),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_262),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g387 ( 
.A(n_386),
.B(n_290),
.CI(n_335),
.CON(n_387),
.SN(n_387)
);


endmodule