module fake_jpeg_25971_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_15),
.B1(n_10),
.B2(n_8),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g13 ( 
.A1(n_11),
.A2(n_1),
.B(n_2),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_15),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_8),
.B1(n_10),
.B2(n_6),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.C(n_22),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_17),
.B1(n_16),
.B2(n_7),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_14),
.C(n_3),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_28),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.C(n_29),
.Y(n_33)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_28),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_3),
.B(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_14),
.Y(n_36)
);


endmodule