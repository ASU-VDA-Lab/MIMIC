module real_jpeg_6154_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_0),
.A2(n_61),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_0),
.A2(n_61),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_0),
.A2(n_61),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_1),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_1),
.Y(n_187)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_1),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_1),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_1),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_2),
.A2(n_269),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_2),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_2),
.A2(n_189),
.B1(n_293),
.B2(n_307),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_2),
.A2(n_293),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_2),
.A2(n_53),
.B1(n_293),
.B2(n_464),
.Y(n_463)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_3),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_3),
.Y(n_250)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_3),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_4),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_4),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_4),
.A2(n_128),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_128),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_4),
.A2(n_128),
.B1(n_424),
.B2(n_427),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_5),
.A2(n_58),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_5),
.A2(n_80),
.B1(n_208),
.B2(n_269),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_5),
.A2(n_182),
.B1(n_208),
.B2(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_5),
.A2(n_208),
.B1(n_344),
.B2(n_346),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_79),
.B1(n_137),
.B2(n_163),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_137),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_20),
.B(n_510),
.Y(n_19)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_8),
.Y(n_512)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_13),
.A2(n_199),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_13),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_13),
.B(n_82),
.C(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_13),
.B(n_118),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_13),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_13),
.B(n_93),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_13),
.B(n_134),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_14),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_15),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_15),
.A2(n_251),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_15),
.A2(n_79),
.B1(n_251),
.B2(n_334),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_15),
.A2(n_172),
.B1(n_251),
.B2(n_439),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_16),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_16),
.A2(n_44),
.B1(n_98),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_16),
.A2(n_98),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_18),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_18),
.A2(n_51),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_18),
.A2(n_51),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_18),
.A2(n_51),
.B1(n_238),
.B2(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_211),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_210),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_156),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_24),
.B(n_156),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_138),
.B2(n_139),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.C(n_99),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_27),
.A2(n_140),
.B1(n_141),
.B2(n_155),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_27),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_27),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_28),
.A2(n_55),
.B1(n_57),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_28),
.A2(n_248),
.B(n_253),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_28),
.A2(n_39),
.B1(n_248),
.B2(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_29),
.B(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_29),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_39),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_35),
.Y(n_154)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_39),
.B(n_266),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_39)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_40),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_42),
.Y(n_345)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_42),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_43),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_43),
.Y(n_414)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_44),
.A2(n_404),
.A3(n_407),
.B1(n_409),
.B2(n_415),
.Y(n_403)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_45),
.Y(n_136)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_48),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_50),
.B(n_56),
.Y(n_205)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_52),
.Y(n_406)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_55),
.A2(n_206),
.B(n_463),
.Y(n_480)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_56),
.B(n_207),
.Y(n_253)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_59),
.A2(n_266),
.B(n_415),
.Y(n_434)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_60),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_63),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_62),
.A2(n_63),
.B1(n_99),
.B2(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_92),
.B(n_94),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_64),
.A2(n_264),
.B(n_267),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_64),
.A2(n_92),
.B1(n_291),
.B2(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_64),
.A2(n_267),
.B(n_333),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_64),
.A2(n_92),
.B1(n_444),
.B2(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_65),
.A2(n_93),
.B1(n_162),
.B2(n_167),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_65),
.A2(n_93),
.B1(n_162),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_65),
.A2(n_93),
.B1(n_198),
.B2(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_65),
.B(n_268),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_81),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_75),
.B2(n_79),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_70),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_70),
.Y(n_203)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_70),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_70),
.Y(n_273)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_71),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_71),
.Y(n_365)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_81),
.A2(n_291),
.B(n_294),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_88),
.B2(n_90),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_86),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_88),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_88),
.Y(n_427)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_92),
.A2(n_294),
.B(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_93),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_97),
.Y(n_445)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_125),
.B1(n_132),
.B2(n_133),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_132),
.B1(n_133),
.B2(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_101),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_101),
.A2(n_132),
.B1(n_171),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_101),
.A2(n_132),
.B1(n_379),
.B2(n_438),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_118),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_108),
.B1(n_111),
.B2(n_113),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_105),
.Y(n_362)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_107),
.Y(n_368)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_110),
.Y(n_442)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_117),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_117),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_117),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_118),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_126),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22x1_ASAP7_75t_L g466 ( 
.A1(n_118),
.A2(n_169),
.B1(n_385),
.B2(n_467),
.Y(n_466)
);

AO22x2_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_121),
.Y(n_238)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_131),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_132),
.B(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_132),
.A2(n_379),
.B(n_384),
.Y(n_378)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_176),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_157),
.B(n_160),
.CI(n_176),
.CON(n_213),
.SN(n_213)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_166),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_169),
.A2(n_338),
.B(n_342),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_169),
.B(n_385),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_169),
.A2(n_342),
.B(n_483),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_174),
.Y(n_380)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B(n_204),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_197),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_204),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_178),
.A2(n_197),
.B1(n_219),
.B2(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_185),
.B(n_188),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_188),
.B1(n_226),
.B2(n_232),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_179),
.A2(n_278),
.B(n_283),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_179),
.A2(n_266),
.B(n_283),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_179),
.A2(n_418),
.B1(n_419),
.B2(n_422),
.Y(n_417)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_180),
.B(n_286),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_180),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_180),
.A2(n_352),
.B1(n_389),
.B2(n_394),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_180),
.A2(n_186),
.B1(n_423),
.B2(n_460),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_181),
.Y(n_322)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_191),
.Y(n_282)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_191),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_197),
.Y(n_454)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_254),
.B(n_509),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_213),
.B(n_214),
.Y(n_509)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_213),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.C(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_220),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_223),
.B(n_469),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_242),
.C(n_247),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_224),
.B(n_452),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_236),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_225),
.B(n_236),
.Y(n_477)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_226),
.Y(n_460)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_229),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_229),
.Y(n_391)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_235),
.Y(n_421)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_237),
.Y(n_458)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_242),
.B(n_247),
.Y(n_452)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_243),
.Y(n_467)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_250),
.B(n_266),
.Y(n_415)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_253),
.Y(n_435)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI311xp33_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_448),
.A3(n_485),
.B1(n_503),
.C1(n_504),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_397),
.B(n_447),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_370),
.B(n_396),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_327),
.B(n_369),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_297),
.B(n_326),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_276),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_262),
.B(n_276),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_271),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_263),
.A2(n_271),
.B1(n_272),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g338 ( 
.A1(n_266),
.A2(n_339),
.B(n_340),
.Y(n_338)
);

INVx3_ASAP7_75t_SL g360 ( 
.A(n_269),
.Y(n_360)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_289),
.C(n_296),
.Y(n_328)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_285),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_295),
.B2(n_296),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_316),
.B(n_325),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_304),
.B(n_315),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_314),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_314),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_310),
.B(n_313),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_313),
.A2(n_351),
.B(n_357),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_323),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_329),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_349),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_336),
.B2(n_337),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_336),
.C(n_349),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI32xp33_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_359),
.A3(n_360),
.B1(n_361),
.B2(n_363),
.Y(n_358)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_358),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_358),
.Y(n_376)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_371),
.B(n_372),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_377),
.B2(n_395),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_376),
.C(n_395),
.Y(n_398)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_386),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_378),
.B(n_387),
.C(n_388),
.Y(n_428)
);

INVx4_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_398),
.B(n_399),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_431),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_400)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_401),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_416),
.B2(n_417),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_403),
.B(n_416),
.Y(n_481)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx6_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_428),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_429),
.C(n_431),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_436),
.B2(n_446),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_432),
.B(n_437),
.C(n_443),
.Y(n_494)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_436),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_443),
.Y(n_436)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_471),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_SL g504 ( 
.A1(n_449),
.A2(n_471),
.B(n_505),
.C(n_508),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_468),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_450),
.B(n_468),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_453),
.C(n_455),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_451),
.B(n_453),
.CI(n_455),
.CON(n_484),
.SN(n_484)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_461),
.C(n_466),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_459),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_461),
.A2(n_462),
.B1(n_466),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_466),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_484),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_477),
.C(n_478),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.C(n_482),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_480),
.B1(n_482),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_484),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_498),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_487),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_495),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_495),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_492),
.C(n_494),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_501),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_492),
.A2(n_493),
.B1(n_494),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_500),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

INVx8_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);


endmodule