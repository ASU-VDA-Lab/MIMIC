module fake_netlist_6_1629_n_2047 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2047);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2047;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_59),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_53),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_50),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_18),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_51),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_7),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_77),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_84),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_75),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_125),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_39),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_65),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_103),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_168),
.Y(n_238)
);

CKINVDCx6p67_ASAP7_75t_R g239 ( 
.A(n_94),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_202),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_134),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_43),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_92),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_133),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_107),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_98),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_73),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_69),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_70),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_88),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_85),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_172),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_70),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_67),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_74),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_163),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_108),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_193),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_191),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_176),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_9),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_137),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_29),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_12),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_26),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_49),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_158),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_148),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_29),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_106),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_113),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_194),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_24),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_138),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_102),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_82),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_16),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_71),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_184),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_157),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_129),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_11),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_60),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_95),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_39),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_128),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_54),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_209),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_182),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_112),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_23),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_131),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_150),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_33),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_25),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_109),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_87),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_104),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_199),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_42),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_81),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_166),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_34),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_208),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_51),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_105),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_27),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_111),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_142),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_155),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_40),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_79),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_200),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_74),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_89),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_159),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_195),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_54),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_167),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_47),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_120),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_205),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_210),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_136),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_114),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_119),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_207),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_21),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_32),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_57),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_122),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_96),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_147),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_139),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_196),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_68),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_6),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_115),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_14),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_156),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_66),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_56),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_154),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_72),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_68),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_110),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_58),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_83),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_161),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_31),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_30),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_153),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_90),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_43),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_40),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_183),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_143),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_23),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_197),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_31),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_20),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_162),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_35),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_3),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_28),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_80),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_3),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_15),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_86),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_24),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_180),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_97),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_4),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_35),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_37),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_164),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_49),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_146),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_132),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_22),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_56),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_149),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_190),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_5),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_62),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_0),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_101),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_64),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_124),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_14),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_71),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_192),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_173),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_4),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_16),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_38),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_46),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_45),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_185),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_188),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_32),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_212),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_255),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_257),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_212),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_212),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_215),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_212),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_262),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_263),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_264),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_398),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_265),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_267),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_212),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_269),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_320),
.B(n_222),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_212),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_229),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_212),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_211),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_212),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_240),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_246),
.B(n_0),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_284),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_290),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_293),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_219),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_274),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_278),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_335),
.B(n_1),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_311),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_396),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_1),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_353),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_353),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_214),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_353),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_383),
.B(n_2),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_408),
.B(n_2),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_251),
.B(n_6),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_358),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_280),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_281),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_344),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_285),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_292),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_294),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_251),
.B(n_7),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_369),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_298),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_258),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_300),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_273),
.B(n_8),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_244),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_372),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_372),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_258),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_372),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_273),
.B(n_8),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_415),
.B(n_10),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_307),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_322),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_324),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_326),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_327),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_258),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_213),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_356),
.B(n_10),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_379),
.B(n_12),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_221),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_227),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_224),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_332),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_242),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_356),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_334),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_214),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_338),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_248),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_252),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_234),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_254),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_216),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_247),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_249),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_339),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_341),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_482),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_228),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_461),
.B(n_356),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_223),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_243),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_420),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_228),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_434),
.A2(n_310),
.B1(n_385),
.B2(n_288),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_482),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_419),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_422),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_223),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_509),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_452),
.A2(n_397),
.B1(n_414),
.B2(n_411),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_490),
.B(n_275),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_275),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_291),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_491),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_291),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_495),
.B(n_225),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_495),
.B(n_317),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_497),
.B(n_225),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_460),
.B(n_391),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_497),
.B(n_317),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_423),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_425),
.B(n_318),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_425),
.B(n_318),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_499),
.B(n_330),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_432),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_435),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_435),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_437),
.B(n_230),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_439),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_468),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_440),
.B(n_453),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_454),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_454),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_455),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_455),
.B(n_330),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_515),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_456),
.A2(n_289),
.B(n_282),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_499),
.B(n_342),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_457),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_457),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_459),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_521),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_342),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_459),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_464),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_467),
.Y(n_588)
);

AND3x2_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_393),
.C(n_321),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_467),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_476),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_479),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_479),
.Y(n_594)
);

AND3x2_ASAP7_75t_L g595 ( 
.A(n_446),
.B(n_393),
.C(n_325),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_504),
.B(n_253),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

INVx6_ASAP7_75t_L g598 ( 
.A(n_473),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_489),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_481),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_483),
.Y(n_601)
);

BUFx8_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_483),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_484),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_484),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_505),
.B(n_256),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_429),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_486),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_486),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_498),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_554),
.A2(n_424),
.B1(n_473),
.B2(n_474),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_596),
.B(n_259),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_536),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_570),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_537),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_554),
.B(n_421),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_529),
.B(n_426),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_557),
.A2(n_279),
.B(n_276),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_570),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_570),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_529),
.B(n_427),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_537),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_533),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_592),
.B(n_428),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_537),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_537),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_556),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_592),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_592),
.B(n_430),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_599),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_560),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_540),
.B(n_431),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_537),
.Y(n_639)
);

AND3x2_ASAP7_75t_L g640 ( 
.A(n_607),
.B(n_502),
.C(n_485),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_536),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_527),
.B(n_243),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_560),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_540),
.B(n_433),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_598),
.B(n_506),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_578),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_538),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_567),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_561),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_596),
.B(n_505),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_538),
.Y(n_655)
);

INVx6_ASAP7_75t_L g656 ( 
.A(n_541),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_598),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_538),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_596),
.B(n_480),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_598),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_607),
.B(n_447),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_564),
.B(n_527),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_537),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_564),
.B(n_527),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_545),
.A2(n_463),
.B1(n_449),
.B2(n_442),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_448),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_538),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_607),
.B(n_465),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_577),
.B(n_466),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_606),
.B(n_503),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_577),
.B(n_469),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_552),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_606),
.B(n_520),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_545),
.B(n_470),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_552),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_565),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_565),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_542),
.A2(n_271),
.B1(n_367),
.B2(n_268),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_606),
.B(n_283),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_571),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_598),
.B(n_287),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_568),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_568),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_598),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_568),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_568),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_571),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_578),
.A2(n_462),
.B1(n_472),
.B2(n_478),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_602),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_559),
.B(n_304),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_528),
.B(n_493),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_568),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_528),
.B(n_494),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_578),
.A2(n_488),
.B1(n_492),
.B2(n_458),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_572),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_574),
.B(n_500),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_552),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_598),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_574),
.B(n_511),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_580),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_580),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_544),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_583),
.B(n_525),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_581),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_557),
.B(n_243),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_548),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_581),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_582),
.B(n_303),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g716 ( 
.A(n_544),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_567),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_562),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_580),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_582),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_583),
.B(n_477),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_602),
.B(n_475),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_562),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_562),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_546),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_559),
.B(n_520),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_589),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_585),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_550),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_585),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_586),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_550),
.B(n_243),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_578),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_602),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_578),
.A2(n_316),
.B1(n_394),
.B2(n_384),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_559),
.B(n_584),
.C(n_579),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_553),
.B(n_496),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_586),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_562),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_580),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_557),
.A2(n_331),
.B1(n_403),
.B2(n_380),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_526),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_580),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_602),
.B(n_471),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_526),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_548),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_526),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_580),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_542),
.A2(n_524),
.B1(n_516),
.B2(n_514),
.Y(n_750)
);

AND2x6_ASAP7_75t_L g751 ( 
.A(n_557),
.B(n_243),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_553),
.B(n_501),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_590),
.Y(n_753)
);

BUFx6f_ASAP7_75t_SL g754 ( 
.A(n_557),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_526),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_314),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_548),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_526),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_535),
.B(n_471),
.C(n_513),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_546),
.B(n_216),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_535),
.A2(n_296),
.B1(n_295),
.B2(n_337),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_546),
.B(n_510),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_591),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_636),
.B(n_579),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_662),
.B(n_591),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_664),
.B(n_594),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_617),
.B(n_594),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_623),
.B(n_603),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_614),
.B(n_602),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_729),
.B(n_589),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_646),
.B(n_603),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_725),
.B(n_604),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_631),
.Y(n_773)
);

AND2x6_ASAP7_75t_SL g774 ( 
.A(n_721),
.B(n_345),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_631),
.Y(n_775)
);

INVx8_ASAP7_75t_L g776 ( 
.A(n_684),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_633),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_616),
.A2(n_752),
.B1(n_738),
.B2(n_697),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_614),
.B(n_541),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_693),
.B(n_604),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_633),
.B(n_605),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_634),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_626),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_637),
.B(n_605),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_637),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_619),
.Y(n_786)
);

AND2x6_ASAP7_75t_SL g787 ( 
.A(n_699),
.B(n_346),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_609),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_643),
.B(n_343),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_645),
.B(n_609),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_650),
.B(n_548),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_548),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_653),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_619),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_666),
.A2(n_445),
.B1(n_450),
.B2(n_451),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_653),
.B(n_587),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_643),
.B(n_348),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_667),
.B(n_587),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_737),
.B(n_657),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_634),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_620),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_626),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_659),
.B(n_579),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_659),
.B(n_584),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_636),
.B(n_584),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_762),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_667),
.B(n_587),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_672),
.B(n_587),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_672),
.B(n_587),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_762),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_620),
.B(n_541),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_678),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_665),
.B(n_595),
.C(n_261),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_676),
.B(n_404),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_621),
.B(n_624),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_621),
.B(n_541),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_624),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_648),
.B(n_541),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_716),
.B(n_436),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_745),
.B(n_354),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_647),
.A2(n_441),
.B1(n_444),
.B2(n_443),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_726),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_700),
.A2(n_360),
.B1(n_373),
.B2(n_374),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_648),
.B(n_541),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_680),
.B(n_593),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_726),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_SL g830 ( 
.A1(n_734),
.A2(n_575),
.B(n_558),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_680),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_734),
.A2(n_558),
.B1(n_575),
.B2(n_378),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_683),
.B(n_593),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_683),
.B(n_593),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_692),
.B(n_593),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_692),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_695),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_695),
.B(n_593),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_671),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_703),
.B(n_600),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_600),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_702),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_654),
.B(n_391),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_671),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_706),
.B(n_600),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_675),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_675),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_711),
.B(n_600),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_627),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_734),
.A2(n_375),
.B(n_371),
.C(n_412),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_711),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_652),
.B(n_510),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_714),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_714),
.Y(n_854)
);

NOR2x1p5_ASAP7_75t_L g855 ( 
.A(n_694),
.B(n_239),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_720),
.B(n_600),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_632),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_720),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_753),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_728),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_647),
.A2(n_558),
.B1(n_575),
.B2(n_352),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_753),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_728),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_731),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_732),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_732),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_709),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_739),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_739),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_687),
.B(n_541),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_763),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_687),
.B(n_541),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_687),
.B(n_558),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_763),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_694),
.B(n_239),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_753),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_654),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_713),
.B(n_558),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_747),
.B(n_575),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_709),
.B(n_717),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_757),
.B(n_575),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_737),
.B(n_580),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_657),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_628),
.B(n_601),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_635),
.B(n_601),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_696),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_612),
.B(n_601),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_709),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_709),
.B(n_391),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_612),
.B(n_601),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_638),
.B(n_230),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_612),
.B(n_601),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_612),
.B(n_601),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_670),
.B(n_231),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_660),
.B(n_305),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_682),
.B(n_601),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_733),
.A2(n_566),
.B(n_539),
.Y(n_897)
);

INVx8_ASAP7_75t_L g898 ( 
.A(n_684),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_696),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_673),
.B(n_512),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_710),
.B(n_231),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_750),
.B(n_611),
.C(n_681),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_761),
.B(n_517),
.C(n_512),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_615),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_696),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_727),
.B(n_233),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_682),
.B(n_539),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_660),
.B(n_266),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_715),
.A2(n_566),
.B(n_539),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_705),
.B(n_266),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_647),
.A2(n_727),
.B1(n_682),
.B2(n_754),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_682),
.B(n_696),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_615),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_743),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_756),
.B(n_566),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_743),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_736),
.B(n_643),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_705),
.B(n_308),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_615),
.B(n_266),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_684),
.A2(n_608),
.B(n_597),
.C(n_569),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_746),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_643),
.B(n_569),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_613),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_759),
.B(n_517),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_615),
.B(n_629),
.Y(n_925)
);

AND2x6_ASAP7_75t_SL g926 ( 
.A(n_647),
.B(n_518),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_L g927 ( 
.A(n_735),
.B(n_661),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_760),
.B(n_742),
.C(n_647),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_643),
.B(n_625),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_643),
.B(n_573),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_613),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_622),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_746),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_684),
.A2(n_409),
.B1(n_312),
.B2(n_365),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_830),
.A2(n_685),
.B(n_644),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_808),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_873),
.A2(n_685),
.B(n_644),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_804),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_873),
.A2(n_685),
.B(n_644),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_876),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_882),
.A2(n_685),
.B(n_644),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_767),
.B(n_625),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_783),
.B(n_735),
.Y(n_943)
);

AO21x1_ASAP7_75t_L g944 ( 
.A1(n_778),
.A2(n_618),
.B(n_333),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_786),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_768),
.A2(n_684),
.B1(n_754),
.B2(n_722),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_795),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_876),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_805),
.B(n_669),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_771),
.B(n_625),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_816),
.B(n_765),
.Y(n_951)
);

OAI321xp33_ASAP7_75t_L g952 ( 
.A1(n_816),
.A2(n_355),
.A3(n_329),
.B1(n_336),
.B2(n_340),
.C(n_386),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_766),
.B(n_625),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_806),
.B(n_639),
.Y(n_954)
);

AOI21x1_ASAP7_75t_L g955 ( 
.A1(n_820),
.A2(n_655),
.B(n_651),
.Y(n_955)
);

AO21x1_ASAP7_75t_L g956 ( 
.A1(n_826),
.A2(n_410),
.B(n_395),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_902),
.A2(n_417),
.B(n_518),
.C(n_250),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_827),
.A2(n_658),
.B(n_655),
.Y(n_958)
);

NOR2x1_ASAP7_75t_L g959 ( 
.A(n_880),
.B(n_639),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_827),
.A2(n_668),
.B(n_658),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_884),
.A2(n_885),
.B(n_780),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_812),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_912),
.A2(n_879),
.B(n_878),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_764),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_852),
.Y(n_965)
);

O2A1O1Ixp5_ASAP7_75t_L g966 ( 
.A1(n_840),
.A2(n_718),
.B(n_677),
.C(n_674),
.Y(n_966)
);

BUFx8_ASAP7_75t_L g967 ( 
.A(n_821),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_840),
.B(n_639),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_772),
.B(n_640),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_845),
.B(n_639),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_770),
.B(n_754),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_801),
.B(n_649),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_774),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_862),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_845),
.B(n_649),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_776),
.B(n_498),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_850),
.A2(n_723),
.B(n_674),
.C(n_668),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_770),
.B(n_649),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_881),
.A2(n_719),
.B(n_691),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_907),
.A2(n_719),
.B(n_691),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_817),
.A2(n_701),
.B(n_677),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_803),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_801),
.A2(n_712),
.B1(n_751),
.B2(n_698),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_801),
.B(n_649),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_832),
.A2(n_679),
.B1(n_686),
.B2(n_749),
.Y(n_985)
);

AND2x4_ASAP7_75t_SL g986 ( 
.A(n_862),
.B(n_534),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_887),
.A2(n_629),
.B(n_615),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_890),
.A2(n_663),
.B(n_629),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_807),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_850),
.A2(n_724),
.B(n_704),
.C(n_718),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_892),
.A2(n_663),
.B(n_629),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_849),
.B(n_758),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_893),
.A2(n_663),
.B(n_629),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_859),
.B(n_851),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_924),
.B(n_679),
.Y(n_995)
);

BUFx2_ASAP7_75t_SL g996 ( 
.A(n_867),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_896),
.A2(n_690),
.B(n_663),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_928),
.A2(n_405),
.B(n_250),
.C(n_245),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_819),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_817),
.A2(n_740),
.B(n_723),
.C(n_724),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_859),
.B(n_853),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_915),
.A2(n_690),
.B(n_663),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_925),
.A2(n_690),
.B(n_686),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_925),
.A2(n_690),
.B(n_686),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_779),
.A2(n_704),
.B(n_701),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_886),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_L g1007 ( 
.A(n_796),
.B(n_237),
.C(n_233),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_SL g1008 ( 
.A1(n_917),
.A2(n_740),
.B(n_755),
.C(n_748),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_870),
.A2(n_872),
.B(n_929),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_832),
.A2(n_686),
.B(n_679),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_791),
.A2(n_688),
.B(n_679),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_773),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_782),
.Y(n_1013)
);

AO21x1_ASAP7_75t_L g1014 ( 
.A1(n_769),
.A2(n_543),
.B(n_534),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_911),
.A2(n_688),
.B1(n_689),
.B2(n_749),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_872),
.A2(n_689),
.B(n_688),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_854),
.B(n_688),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_862),
.B(n_689),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_802),
.A2(n_920),
.B(n_793),
.Y(n_1019)
);

AOI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_891),
.A2(n_270),
.B(n_260),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_793),
.A2(n_707),
.B(n_698),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_860),
.B(n_698),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_865),
.A2(n_913),
.B(n_904),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_862),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_926),
.Y(n_1025)
);

O2A1O1Ixp5_ASAP7_75t_L g1026 ( 
.A1(n_909),
.A2(n_707),
.B(n_741),
.C(n_744),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_863),
.B(n_707),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_866),
.B(n_730),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_868),
.B(n_869),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_792),
.A2(n_741),
.B(n_730),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_857),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_775),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_775),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_871),
.B(n_730),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_843),
.B(n_595),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_904),
.A2(n_741),
.B(n_730),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_L g1037 ( 
.A(n_857),
.B(n_741),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_777),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_877),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_861),
.A2(n_744),
.B1(n_749),
.B2(n_238),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_782),
.B(n_744),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_785),
.B(n_744),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_839),
.B(n_749),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_785),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_906),
.B(n_844),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_899),
.A2(n_416),
.B1(n_238),
.B2(n_241),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_904),
.A2(n_708),
.B(n_630),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_794),
.B(n_622),
.Y(n_1048)
);

CKINVDCx10_ASAP7_75t_R g1049 ( 
.A(n_822),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_798),
.A2(n_809),
.B(n_800),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_900),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_814),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_906),
.B(n_272),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_822),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_846),
.B(n_748),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_891),
.B(n_286),
.C(n_277),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_814),
.B(n_755),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_822),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_782),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_824),
.B(n_758),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_888),
.B(n_349),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_904),
.A2(n_708),
.B(n_630),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_824),
.B(n_641),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_889),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_905),
.A2(n_237),
.B1(n_241),
.B2(n_315),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_847),
.B(n_217),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_SL g1067 ( 
.A1(n_810),
.A2(n_642),
.B(n_532),
.C(n_547),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_823),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_782),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_831),
.B(n_573),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_894),
.B(n_350),
.Y(n_1071)
);

OAI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_825),
.A2(n_235),
.B1(n_236),
.B2(n_232),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_836),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_837),
.B(n_573),
.Y(n_1074)
);

INVx11_ASAP7_75t_L g1075 ( 
.A(n_927),
.Y(n_1075)
);

AOI22x1_ASAP7_75t_L g1076 ( 
.A1(n_837),
.A2(n_400),
.B1(n_399),
.B2(n_416),
.Y(n_1076)
);

NOR2xp67_ASAP7_75t_L g1077 ( 
.A(n_894),
.B(n_901),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_842),
.B(n_576),
.Y(n_1078)
);

NAND2x1_ASAP7_75t_L g1079 ( 
.A(n_913),
.B(n_797),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_829),
.B(n_299),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_842),
.A2(n_874),
.B(n_858),
.C(n_864),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_858),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_779),
.A2(n_818),
.B(n_813),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_864),
.B(n_576),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_874),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_L g1086 ( 
.A1(n_901),
.A2(n_226),
.B(n_218),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_781),
.A2(n_576),
.B(n_588),
.C(n_608),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_811),
.A2(n_588),
.B(n_608),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_797),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_883),
.B(n_784),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_895),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_903),
.A2(n_788),
.B(n_790),
.C(n_815),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_883),
.B(n_588),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_895),
.A2(n_751),
.B1(n_712),
.B2(n_543),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_913),
.A2(n_708),
.B(n_630),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_813),
.A2(n_708),
.B(n_630),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_828),
.A2(n_597),
.B(n_532),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_875),
.B(n_301),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_895),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_914),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_918),
.A2(n_776),
.B1(n_898),
.B2(n_797),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_918),
.A2(n_751),
.B1(n_712),
.B2(n_543),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_SL g1103 ( 
.A1(n_833),
.A2(n_531),
.B(n_547),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_934),
.A2(n_597),
.B(n_530),
.C(n_531),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_797),
.B(n_918),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_787),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_834),
.B(n_266),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_835),
.B(n_534),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_838),
.B(n_302),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_841),
.B(n_534),
.Y(n_1110)
);

AND2x6_ASAP7_75t_SL g1111 ( 
.A(n_855),
.B(n_543),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_923),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_848),
.A2(n_751),
.B(n_712),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_856),
.B(n_549),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_923),
.B(n_549),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_916),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1077),
.B(n_951),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1069),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_965),
.B(n_921),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1045),
.B(n_776),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_964),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1051),
.B(n_1053),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_961),
.A2(n_898),
.B(n_930),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_967),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_L g1125 ( 
.A(n_1031),
.B(n_818),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1045),
.B(n_931),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_957),
.A2(n_908),
.B(n_910),
.C(n_919),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1053),
.B(n_931),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_949),
.B(n_922),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_995),
.A2(n_910),
.B1(n_908),
.B2(n_933),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1099),
.B(n_932),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_995),
.A2(n_932),
.B1(n_919),
.B2(n_897),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1112),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_955),
.A2(n_610),
.B(n_630),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_938),
.B(n_1056),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1101),
.A2(n_376),
.B1(n_388),
.B2(n_399),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1097),
.A2(n_935),
.B(n_1005),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1112),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1092),
.A2(n_799),
.B(n_789),
.C(n_549),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_968),
.A2(n_530),
.B(n_708),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_978),
.B(n_549),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1069),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_967),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_978),
.B(n_549),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1068),
.A2(n_357),
.B1(n_315),
.B2(n_366),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_SL g1146 ( 
.A(n_1007),
.B(n_411),
.C(n_245),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_970),
.A2(n_975),
.B(n_953),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_L g1148 ( 
.A1(n_944),
.A2(n_555),
.B(n_551),
.C(n_610),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1092),
.A2(n_551),
.B(n_555),
.C(n_370),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1090),
.B(n_551),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1007),
.A2(n_751),
.B1(n_712),
.B2(n_266),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_945),
.B(n_551),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_957),
.A2(n_555),
.B(n_610),
.C(n_712),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_947),
.B(n_555),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_974),
.B(n_297),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1064),
.B(n_363),
.Y(n_1156)
);

INVxp33_ASAP7_75t_L g1157 ( 
.A(n_936),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_964),
.B(n_306),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1031),
.B(n_610),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_982),
.B(n_363),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_971),
.B(n_366),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_941),
.A2(n_297),
.B(n_376),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_1069),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1105),
.A2(n_370),
.B1(n_388),
.B2(n_389),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_999),
.B(n_389),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_R g1166 ( 
.A(n_943),
.B(n_400),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_L g1167 ( 
.A(n_1020),
.B(n_418),
.C(n_359),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1069),
.Y(n_1168)
);

OAI22x1_ASAP7_75t_L g1169 ( 
.A1(n_1058),
.A2(n_218),
.B1(n_217),
.B2(n_220),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_971),
.B(n_406),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_940),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1071),
.A2(n_406),
.B1(n_712),
.B2(n_751),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1006),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1109),
.B(n_751),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1109),
.B(n_309),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1089),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_974),
.B(n_297),
.Y(n_1177)
);

AND2x2_ASAP7_75t_SL g1178 ( 
.A(n_1098),
.B(n_297),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_942),
.A2(n_297),
.B(n_656),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_950),
.A2(n_656),
.B(n_313),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_989),
.B(n_319),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_979),
.A2(n_656),
.B(n_323),
.Y(n_1182)
);

NAND2x1_ASAP7_75t_L g1183 ( 
.A(n_1059),
.B(n_656),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_936),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1075),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_123),
.B(n_206),
.Y(n_1186)
);

NOR3xp33_ASAP7_75t_L g1187 ( 
.A(n_1098),
.B(n_969),
.C(n_1086),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_962),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1032),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1108),
.A2(n_328),
.B(n_347),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1089),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_989),
.B(n_962),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1110),
.A2(n_414),
.B(n_405),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1033),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1091),
.B(n_220),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1026),
.A2(n_93),
.B(n_203),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1024),
.B(n_76),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_994),
.A2(n_402),
.B1(n_401),
.B2(n_392),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_SL g1199 ( 
.A1(n_1107),
.A2(n_402),
.B(n_401),
.C(n_392),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1039),
.B(n_969),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1114),
.A2(n_387),
.B(n_382),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1011),
.A2(n_387),
.B(n_382),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1054),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1024),
.B(n_189),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1029),
.B(n_381),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_956),
.A2(n_381),
.B1(n_377),
.B2(n_368),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_998),
.A2(n_377),
.B(n_368),
.C(n_364),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1030),
.A2(n_364),
.B(n_362),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_948),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1058),
.B(n_362),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1025),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1089),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1001),
.A2(n_946),
.B1(n_1082),
.B2(n_1085),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1089),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_954),
.B(n_361),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1035),
.B(n_361),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1080),
.B(n_236),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_998),
.B(n_235),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_SL g1219 ( 
.A(n_996),
.B(n_232),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_976),
.B(n_186),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_1106),
.B(n_226),
.C(n_15),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_SL g1222 ( 
.A(n_1080),
.B(n_13),
.C(n_17),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1043),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_952),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1012),
.B(n_1038),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1044),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1052),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_976),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1072),
.B(n_19),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1073),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_976),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_959),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1055),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_992),
.B(n_179),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1043),
.B(n_140),
.Y(n_1235)
);

INVx5_ASAP7_75t_L g1236 ( 
.A(n_1059),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1081),
.A2(n_26),
.B(n_30),
.C(n_33),
.Y(n_1237)
);

AND2x4_ASAP7_75t_SL g1238 ( 
.A(n_1013),
.B(n_178),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_980),
.A2(n_175),
.B(n_170),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1072),
.B(n_1066),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1055),
.B(n_165),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1100),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1076),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1103),
.A2(n_36),
.B(n_41),
.C(n_46),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1013),
.Y(n_1245)
);

O2A1O1Ixp5_ASAP7_75t_L g1246 ( 
.A1(n_1014),
.A2(n_152),
.B(n_151),
.C(n_145),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_973),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1116),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1048),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1061),
.B(n_144),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1093),
.B(n_48),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1046),
.B(n_48),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1050),
.A2(n_118),
.B(n_130),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_972),
.B(n_52),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1065),
.B(n_52),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1079),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_986),
.B(n_135),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1023),
.A2(n_126),
.B(n_100),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_1111),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1088),
.A2(n_937),
.B(n_939),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1026),
.A2(n_127),
.B(n_99),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1041),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_972),
.B(n_53),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1070),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_958),
.A2(n_91),
.B(n_57),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_984),
.B(n_55),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_SL g1267 ( 
.A(n_1040),
.B(n_58),
.C(n_59),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1074),
.Y(n_1268)
);

OAI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_984),
.A2(n_61),
.B(n_62),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1049),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_960),
.A2(n_61),
.B(n_63),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1002),
.A2(n_63),
.B(n_64),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1037),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1083),
.B(n_65),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1018),
.A2(n_66),
.B(n_67),
.C(n_69),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1078),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1185),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1122),
.B(n_1018),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1189),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1217),
.A2(n_1009),
.B(n_1087),
.C(n_990),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1148),
.A2(n_966),
.B(n_1107),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1260),
.A2(n_1015),
.A3(n_985),
.B(n_993),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1134),
.A2(n_966),
.B(n_988),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1178),
.A2(n_977),
.B(n_983),
.C(n_1104),
.Y(n_1284)
);

AOI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1260),
.A2(n_1084),
.B(n_1057),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1228),
.B(n_1057),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1157),
.B(n_1027),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1117),
.A2(n_1115),
.B(n_1010),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1194),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1128),
.A2(n_1022),
.B(n_1017),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1149),
.A2(n_997),
.A3(n_987),
.B(n_991),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1240),
.A2(n_1060),
.B1(n_1028),
.B2(n_1034),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1137),
.A2(n_1004),
.B(n_1003),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1187),
.A2(n_1102),
.B(n_1094),
.C(n_1113),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1229),
.A2(n_1067),
.B(n_1008),
.C(n_1042),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1175),
.A2(n_1000),
.B(n_1021),
.C(n_1016),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1129),
.A2(n_981),
.B(n_1063),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1215),
.B(n_1041),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1242),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1252),
.B(n_1067),
.C(n_1008),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1247),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1199),
.A2(n_1036),
.B(n_1096),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1228),
.B(n_1047),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1257),
.A2(n_1095),
.B(n_1062),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1118),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1255),
.A2(n_1146),
.B1(n_1222),
.B2(n_1200),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1248),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1184),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_L g1309 ( 
.A(n_1124),
.Y(n_1309)
);

NAND3x1_ASAP7_75t_L g1310 ( 
.A(n_1221),
.B(n_1192),
.C(n_1210),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1167),
.A2(n_73),
.B(n_1153),
.C(n_1207),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1228),
.B(n_1235),
.Y(n_1312)
);

AO22x2_ASAP7_75t_L g1313 ( 
.A1(n_1222),
.A2(n_1146),
.B1(n_1213),
.B2(n_1202),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1143),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1147),
.A2(n_1123),
.B(n_1139),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1118),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1121),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1173),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1270),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1211),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1123),
.A2(n_1261),
.B(n_1196),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1244),
.A2(n_1161),
.B(n_1170),
.C(n_1216),
.Y(n_1322)
);

AOI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1158),
.A2(n_1181),
.B(n_1207),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1147),
.A2(n_1174),
.B(n_1141),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1120),
.A2(n_1126),
.B1(n_1233),
.B2(n_1144),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1241),
.A2(n_1250),
.B(n_1234),
.C(n_1263),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1203),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1119),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1188),
.B(n_1205),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1218),
.A2(n_1251),
.B(n_1274),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1132),
.A2(n_1236),
.B(n_1150),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1236),
.B(n_1212),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1224),
.A2(n_1267),
.B(n_1237),
.C(n_1195),
.Y(n_1333)
);

NOR2xp67_ASAP7_75t_SL g1334 ( 
.A(n_1236),
.B(n_1212),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1135),
.B(n_1259),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1226),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1230),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1166),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1220),
.A2(n_1231),
.B1(n_1257),
.B2(n_1136),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1145),
.B(n_1159),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1224),
.A2(n_1237),
.B(n_1275),
.C(n_1156),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1179),
.A2(n_1140),
.B(n_1186),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1190),
.B(n_1243),
.C(n_1201),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1130),
.A2(n_1180),
.B(n_1253),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1190),
.B(n_1201),
.C(n_1193),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1160),
.B(n_1165),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1148),
.A2(n_1271),
.B(n_1265),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_SL g1348 ( 
.A(n_1220),
.B(n_1219),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1227),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1180),
.A2(n_1253),
.B(n_1140),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1153),
.A2(n_1276),
.B(n_1264),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1232),
.A2(n_1249),
.B1(n_1214),
.B2(n_1212),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1162),
.A2(n_1127),
.B(n_1254),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_SL g1354 ( 
.A1(n_1266),
.A2(n_1269),
.B(n_1225),
.C(n_1268),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_SL g1355 ( 
.A1(n_1131),
.A2(n_1127),
.B(n_1239),
.C(n_1258),
.Y(n_1355)
);

AOI222xp33_ASAP7_75t_L g1356 ( 
.A1(n_1169),
.A2(n_1223),
.B1(n_1206),
.B2(n_1198),
.C1(n_1164),
.C2(n_1235),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1171),
.Y(n_1357)
);

AOI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1179),
.A2(n_1162),
.B(n_1182),
.Y(n_1358)
);

OAI22x1_ASAP7_75t_L g1359 ( 
.A1(n_1273),
.A2(n_1245),
.B1(n_1204),
.B2(n_1197),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1159),
.B(n_1133),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1193),
.A2(n_1208),
.B(n_1202),
.C(n_1246),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1208),
.B(n_1209),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1182),
.A2(n_1239),
.B(n_1214),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1272),
.A2(n_1258),
.A3(n_1154),
.B(n_1152),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1125),
.A2(n_1138),
.B1(n_1151),
.B2(n_1262),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1214),
.A2(n_1256),
.B(n_1183),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1262),
.B(n_1238),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1272),
.A2(n_1204),
.B(n_1197),
.C(n_1155),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1176),
.B(n_1118),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1172),
.A2(n_1256),
.B(n_1191),
.C(n_1177),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1191),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1142),
.A2(n_1163),
.B(n_1168),
.C(n_1191),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1168),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1178),
.A2(n_778),
.B1(n_902),
.B2(n_1217),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1121),
.B(n_965),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1189),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1097),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1228),
.B(n_1031),
.Y(n_1378)
);

CKINVDCx11_ASAP7_75t_R g1379 ( 
.A(n_1124),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1122),
.B(n_965),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1228),
.B(n_1031),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1217),
.A2(n_902),
.B(n_1053),
.C(n_616),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1122),
.B(n_778),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1217),
.A2(n_902),
.B(n_1053),
.C(n_616),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1217),
.A2(n_902),
.B(n_1053),
.C(n_616),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1260),
.A2(n_961),
.B(n_963),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1228),
.B(n_1031),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1260),
.A2(n_1147),
.B(n_1137),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1097),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1097),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1118),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1097),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1210),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1217),
.A2(n_778),
.B(n_951),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1217),
.A2(n_1053),
.B(n_616),
.C(n_951),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1122),
.B(n_951),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_SL g1397 ( 
.A1(n_1244),
.A2(n_957),
.B(n_951),
.C(n_778),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1122),
.B(n_778),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_SL g1399 ( 
.A1(n_1244),
.A2(n_957),
.B(n_951),
.C(n_778),
.Y(n_1399)
);

AOI221x1_ASAP7_75t_L g1400 ( 
.A1(n_1222),
.A2(n_902),
.B1(n_1007),
.B2(n_1187),
.C(n_1146),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1122),
.B(n_778),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1236),
.B(n_1212),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1121),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1097),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1217),
.A2(n_778),
.B(n_951),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1260),
.A2(n_961),
.B(n_963),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1122),
.B(n_778),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1236),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1097),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1217),
.A2(n_778),
.B(n_1077),
.C(n_1178),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1189),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1122),
.B(n_951),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1122),
.B(n_951),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1184),
.Y(n_1414)
);

AOI221x1_ASAP7_75t_L g1415 ( 
.A1(n_1222),
.A2(n_902),
.B1(n_1007),
.B2(n_1187),
.C(n_1146),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1260),
.A2(n_961),
.B(n_963),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1122),
.B(n_778),
.Y(n_1417)
);

AO32x2_ASAP7_75t_L g1418 ( 
.A1(n_1213),
.A2(n_826),
.A3(n_1130),
.B1(n_1132),
.B2(n_946),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1120),
.A2(n_1175),
.B(n_951),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1178),
.A2(n_778),
.B1(n_902),
.B2(n_1217),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1122),
.B(n_778),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1122),
.B(n_778),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1118),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1122),
.B(n_951),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1185),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1260),
.A2(n_961),
.B(n_963),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1148),
.A2(n_1260),
.B(n_1147),
.Y(n_1427)
);

AND2x6_ASAP7_75t_L g1428 ( 
.A(n_1220),
.B(n_1257),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1118),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1122),
.B(n_951),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1121),
.B(n_965),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1414),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1396),
.B(n_1412),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1308),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1391),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1374),
.A2(n_1420),
.B1(n_1398),
.B2(n_1407),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1391),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1374),
.A2(n_1420),
.B1(n_1421),
.B2(n_1306),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1379),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1383),
.A2(n_1422),
.B1(n_1417),
.B2(n_1401),
.Y(n_1440)
);

BUFx8_ASAP7_75t_L g1441 ( 
.A(n_1327),
.Y(n_1441)
);

BUFx12f_ASAP7_75t_L g1442 ( 
.A(n_1320),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1394),
.A2(n_1405),
.B1(n_1323),
.B2(n_1306),
.Y(n_1443)
);

BUFx8_ASAP7_75t_SL g1444 ( 
.A(n_1301),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1425),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1411),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1356),
.A2(n_1424),
.B1(n_1413),
.B2(n_1430),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1328),
.B(n_1380),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1313),
.A2(n_1343),
.B1(n_1339),
.B2(n_1346),
.Y(n_1449)
);

CKINVDCx14_ASAP7_75t_R g1450 ( 
.A(n_1309),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1279),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1313),
.A2(n_1343),
.B1(n_1348),
.B2(n_1278),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1428),
.A2(n_1345),
.B1(n_1353),
.B2(n_1325),
.Y(n_1453)
);

BUFx4_ASAP7_75t_R g1454 ( 
.A(n_1393),
.Y(n_1454)
);

BUFx12f_ASAP7_75t_L g1455 ( 
.A(n_1277),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1376),
.Y(n_1456)
);

NAND2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1334),
.B(n_1402),
.Y(n_1457)
);

INVx6_ASAP7_75t_L g1458 ( 
.A(n_1378),
.Y(n_1458)
);

CKINVDCx11_ASAP7_75t_R g1459 ( 
.A(n_1314),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1336),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1428),
.A2(n_1345),
.B1(n_1329),
.B2(n_1340),
.Y(n_1461)
);

BUFx4f_ASAP7_75t_SL g1462 ( 
.A(n_1381),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1319),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1428),
.A2(n_1393),
.B1(n_1382),
.B2(n_1384),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_1338),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1337),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1410),
.A2(n_1385),
.B1(n_1310),
.B2(n_1431),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1428),
.A2(n_1300),
.B1(n_1362),
.B2(n_1344),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1300),
.A2(n_1287),
.B1(n_1307),
.B2(n_1299),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1349),
.A2(n_1357),
.B1(n_1395),
.B2(n_1318),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1375),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1351),
.A2(n_1288),
.B1(n_1298),
.B2(n_1312),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1381),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1387),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1371),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1285),
.Y(n_1476)
);

CKINVDCx11_ASAP7_75t_R g1477 ( 
.A(n_1312),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1309),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1286),
.A2(n_1359),
.B1(n_1400),
.B2(n_1415),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1403),
.A2(n_1317),
.B1(n_1365),
.B2(n_1361),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1360),
.B(n_1286),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1369),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1367),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1305),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1335),
.A2(n_1399),
.B1(n_1397),
.B2(n_1326),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1322),
.B(n_1333),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1290),
.A2(n_1315),
.B1(n_1427),
.B2(n_1303),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1373),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1352),
.A2(n_1303),
.B1(n_1350),
.B2(n_1363),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1316),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1429),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1388),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1388),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1370),
.A2(n_1294),
.B(n_1368),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1292),
.A2(n_1408),
.B1(n_1331),
.B2(n_1332),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1408),
.A2(n_1311),
.B1(n_1427),
.B2(n_1341),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1297),
.A2(n_1292),
.B1(n_1324),
.B2(n_1426),
.Y(n_1497)
);

BUFx2_ASAP7_75t_R g1498 ( 
.A(n_1330),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1284),
.A2(n_1280),
.B(n_1416),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1302),
.A2(n_1347),
.B1(n_1281),
.B2(n_1418),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1354),
.B(n_1423),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1423),
.A2(n_1342),
.B1(n_1355),
.B2(n_1419),
.Y(n_1502)
);

BUFx8_ASAP7_75t_L g1503 ( 
.A(n_1372),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1295),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1366),
.A2(n_1321),
.B1(n_1293),
.B2(n_1304),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1296),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1364),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1283),
.A2(n_1389),
.B1(n_1404),
.B2(n_1392),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1364),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1291),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1358),
.A2(n_1282),
.B1(n_1291),
.B2(n_1377),
.Y(n_1511)
);

BUFx10_ASAP7_75t_L g1512 ( 
.A(n_1291),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1390),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1409),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1379),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1380),
.B(n_1383),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1334),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1374),
.A2(n_778),
.B1(n_1420),
.B2(n_1398),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1379),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1379),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1386),
.A2(n_1416),
.B(n_1406),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1289),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1383),
.A2(n_1178),
.B1(n_1401),
.B2(n_1398),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1383),
.A2(n_1178),
.B1(n_1401),
.B2(n_1398),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1289),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1289),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1383),
.A2(n_1178),
.B1(n_1401),
.B2(n_1398),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1379),
.Y(n_1530)
);

BUFx8_ASAP7_75t_SL g1531 ( 
.A(n_1301),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1308),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1383),
.A2(n_1178),
.B1(n_1401),
.B2(n_1398),
.Y(n_1537)
);

BUFx4f_ASAP7_75t_L g1538 ( 
.A(n_1428),
.Y(n_1538)
);

CKINVDCx11_ASAP7_75t_R g1539 ( 
.A(n_1379),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_SL g1540 ( 
.A(n_1425),
.Y(n_1540)
);

BUFx8_ASAP7_75t_SL g1541 ( 
.A(n_1301),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1383),
.A2(n_778),
.B1(n_1401),
.B2(n_1398),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1386),
.A2(n_1416),
.B(n_1406),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1374),
.A2(n_778),
.B1(n_1178),
.B2(n_1420),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1289),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1374),
.A2(n_778),
.B1(n_1420),
.B2(n_1398),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1380),
.B(n_1383),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1308),
.Y(n_1549)
);

CKINVDCx16_ASAP7_75t_R g1550 ( 
.A(n_1301),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1374),
.A2(n_778),
.B1(n_1420),
.B2(n_1398),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_SL g1552 ( 
.A(n_1308),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1308),
.Y(n_1553)
);

CKINVDCx6p67_ASAP7_75t_R g1554 ( 
.A(n_1379),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1289),
.Y(n_1555)
);

CKINVDCx11_ASAP7_75t_R g1556 ( 
.A(n_1379),
.Y(n_1556)
);

INVx8_ASAP7_75t_L g1557 ( 
.A(n_1391),
.Y(n_1557)
);

CKINVDCx6p67_ASAP7_75t_R g1558 ( 
.A(n_1379),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1308),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1383),
.A2(n_778),
.B1(n_1401),
.B2(n_1398),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1383),
.A2(n_1178),
.B1(n_1401),
.B2(n_1398),
.Y(n_1562)
);

BUFx12f_ASAP7_75t_L g1563 ( 
.A(n_1379),
.Y(n_1563)
);

BUFx4_ASAP7_75t_R g1564 ( 
.A(n_1393),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1391),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1383),
.A2(n_1401),
.B1(n_1407),
.B2(n_1398),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1514),
.B(n_1510),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1526),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1451),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1476),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1509),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1476),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1514),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1451),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1504),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1435),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1521),
.A2(n_1543),
.B(n_1511),
.Y(n_1577)
);

CKINVDCx11_ASAP7_75t_R g1578 ( 
.A(n_1439),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1443),
.A2(n_1524),
.B(n_1523),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1513),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1443),
.B(n_1452),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1507),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1452),
.B(n_1449),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1507),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1538),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1492),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1492),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1542),
.A2(n_1561),
.B1(n_1436),
.B2(n_1544),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1444),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1494),
.B(n_1499),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1486),
.B(n_1449),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1448),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1525),
.B(n_1526),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1432),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1512),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1493),
.A2(n_1497),
.B(n_1487),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1497),
.A2(n_1487),
.B(n_1468),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1512),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1495),
.A2(n_1546),
.B(n_1518),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1456),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1460),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1500),
.A2(n_1453),
.B(n_1468),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1506),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1538),
.B(n_1485),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1506),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1555),
.B(n_1516),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1506),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1466),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1547),
.B(n_1479),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1446),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1522),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1527),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1528),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1545),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1503),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1503),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1501),
.Y(n_1618)
);

OR2x6_ASAP7_75t_L g1619 ( 
.A(n_1480),
.B(n_1457),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1470),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1534),
.B(n_1536),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1470),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1500),
.A2(n_1453),
.B(n_1479),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1475),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1472),
.A2(n_1464),
.B(n_1461),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1502),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1488),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1471),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1481),
.B(n_1482),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1461),
.B(n_1548),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1496),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1469),
.B(n_1534),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1437),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1529),
.B(n_1562),
.C(n_1537),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1440),
.A2(n_1566),
.B1(n_1560),
.B2(n_1536),
.C(n_1447),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1472),
.A2(n_1464),
.B(n_1457),
.Y(n_1637)
);

BUFx4f_ASAP7_75t_L g1638 ( 
.A(n_1557),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1508),
.Y(n_1639)
);

BUFx4f_ASAP7_75t_SL g1640 ( 
.A(n_1563),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1467),
.B(n_1469),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1531),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1438),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1489),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1441),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1551),
.A2(n_1566),
.B1(n_1560),
.B2(n_1447),
.Y(n_1646)
);

CKINVDCx6p67_ASAP7_75t_R g1647 ( 
.A(n_1445),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1505),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1498),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1433),
.A2(n_1490),
.B(n_1491),
.Y(n_1650)
);

CKINVDCx10_ASAP7_75t_R g1651 ( 
.A(n_1550),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_1541),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1517),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1441),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1450),
.A2(n_1483),
.B1(n_1462),
.B2(n_1552),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1435),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1474),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1473),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_L g1659 ( 
.A(n_1579),
.B(n_1473),
.C(n_1477),
.Y(n_1659)
);

INVx5_ASAP7_75t_SL g1660 ( 
.A(n_1590),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1592),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1635),
.A2(n_1557),
.B(n_1450),
.C(n_1564),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1654),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1609),
.B(n_1458),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1636),
.B(n_1540),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1588),
.A2(n_1552),
.B1(n_1535),
.B2(n_1549),
.C(n_1434),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1646),
.A2(n_1559),
.B(n_1553),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1635),
.A2(n_1633),
.B1(n_1593),
.B2(n_1622),
.C(n_1621),
.Y(n_1668)
);

O2A1O1Ixp33_ASAP7_75t_SL g1669 ( 
.A1(n_1641),
.A2(n_1564),
.B(n_1454),
.C(n_1557),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1655),
.A2(n_1563),
.B1(n_1540),
.B2(n_1462),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1609),
.B(n_1484),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1609),
.Y(n_1672)
);

OAI211xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1643),
.A2(n_1478),
.B(n_1459),
.C(n_1445),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1641),
.A2(n_1568),
.B1(n_1603),
.B2(n_1590),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1582),
.B(n_1559),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1626),
.A2(n_1454),
.B(n_1565),
.C(n_1463),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1651),
.Y(n_1677)
);

BUFx8_ASAP7_75t_L g1678 ( 
.A(n_1654),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1619),
.B(n_1455),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1600),
.B(n_1465),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1590),
.A2(n_1599),
.B1(n_1633),
.B2(n_1631),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1600),
.B(n_1465),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1643),
.B(n_1558),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1569),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_SL g1686 ( 
.A1(n_1591),
.A2(n_1554),
.B(n_1556),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1650),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1631),
.B(n_1442),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1577),
.A2(n_1515),
.B(n_1519),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1601),
.B(n_1539),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1569),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1601),
.B(n_1520),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1607),
.B(n_1530),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_L g1694 ( 
.A(n_1637),
.B(n_1650),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1610),
.B(n_1602),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1573),
.B(n_1584),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1610),
.B(n_1602),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1573),
.B(n_1584),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1651),
.B(n_1594),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1602),
.B(n_1607),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1625),
.B(n_1611),
.Y(n_1701)
);

OR2x6_ASAP7_75t_L g1702 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1602),
.B(n_1624),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1653),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1589),
.B(n_1642),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1626),
.A2(n_1581),
.B(n_1637),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1573),
.B(n_1567),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_SL g1708 ( 
.A1(n_1591),
.A2(n_1575),
.B(n_1632),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_SL g1709 ( 
.A1(n_1649),
.A2(n_1632),
.B(n_1618),
.C(n_1644),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1624),
.B(n_1639),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1657),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1573),
.B(n_1567),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1624),
.B(n_1639),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1580),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1580),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1624),
.B(n_1574),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1649),
.A2(n_1605),
.B1(n_1608),
.B2(n_1606),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1599),
.A2(n_1644),
.B(n_1619),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1583),
.A2(n_1627),
.B(n_1648),
.C(n_1623),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1605),
.A2(n_1606),
.B1(n_1608),
.B2(n_1619),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1570),
.B(n_1572),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1654),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1597),
.A2(n_1653),
.B(n_1619),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_SL g1725 ( 
.A(n_1599),
.B(n_1598),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1570),
.B(n_1572),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1597),
.A2(n_1620),
.B(n_1648),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1652),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1630),
.B(n_1613),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1665),
.B(n_1647),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1661),
.B(n_1629),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1672),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1728),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1678),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.B(n_1695),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1674),
.A2(n_1605),
.B1(n_1604),
.B2(n_1620),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1707),
.B(n_1567),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1719),
.B(n_1585),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1672),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1714),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1700),
.B(n_1695),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1685),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1668),
.A2(n_1604),
.B1(n_1647),
.B2(n_1658),
.Y(n_1744)
);

AND2x4_ASAP7_75t_SL g1745 ( 
.A(n_1680),
.B(n_1567),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1697),
.B(n_1586),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1688),
.B(n_1645),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1697),
.B(n_1596),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1696),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1685),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1704),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1691),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1710),
.B(n_1713),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1713),
.B(n_1596),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1691),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1716),
.B(n_1598),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1679),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1716),
.B(n_1729),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1671),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1727),
.B(n_1618),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1706),
.B(n_1604),
.C(n_1628),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1722),
.Y(n_1762)
);

AOI222xp33_ASAP7_75t_L g1763 ( 
.A1(n_1659),
.A2(n_1640),
.B1(n_1578),
.B2(n_1613),
.C1(n_1614),
.C2(n_1615),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1721),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1687),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1701),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1664),
.B(n_1614),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1703),
.B(n_1587),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1707),
.B(n_1712),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1678),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1712),
.B(n_1595),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1703),
.B(n_1571),
.Y(n_1772)
);

INVx5_ASAP7_75t_L g1773 ( 
.A(n_1680),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1732),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1740),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1744),
.A2(n_1662),
.B1(n_1666),
.B2(n_1676),
.C(n_1688),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1741),
.B(n_1696),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1735),
.B(n_1694),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1735),
.B(n_1694),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1749),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1761),
.B(n_1724),
.C(n_1682),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1734),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1741),
.B(n_1711),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1772),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1738),
.A2(n_1662),
.B1(n_1676),
.B2(n_1680),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1763),
.A2(n_1702),
.B1(n_1680),
.B2(n_1684),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.B(n_1698),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1753),
.B(n_1698),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_SL g1789 ( 
.A(n_1760),
.B(n_1667),
.C(n_1717),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1739),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1731),
.A2(n_1718),
.B(n_1692),
.C(n_1693),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1767),
.B(n_1681),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1750),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1750),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1736),
.A2(n_1708),
.B1(n_1709),
.B2(n_1669),
.C(n_1681),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1758),
.B(n_1698),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1747),
.A2(n_1702),
.B1(n_1720),
.B2(n_1660),
.Y(n_1798)
);

OR2x6_ASAP7_75t_L g1799 ( 
.A(n_1734),
.B(n_1702),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1758),
.B(n_1690),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1733),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1773),
.B(n_1689),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1746),
.B(n_1768),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1740),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1769),
.B(n_1690),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1751),
.B(n_1683),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1768),
.B(n_1726),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1752),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1734),
.A2(n_1702),
.B1(n_1660),
.B2(n_1670),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1752),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1737),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1769),
.B(n_1725),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1771),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1759),
.B(n_1683),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1773),
.A2(n_1709),
.B(n_1669),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1755),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1770),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1742),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1756),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1775),
.B(n_1764),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1793),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1793),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1804),
.B(n_1764),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1790),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1818),
.B(n_1757),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1813),
.B(n_1748),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1784),
.B(n_1765),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1794),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1794),
.B(n_1766),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1808),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1811),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1790),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1780),
.B(n_1754),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1780),
.B(n_1754),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1808),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1802),
.B(n_1773),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1802),
.B(n_1773),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1802),
.B(n_1773),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1797),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1811),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1810),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1816),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1785),
.B(n_1677),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1811),
.B(n_1773),
.Y(n_1844)
);

INVx3_ASAP7_75t_SL g1845 ( 
.A(n_1817),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1791),
.B(n_1730),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1803),
.B(n_1762),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1812),
.B(n_1762),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1812),
.B(n_1762),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_1782),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1774),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1774),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1821),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1827),
.B(n_1803),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1827),
.B(n_1783),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1836),
.B(n_1777),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1824),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1836),
.B(n_1777),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1824),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1824),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1821),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1836),
.B(n_1787),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1822),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1822),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1828),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1836),
.B(n_1799),
.Y(n_1866)
);

OAI21xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1846),
.A2(n_1805),
.B(n_1800),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1828),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1836),
.B(n_1787),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1827),
.B(n_1783),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1850),
.B(n_1800),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1825),
.B(n_1778),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1778),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1788),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1837),
.B(n_1788),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1847),
.B(n_1779),
.Y(n_1876)
);

INVxp67_ASAP7_75t_SL g1877 ( 
.A(n_1850),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1850),
.B(n_1814),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1832),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1846),
.B(n_1814),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1830),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1845),
.B(n_1806),
.Y(n_1883)
);

NOR5xp2_ASAP7_75t_L g1884 ( 
.A(n_1845),
.B(n_1781),
.C(n_1776),
.D(n_1673),
.E(n_1819),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1845),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1830),
.Y(n_1887)
);

INVxp67_ASAP7_75t_SL g1888 ( 
.A(n_1829),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1837),
.B(n_1805),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1832),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1832),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1847),
.B(n_1779),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1835),
.Y(n_1893)
);

AOI32xp33_ASAP7_75t_L g1894 ( 
.A1(n_1843),
.A2(n_1786),
.A3(n_1795),
.B1(n_1809),
.B2(n_1817),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1847),
.B(n_1807),
.Y(n_1895)
);

NAND2x1_ASAP7_75t_L g1896 ( 
.A(n_1838),
.B(n_1799),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1835),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1845),
.B(n_1792),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1855),
.B(n_1820),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1853),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1877),
.B(n_1848),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1881),
.B(n_1848),
.Y(n_1902)
);

AND2x2_ASAP7_75t_SL g1903 ( 
.A(n_1884),
.B(n_1817),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1855),
.B(n_1820),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1889),
.B(n_1838),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1853),
.Y(n_1906)
);

NOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1886),
.B(n_1770),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1871),
.B(n_1677),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1878),
.B(n_1848),
.Y(n_1909)
);

AND2x4_ASAP7_75t_SL g1910 ( 
.A(n_1866),
.B(n_1799),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1867),
.A2(n_1843),
.B(n_1883),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1861),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1889),
.B(n_1838),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1870),
.B(n_1823),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1861),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1870),
.Y(n_1916)
);

INVxp67_ASAP7_75t_SL g1917 ( 
.A(n_1896),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1863),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1898),
.B(n_1849),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1856),
.B(n_1838),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1863),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1888),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1854),
.B(n_1823),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1857),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1866),
.B(n_1728),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1894),
.B(n_1849),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1856),
.B(n_1838),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1894),
.B(n_1849),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1857),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1854),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1864),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1866),
.B(n_1801),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1896),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1859),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1864),
.Y(n_1935)
);

NOR4xp25_ASAP7_75t_L g1936 ( 
.A(n_1926),
.B(n_1789),
.C(n_1865),
.D(n_1893),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1916),
.B(n_1858),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1935),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1903),
.A2(n_1686),
.B1(n_1782),
.B2(n_1885),
.Y(n_1940)
);

AOI222xp33_ASAP7_75t_L g1941 ( 
.A1(n_1903),
.A2(n_1880),
.B1(n_1869),
.B2(n_1862),
.C1(n_1858),
.C2(n_1874),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1925),
.B(n_1908),
.Y(n_1942)
);

OAI32xp33_ASAP7_75t_L g1943 ( 
.A1(n_1928),
.A2(n_1872),
.A3(n_1873),
.B1(n_1892),
.B2(n_1876),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1900),
.Y(n_1944)
);

OAI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1911),
.A2(n_1798),
.B1(n_1873),
.B2(n_1872),
.C(n_1815),
.Y(n_1945)
);

AOI322xp5_ASAP7_75t_L g1946 ( 
.A1(n_1903),
.A2(n_1862),
.A3(n_1885),
.B1(n_1880),
.B2(n_1875),
.C1(n_1874),
.C2(n_1869),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1920),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1900),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1907),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1916),
.B(n_1875),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1922),
.A2(n_1770),
.B1(n_1660),
.B2(n_1799),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1932),
.A2(n_1844),
.B1(n_1745),
.B2(n_1893),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1906),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1933),
.A2(n_1917),
.B1(n_1910),
.B2(n_1907),
.Y(n_1954)
);

AOI21xp33_ASAP7_75t_L g1955 ( 
.A1(n_1901),
.A2(n_1868),
.B(n_1865),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1906),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1902),
.B(n_1833),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1910),
.A2(n_1705),
.B(n_1699),
.Y(n_1958)
);

AOI21xp33_ASAP7_75t_L g1959 ( 
.A1(n_1899),
.A2(n_1882),
.B(n_1868),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1920),
.B(n_1678),
.Y(n_1960)
);

AOI211x1_ASAP7_75t_L g1961 ( 
.A1(n_1927),
.A2(n_1834),
.B(n_1833),
.C(n_1826),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1909),
.B(n_1895),
.Y(n_1962)
);

AOI21xp33_ASAP7_75t_SL g1963 ( 
.A1(n_1899),
.A2(n_1844),
.B(n_1895),
.Y(n_1963)
);

OAI322xp33_ASAP7_75t_L g1964 ( 
.A1(n_1904),
.A2(n_1876),
.A3(n_1892),
.B1(n_1897),
.B2(n_1882),
.C1(n_1887),
.C2(n_1891),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1936),
.B(n_1927),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1937),
.B(n_1919),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1944),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1948),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1941),
.A2(n_1913),
.B1(n_1905),
.B2(n_1844),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1953),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_SL g1971 ( 
.A1(n_1943),
.A2(n_1905),
.B1(n_1913),
.B2(n_1912),
.Y(n_1971)
);

A2O1A1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1946),
.A2(n_1617),
.B(n_1616),
.C(n_1689),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1942),
.A2(n_1915),
.B(n_1912),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1947),
.B(n_1940),
.Y(n_1974)
);

A2O1A1Ixp33_ASAP7_75t_SL g1975 ( 
.A1(n_1954),
.A2(n_1921),
.B(n_1918),
.C(n_1915),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1945),
.A2(n_1918),
.B1(n_1931),
.B2(n_1921),
.Y(n_1976)
);

NAND2x1_ASAP7_75t_L g1977 ( 
.A(n_1940),
.B(n_1931),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1939),
.Y(n_1978)
);

NAND3x2_ASAP7_75t_L g1979 ( 
.A(n_1962),
.B(n_1914),
.C(n_1904),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1949),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1956),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1950),
.B(n_1923),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1938),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1960),
.B(n_1914),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1964),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1951),
.B(n_1923),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1985),
.A2(n_1952),
.B1(n_1951),
.B2(n_1957),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1967),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1980),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1968),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1977),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1978),
.B(n_1958),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1978),
.A2(n_1975),
.B1(n_1965),
.B2(n_1973),
.C(n_1983),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1970),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1981),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1982),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1974),
.B(n_1963),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1984),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1971),
.A2(n_1969),
.B1(n_1976),
.B2(n_1986),
.Y(n_1999)
);

NAND3xp33_ASAP7_75t_L g2000 ( 
.A(n_1993),
.B(n_1975),
.C(n_1971),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1989),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1999),
.A2(n_1976),
.B(n_1972),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1998),
.B(n_1966),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1997),
.B(n_1961),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1991),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1992),
.B(n_1972),
.Y(n_2006)
);

NOR4xp75_ASAP7_75t_L g2007 ( 
.A(n_1995),
.B(n_1979),
.C(n_1955),
.D(n_1959),
.Y(n_2007)
);

OAI211xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1993),
.A2(n_1934),
.B(n_1929),
.C(n_1924),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1992),
.A2(n_1844),
.B1(n_1929),
.B2(n_1924),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1987),
.A2(n_1844),
.B1(n_1840),
.B2(n_1831),
.Y(n_2010)
);

OAI211xp5_ASAP7_75t_SL g2011 ( 
.A1(n_2002),
.A2(n_1996),
.B(n_1989),
.C(n_1990),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_2000),
.B(n_1995),
.C(n_1994),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_2006),
.A2(n_1988),
.B(n_1934),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2005),
.Y(n_2014)
);

NAND4xp25_ASAP7_75t_SL g2015 ( 
.A(n_2004),
.B(n_1897),
.C(n_1887),
.D(n_1890),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_2008),
.A2(n_1891),
.B1(n_1890),
.B2(n_1879),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2003),
.Y(n_2017)
);

XNOR2xp5_ASAP7_75t_L g2018 ( 
.A(n_2014),
.B(n_2007),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_2017),
.Y(n_2019)
);

OAI221xp5_ASAP7_75t_L g2020 ( 
.A1(n_2011),
.A2(n_2009),
.B1(n_2010),
.B2(n_2001),
.C(n_1663),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_2012),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2013),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_2015),
.A2(n_1723),
.B1(n_1663),
.B2(n_1675),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_2016),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_2014),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2025),
.Y(n_2026)
);

XNOR2xp5_ASAP7_75t_L g2027 ( 
.A(n_2018),
.B(n_1616),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2025),
.Y(n_2028)
);

NOR2x1_ASAP7_75t_L g2029 ( 
.A(n_2022),
.B(n_1616),
.Y(n_2029)
);

NAND4xp75_ASAP7_75t_L g2030 ( 
.A(n_2021),
.B(n_1879),
.C(n_1860),
.D(n_1859),
.Y(n_2030)
);

NOR2x1p5_ASAP7_75t_L g2031 ( 
.A(n_2020),
.B(n_1617),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2027),
.A2(n_2024),
.B(n_2019),
.C(n_2023),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2026),
.B(n_1860),
.Y(n_2033)
);

AOI22x1_ASAP7_75t_L g2034 ( 
.A1(n_2031),
.A2(n_1840),
.B1(n_1831),
.B2(n_1675),
.Y(n_2034)
);

O2A1O1Ixp33_ASAP7_75t_L g2035 ( 
.A1(n_2032),
.A2(n_2028),
.B(n_2033),
.C(n_2029),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2035),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2036),
.Y(n_2037)
);

AOI211xp5_ASAP7_75t_L g2038 ( 
.A1(n_2036),
.A2(n_2034),
.B(n_2030),
.C(n_1617),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_2037),
.A2(n_1840),
.B1(n_1831),
.B2(n_1723),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_2038),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_2040),
.A2(n_1675),
.B(n_1638),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2039),
.A2(n_1831),
.B1(n_1840),
.B2(n_1839),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_2041),
.A2(n_1638),
.B(n_1831),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_2043),
.A2(n_2042),
.B(n_1638),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_2044),
.A2(n_1840),
.B1(n_1834),
.B2(n_1833),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2045),
.A2(n_1852),
.B1(n_1851),
.B2(n_1841),
.C(n_1842),
.Y(n_2046)
);

AOI211xp5_ASAP7_75t_L g2047 ( 
.A1(n_2046),
.A2(n_1634),
.B(n_1656),
.C(n_1576),
.Y(n_2047)
);


endmodule