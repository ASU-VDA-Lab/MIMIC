module fake_jpeg_12419_n_94 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_12),
.B(n_27),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_31),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_58),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_39),
.B1(n_13),
.B2(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_11),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_68),
.B(n_9),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_6),
.B(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_R g75 ( 
.A(n_62),
.B(n_8),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.C(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_8),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_67),
.C(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_74),
.B1(n_72),
.B2(n_76),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_SL g88 ( 
.A1(n_86),
.A2(n_87),
.A3(n_75),
.B1(n_63),
.B2(n_85),
.C1(n_82),
.C2(n_84),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_74),
.B1(n_66),
.B2(n_73),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_15),
.B(n_18),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_19),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_20),
.B(n_23),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_25),
.B(n_29),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g94 ( 
.A(n_93),
.Y(n_94)
);


endmodule