module fake_ariane_1341_n_1665 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1665);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1665;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1468;
wire n_1253;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g159 ( 
.A(n_43),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_19),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_32),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_46),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_105),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_23),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_5),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_36),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_41),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_49),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_93),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_66),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

BUFx2_ASAP7_75t_SL g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_95),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_39),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_45),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_17),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_4),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_44),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_8),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_60),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_118),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_51),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_40),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_51),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_83),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_121),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_9),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_59),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_103),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_20),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_91),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_134),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_120),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_77),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_32),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_21),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_7),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_72),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_5),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_92),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_71),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_73),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_37),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_130),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_86),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_99),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_49),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_48),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_52),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_138),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_19),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_87),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_108),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_25),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_18),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_84),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_13),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_24),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_109),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_96),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_26),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_44),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_135),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_14),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_58),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_18),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_29),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_24),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_56),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_36),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_122),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_128),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_75),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_3),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_11),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_107),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_1),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_39),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_101),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_23),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_158),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_94),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_97),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_63),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_25),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_21),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_153),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_156),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_53),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_123),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_64),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_119),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_125),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_13),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_148),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_27),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_22),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_26),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_82),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_76),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_202),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_R g318 ( 
.A(n_172),
.B(n_79),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_177),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_274),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_197),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_197),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_179),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_209),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_291),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_209),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_236),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_171),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_231),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_203),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_200),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_207),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_191),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_231),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_208),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_212),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_218),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_191),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_216),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_200),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_218),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_222),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_284),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_226),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_237),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_226),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_240),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_248),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_163),
.B(n_0),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_257),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_255),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_263),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_309),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_264),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_257),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_173),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_181),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_185),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_187),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_235),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_164),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_189),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_211),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_247),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_252),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_256),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_258),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_259),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_260),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_265),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_272),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_267),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_220),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_271),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_165),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_280),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_278),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_165),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_285),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_327),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_342),
.B(n_166),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_339),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_342),
.B(n_160),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_326),
.B(n_182),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_228),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_228),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_345),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_346),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_351),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_350),
.B(n_323),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_334),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_354),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_357),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_R g426 ( 
.A(n_359),
.B(n_206),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_324),
.B(n_269),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_340),
.B(n_269),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_363),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_352),
.B(n_184),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_311),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_364),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_353),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_366),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_334),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_382),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_318),
.B(n_220),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_356),
.B(n_311),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_356),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_388),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_358),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_362),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_362),
.B(n_227),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_337),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_333),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_335),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_335),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_322),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_399),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_438),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_385),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_420),
.B(n_376),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_420),
.A2(n_319),
.B1(n_361),
.B2(n_227),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_426),
.B(n_160),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_420),
.A2(n_312),
.B1(n_297),
.B2(n_296),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_415),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_452),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_420),
.B(n_368),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_401),
.B(n_162),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_397),
.B(n_368),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_405),
.B(n_162),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_410),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_399),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_416),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_433),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_369),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_392),
.B(n_369),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_392),
.B(n_370),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_433),
.Y(n_492)
);

AO22x2_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_159),
.B1(n_294),
.B2(n_391),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_393),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_394),
.B(n_370),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_417),
.B(n_169),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_371),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_436),
.B(n_427),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_394),
.B(n_400),
.C(n_396),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_403),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_449),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_402),
.B(n_371),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_432),
.B(n_374),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_402),
.Y(n_512)
);

AND3x2_ASAP7_75t_L g513 ( 
.A(n_454),
.B(n_243),
.C(n_374),
.Y(n_513)
);

NOR3xp33_ASAP7_75t_L g514 ( 
.A(n_421),
.B(n_168),
.C(n_167),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_432),
.B(n_375),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_430),
.B(n_375),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_456),
.A2(n_280),
.B1(n_389),
.B2(n_386),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_456),
.A2(n_280),
.B1(n_389),
.B2(n_386),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_451),
.B(n_377),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_437),
.B(n_377),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_404),
.B(n_378),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_404),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_422),
.B(n_169),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_421),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_413),
.B(n_378),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_423),
.B(n_176),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_413),
.B(n_301),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_409),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_414),
.B(n_379),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_462),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_444),
.A2(n_298),
.B1(n_167),
.B2(n_170),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_452),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_418),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_449),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_379),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_437),
.B(n_380),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_409),
.B(n_380),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_437),
.B(n_447),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_456),
.A2(n_391),
.B1(n_384),
.B2(n_381),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_435),
.B(n_381),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_439),
.B(n_443),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_429),
.B(n_384),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_449),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_456),
.A2(n_224),
.B1(n_348),
.B2(n_347),
.Y(n_555)
);

OA22x2_ASAP7_75t_L g556 ( 
.A1(n_437),
.A2(n_338),
.B1(n_348),
.B2(n_347),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_445),
.B(n_192),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_431),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_409),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_409),
.B(n_176),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_412),
.B(n_178),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_412),
.B(n_178),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_R g565 ( 
.A(n_403),
.B(n_341),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_447),
.B(n_338),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_450),
.B(n_168),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_440),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_441),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_446),
.B(n_180),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_442),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_412),
.B(n_434),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_442),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_448),
.B(n_239),
.C(n_195),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_447),
.A2(n_412),
.B1(n_434),
.B2(n_463),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_434),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_447),
.B(n_180),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_L g583 ( 
.A1(n_444),
.A2(n_170),
.B1(n_174),
.B2(n_290),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_186),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_453),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_395),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_453),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_455),
.B(n_186),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_455),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_461),
.B(n_344),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_457),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_450),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_461),
.B(n_344),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_457),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_398),
.B(n_188),
.Y(n_597)
);

INVx4_ASAP7_75t_SL g598 ( 
.A(n_463),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_420),
.B(n_188),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_420),
.B(n_174),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_458),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_458),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_426),
.B(n_190),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_426),
.B(n_190),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_438),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_426),
.B(n_238),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_415),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_438),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_452),
.B(n_175),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_410),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_410),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_410),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_420),
.B(n_238),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_509),
.B(n_279),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_507),
.B(n_355),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_509),
.B(n_279),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_508),
.A2(n_213),
.B(n_276),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_500),
.B(n_283),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_475),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_467),
.B(n_283),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_506),
.B(n_175),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_547),
.B(n_286),
.Y(n_622)
);

AND2x6_ASAP7_75t_SL g623 ( 
.A(n_557),
.B(n_464),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_483),
.B(n_286),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_506),
.B(n_288),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_507),
.B(n_365),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_511),
.B(n_288),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_494),
.B(n_193),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_592),
.B(n_293),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_511),
.B(n_293),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_556),
.A2(n_183),
.B1(n_281),
.B2(n_290),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_494),
.B(n_193),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_468),
.B(n_194),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_516),
.A2(n_295),
.B1(n_314),
.B2(n_310),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_519),
.A2(n_295),
.B1(n_314),
.B2(n_310),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_489),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_475),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_499),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_302),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_515),
.B(n_302),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_531),
.A2(n_306),
.B1(n_307),
.B2(n_201),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_515),
.B(n_306),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_508),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_482),
.B(n_194),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_479),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_499),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_592),
.B(n_196),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_468),
.B(n_307),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_466),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_466),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_196),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_509),
.B(n_198),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_541),
.B(n_281),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_538),
.B(n_282),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_541),
.B(n_282),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_541),
.B(n_287),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_538),
.B(n_554),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_523),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_527),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_538),
.B(n_287),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_527),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_576),
.A2(n_246),
.B(n_204),
.C(n_205),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_554),
.B(n_292),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_554),
.B(n_292),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_470),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_537),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_576),
.B(n_298),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_303),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_489),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_531),
.B(n_303),
.Y(n_671)
);

AND2x6_ASAP7_75t_SL g672 ( 
.A(n_489),
.B(n_497),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_537),
.A2(n_199),
.B(n_254),
.C(n_261),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_470),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_560),
.B(n_305),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_560),
.B(n_305),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_605),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_479),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_589),
.B(n_308),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_589),
.A2(n_308),
.B1(n_219),
.B2(n_304),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_589),
.B(n_210),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_489),
.B(n_1),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_481),
.B(n_214),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_521),
.B(n_540),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_592),
.B(n_215),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_L g686 ( 
.A(n_592),
.B(n_581),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_552),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_556),
.A2(n_221),
.B1(n_229),
.B2(n_300),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_605),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_592),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_561),
.B(n_223),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_551),
.B(n_251),
.C(n_299),
.Y(n_692)
);

CKINVDCx11_ASAP7_75t_R g693 ( 
.A(n_487),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_608),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_497),
.B(n_6),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_487),
.B(n_217),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_520),
.B(n_225),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_520),
.B(n_230),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_595),
.B(n_301),
.Y(n_699)
);

OAI221xp5_ASAP7_75t_L g700 ( 
.A1(n_469),
.A2(n_270),
.B1(n_273),
.B2(n_250),
.C(n_277),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_552),
.A2(n_6),
.B(n_9),
.C(n_10),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_472),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_520),
.B(n_315),
.Y(n_703)
);

AND2x6_ASAP7_75t_SL g704 ( 
.A(n_497),
.B(n_10),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_608),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_497),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_586),
.B(n_244),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_540),
.B(n_245),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_505),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_562),
.B(n_12),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_544),
.B(n_242),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_253),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_505),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_502),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_599),
.B(n_268),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_580),
.A2(n_266),
.B1(n_262),
.B2(n_241),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_613),
.B(n_301),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_602),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_563),
.B(n_14),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_595),
.B(n_543),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_R g722 ( 
.A(n_526),
.B(n_62),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_567),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_572),
.B(n_574),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_595),
.B(n_301),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_577),
.A2(n_301),
.B1(n_275),
.B2(n_27),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_572),
.B(n_301),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_574),
.B(n_301),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_595),
.B(n_275),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_484),
.B(n_15),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_536),
.A2(n_275),
.B1(n_16),
.B2(n_28),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_556),
.A2(n_275),
.B1(n_28),
.B2(n_29),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_564),
.B(n_15),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_587),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_496),
.B(n_30),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_587),
.B(n_30),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_536),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_594),
.B(n_31),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_609),
.B(n_275),
.C(n_37),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_594),
.B(n_34),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_596),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_526),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_609),
.B(n_34),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_586),
.B(n_38),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_472),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_596),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_568),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_473),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_476),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_493),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_586),
.B(n_47),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_568),
.B(n_490),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_476),
.Y(n_753)
);

BUFx6f_ASAP7_75t_SL g754 ( 
.A(n_565),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_512),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_512),
.Y(n_756)
);

OR2x6_ASAP7_75t_L g757 ( 
.A(n_581),
.B(n_50),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_524),
.B(n_50),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_535),
.B(n_52),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_491),
.B(n_57),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_600),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_478),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_525),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_525),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_495),
.B(n_68),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_602),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_532),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_583),
.B(n_69),
.C(n_70),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_595),
.B(n_74),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_510),
.B(n_78),
.Y(n_770)
);

O2A1O1Ixp5_ASAP7_75t_L g771 ( 
.A1(n_532),
.A2(n_85),
.B(n_89),
.C(n_100),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_600),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_522),
.B(n_104),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_493),
.A2(n_106),
.B1(n_117),
.B2(n_126),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_542),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_542),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_543),
.B(n_133),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_514),
.B(n_140),
.C(n_144),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_678),
.B(n_601),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_724),
.A2(n_502),
.B(n_558),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_615),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_752),
.B(n_546),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_637),
.B(n_564),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_719),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_620),
.B(n_618),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_670),
.B(n_598),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_725),
.A2(n_548),
.B(n_559),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_737),
.B(n_571),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_730),
.A2(n_573),
.B(n_591),
.C(n_578),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_622),
.B(n_555),
.Y(n_790)
);

INVx11_ASAP7_75t_L g791 ( 
.A(n_693),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_623),
.B(n_529),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_650),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_679),
.B(n_533),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_730),
.A2(n_591),
.B(n_585),
.C(n_578),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_727),
.A2(n_611),
.B(n_485),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_759),
.A2(n_597),
.B(n_584),
.C(n_588),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_679),
.B(n_539),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_658),
.A2(n_478),
.B(n_492),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_658),
.A2(n_492),
.B(n_488),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_766),
.B(n_579),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_626),
.B(n_493),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_706),
.A2(n_606),
.B1(n_604),
.B2(n_471),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_690),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_725),
.A2(n_607),
.B(n_504),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_653),
.A2(n_607),
.B(n_488),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_690),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_702),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_653),
.A2(n_616),
.B(n_614),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_733),
.B(n_684),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_733),
.B(n_582),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_614),
.A2(n_504),
.B(n_530),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_644),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_616),
.A2(n_530),
.B(n_465),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_709),
.A2(n_585),
.B(n_573),
.Y(n_815)
);

INVx8_ASAP7_75t_L g816 ( 
.A(n_742),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_735),
.A2(n_553),
.B(n_528),
.C(n_579),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_772),
.A2(n_603),
.B1(n_575),
.B2(n_517),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_735),
.B(n_590),
.C(n_593),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_742),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_728),
.A2(n_765),
.B(n_760),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_646),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_758),
.A2(n_534),
.B(n_549),
.C(n_590),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_772),
.A2(n_518),
.B1(n_549),
.B2(n_534),
.Y(n_824)
);

BUFx2_ASAP7_75t_SL g825 ( 
.A(n_754),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_624),
.B(n_593),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_704),
.Y(n_827)
);

OAI321xp33_ASAP7_75t_L g828 ( 
.A1(n_750),
.A2(n_474),
.A3(n_570),
.B1(n_569),
.B2(n_493),
.C(n_465),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_650),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_655),
.B(n_569),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_629),
.B(n_543),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_742),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_772),
.A2(n_534),
.B1(n_549),
.B2(n_501),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_721),
.A2(n_611),
.B(n_485),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_655),
.B(n_661),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_633),
.B(n_513),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_661),
.B(n_570),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_659),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_645),
.B(n_503),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_709),
.A2(n_611),
.B(n_480),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_634),
.B(n_486),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_660),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_627),
.B(n_486),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_770),
.A2(n_480),
.B(n_485),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_758),
.B(n_503),
.C(n_501),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_773),
.A2(n_480),
.B(n_501),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_681),
.A2(n_503),
.B(n_477),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_648),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_651),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_718),
.A2(n_477),
.B(n_498),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_664),
.A2(n_498),
.B(n_612),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_645),
.B(n_477),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_635),
.B(n_612),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_731),
.A2(n_598),
.B(n_545),
.C(n_566),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_631),
.B(n_598),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_702),
.Y(n_856)
);

BUFx4f_ASAP7_75t_L g857 ( 
.A(n_757),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_665),
.A2(n_612),
.B(n_610),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_636),
.B(n_612),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_641),
.B(n_643),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_714),
.A2(n_610),
.B(n_545),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_649),
.B(n_566),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_662),
.A2(n_610),
.B(n_566),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_729),
.A2(n_610),
.B(n_545),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_744),
.B(n_545),
.C(n_566),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_621),
.B(n_691),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_648),
.B(n_632),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_667),
.A2(n_566),
.B(n_545),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_682),
.A2(n_145),
.B1(n_695),
.B2(n_711),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_711),
.A2(n_720),
.B(n_691),
.C(n_734),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_672),
.B(n_743),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_686),
.B(n_696),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_720),
.A2(n_741),
.B(n_710),
.C(n_687),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_632),
.B(n_628),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_723),
.A2(n_746),
.B(n_753),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_748),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_666),
.Y(n_877)
);

CKINVDCx10_ASAP7_75t_R g878 ( 
.A(n_754),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_708),
.B(n_668),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_722),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_714),
.A2(n_756),
.B(n_776),
.Y(n_881)
);

AOI21xp33_ASAP7_75t_L g882 ( 
.A1(n_700),
.A2(n_712),
.B(n_713),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_625),
.B(n_652),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_669),
.B(n_688),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_680),
.A2(n_656),
.B(n_657),
.C(n_654),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_755),
.A2(n_763),
.B(n_756),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_717),
.B(n_716),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_736),
.A2(n_740),
.B(n_738),
.C(n_671),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_688),
.B(n_683),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_757),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_739),
.A2(n_732),
.B(n_726),
.C(n_761),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_755),
.A2(n_776),
.B(n_763),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_749),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_764),
.A2(n_775),
.B(n_767),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_762),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_775),
.A2(n_777),
.B(n_630),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_777),
.A2(n_675),
.B(n_676),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_685),
.A2(n_689),
.B(n_677),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_732),
.A2(n_747),
.B1(n_774),
.B2(n_745),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_642),
.B(n_647),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_757),
.B(n_750),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_666),
.A2(n_674),
.B(n_705),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_751),
.B(n_697),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_701),
.A2(n_663),
.B(n_715),
.C(n_673),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_674),
.A2(n_677),
.B(n_694),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_698),
.B(n_707),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_689),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_694),
.A2(n_705),
.B(n_619),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_703),
.B(n_774),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_638),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_638),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_640),
.B(n_692),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_699),
.A2(n_769),
.B(n_639),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_768),
.B(n_778),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_617),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_769),
.A2(n_639),
.B(n_771),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_730),
.A2(n_758),
.B(n_735),
.C(n_720),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_711),
.A2(n_720),
.B(n_616),
.C(n_614),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_637),
.B(n_507),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_620),
.A2(n_759),
.B(n_731),
.C(n_622),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_752),
.B(n_500),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_644),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_658),
.A2(n_724),
.B(n_653),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_724),
.A2(n_658),
.B(n_653),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_724),
.A2(n_658),
.B(n_653),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_658),
.A2(n_724),
.B(n_653),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_724),
.A2(n_620),
.B1(n_658),
.B2(n_644),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_724),
.A2(n_658),
.B(n_653),
.Y(n_928)
);

AOI21x1_ASAP7_75t_L g929 ( 
.A1(n_721),
.A2(n_725),
.B(n_760),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_678),
.B(n_321),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_615),
.B(n_507),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_724),
.A2(n_620),
.B1(n_658),
.B2(n_644),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_629),
.A2(n_633),
.B(n_620),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_690),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_724),
.A2(n_502),
.B(n_725),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_752),
.B(n_500),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_637),
.B(n_507),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_724),
.A2(n_620),
.B1(n_658),
.B2(n_644),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_730),
.A2(n_758),
.B(n_735),
.C(n_720),
.Y(n_939)
);

CKINVDCx10_ASAP7_75t_R g940 ( 
.A(n_754),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_678),
.B(n_321),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_629),
.B(n_547),
.C(n_416),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_752),
.B(n_500),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_658),
.A2(n_724),
.B(n_653),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_752),
.B(n_500),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_658),
.A2(n_724),
.B(n_653),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_752),
.B(n_500),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_724),
.A2(n_658),
.B(n_653),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_646),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_620),
.A2(n_759),
.B(n_731),
.C(n_622),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_678),
.B(n_321),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_752),
.B(n_500),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_724),
.A2(n_658),
.B(n_653),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_752),
.B(n_500),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_724),
.A2(n_658),
.B(n_653),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_678),
.B(n_321),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_644),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_917),
.A2(n_939),
.B(n_780),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_793),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_816),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_938),
.A2(n_821),
.B(n_866),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_916),
.A2(n_844),
.B(n_881),
.Y(n_962)
);

OAI22x1_ASAP7_75t_L g963 ( 
.A1(n_901),
.A2(n_869),
.B1(n_871),
.B2(n_909),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_852),
.A2(n_926),
.B(n_923),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_779),
.A2(n_930),
.B1(n_951),
.B2(n_956),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_931),
.B(n_781),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_807),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_881),
.A2(n_894),
.B(n_913),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_942),
.B(n_933),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_816),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_944),
.A2(n_946),
.B(n_925),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_894),
.A2(n_913),
.B(n_902),
.Y(n_972)
);

OAI21x1_ASAP7_75t_SL g973 ( 
.A1(n_875),
.A2(n_897),
.B(n_888),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_813),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_924),
.A2(n_928),
.B(n_925),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_829),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_870),
.A2(n_798),
.B(n_794),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_921),
.A2(n_952),
.B1(n_943),
.B2(n_947),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_924),
.A2(n_948),
.B(n_928),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_936),
.A2(n_945),
.B1(n_954),
.B2(n_899),
.Y(n_980)
);

AOI21x1_ASAP7_75t_SL g981 ( 
.A1(n_785),
.A2(n_879),
.B(n_826),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_948),
.A2(n_955),
.B(n_953),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_849),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_880),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_891),
.B(n_857),
.Y(n_985)
);

INVx3_ASAP7_75t_SL g986 ( 
.A(n_816),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_784),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_878),
.Y(n_988)
);

AO31x2_ASAP7_75t_L g989 ( 
.A1(n_789),
.A2(n_795),
.A3(n_897),
.B(n_873),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_782),
.B(n_860),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_825),
.Y(n_991)
);

AOI22x1_ASAP7_75t_L g992 ( 
.A1(n_953),
.A2(n_955),
.B1(n_809),
.B2(n_800),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_822),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_819),
.B(n_883),
.Y(n_994)
);

NOR2x1_ASAP7_75t_SL g995 ( 
.A(n_807),
.B(n_831),
.Y(n_995)
);

AND3x2_ASAP7_75t_L g996 ( 
.A(n_941),
.B(n_836),
.C(n_792),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_920),
.A2(n_950),
.B(n_882),
.C(n_887),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_810),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_830),
.A2(n_837),
.B(n_839),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_846),
.A2(n_896),
.B(n_780),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_902),
.A2(n_929),
.B(n_846),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_788),
.B(n_802),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_935),
.A2(n_918),
.B(n_823),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_896),
.A2(n_847),
.B(n_858),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_808),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_820),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_949),
.Y(n_1007)
);

AND3x4_ASAP7_75t_L g1008 ( 
.A(n_890),
.B(n_810),
.C(n_791),
.Y(n_1008)
);

AOI21x1_ASAP7_75t_L g1009 ( 
.A1(n_851),
.A2(n_914),
.B(n_858),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_898),
.A2(n_905),
.B(n_908),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_838),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_864),
.A2(n_892),
.B(n_886),
.Y(n_1012)
);

AO21x1_ASAP7_75t_L g1013 ( 
.A1(n_853),
.A2(n_859),
.B(n_889),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_787),
.A2(n_817),
.B(n_799),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_814),
.A2(n_812),
.B(n_862),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_885),
.A2(n_797),
.B(n_790),
.C(n_904),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_940),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_915),
.A2(n_884),
.B(n_854),
.C(n_867),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_806),
.A2(n_815),
.B(n_805),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_786),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_842),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_922),
.B(n_957),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_861),
.A2(n_850),
.B(n_855),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_876),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_893),
.B(n_895),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_857),
.A2(n_818),
.B1(n_841),
.B2(n_906),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_834),
.A2(n_863),
.B(n_868),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_786),
.B(n_856),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_910),
.B(n_911),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_843),
.A2(n_840),
.B(n_912),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_804),
.A2(n_934),
.B(n_877),
.Y(n_1031)
);

AOI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_828),
.A2(n_900),
.B(n_874),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_848),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_845),
.A2(n_811),
.B(n_934),
.Y(n_1034)
);

OA21x2_ASAP7_75t_L g1035 ( 
.A1(n_865),
.A2(n_824),
.B(n_833),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_801),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_907),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_803),
.A2(n_872),
.B(n_903),
.C(n_804),
.Y(n_1038)
);

CKINVDCx11_ASAP7_75t_R g1039 ( 
.A(n_827),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_783),
.A2(n_937),
.B(n_919),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_907),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_SL g1042 ( 
.A(n_906),
.B(n_808),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_907),
.B(n_808),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_906),
.B(n_856),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_872),
.A2(n_856),
.B(n_832),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_921),
.B(n_936),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_899),
.B(n_901),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_810),
.B(n_848),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_810),
.B(n_848),
.Y(n_1049)
);

AO31x2_ASAP7_75t_L g1050 ( 
.A1(n_821),
.A2(n_916),
.A3(n_939),
.B(n_917),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_786),
.B(n_690),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_835),
.A2(n_932),
.B(n_927),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_822),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_901),
.A2(n_626),
.B1(n_615),
.B2(n_931),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_921),
.B(n_936),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_835),
.A2(n_932),
.B(n_927),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_779),
.B(n_507),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_835),
.A2(n_932),
.B(n_927),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_779),
.A2(n_494),
.B1(n_507),
.B2(n_866),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_921),
.B(n_936),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_835),
.A2(n_932),
.B(n_927),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_793),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_779),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_816),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_835),
.A2(n_866),
.B(n_899),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_901),
.A2(n_869),
.B1(n_871),
.B2(n_695),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_808),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_SL g1068 ( 
.A(n_807),
.B(n_690),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_917),
.A2(n_939),
.B(n_780),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_917),
.A2(n_939),
.B(n_780),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_816),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_796),
.A2(n_916),
.B(n_844),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_821),
.A2(n_916),
.A3(n_939),
.B(n_917),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_931),
.B(n_615),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_813),
.Y(n_1075)
);

INVx3_ASAP7_75t_SL g1076 ( 
.A(n_816),
.Y(n_1076)
);

BUFx4f_ASAP7_75t_SL g1077 ( 
.A(n_822),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_807),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_921),
.B(n_936),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_917),
.B(n_939),
.C(n_866),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_813),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_835),
.A2(n_932),
.B(n_927),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_917),
.A2(n_939),
.B(n_780),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_835),
.A2(n_932),
.B(n_927),
.Y(n_1084)
);

AO21x1_ASAP7_75t_L g1085 ( 
.A1(n_835),
.A2(n_866),
.B(n_899),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_821),
.A2(n_916),
.A3(n_939),
.B(n_917),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_793),
.Y(n_1087)
);

NAND2x1_ASAP7_75t_L g1088 ( 
.A(n_807),
.B(n_690),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_921),
.B(n_936),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1074),
.B(n_966),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1057),
.B(n_1063),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_1005),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_987),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_978),
.B(n_1046),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1042),
.B(n_1044),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_994),
.A2(n_980),
.B(n_978),
.C(n_1084),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_974),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1011),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1077),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1002),
.B(n_1059),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_986),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_1028),
.B(n_1048),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_988),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1054),
.B(n_965),
.Y(n_1104)
);

AND2x6_ASAP7_75t_L g1105 ( 
.A(n_1020),
.B(n_1049),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1046),
.B(n_1055),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_991),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1055),
.B(n_1060),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1021),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1076),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1017),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1047),
.A2(n_985),
.B1(n_994),
.B2(n_980),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_1080),
.A2(n_1061),
.B(n_1084),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_970),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1060),
.B(n_1079),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1024),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_984),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1061),
.A2(n_1082),
.B(n_961),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_961),
.A2(n_964),
.B(n_999),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1047),
.A2(n_985),
.B1(n_1085),
.B2(n_1065),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1075),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_993),
.B(n_1053),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1079),
.B(n_1089),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1005),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_990),
.B(n_1089),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_970),
.B(n_960),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1081),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_SL g1129 ( 
.A1(n_1066),
.A2(n_963),
.B1(n_1083),
.B2(n_958),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_1007),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_997),
.A2(n_977),
.B(n_1016),
.C(n_990),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_998),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_977),
.A2(n_971),
.B(n_982),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1032),
.A2(n_1036),
.B1(n_1087),
.B2(n_976),
.Y(n_1134)
);

AND2x6_ASAP7_75t_L g1135 ( 
.A(n_967),
.B(n_1078),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_993),
.B(n_1053),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1022),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1043),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_1008),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1005),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1022),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_SL g1142 ( 
.A(n_1026),
.B(n_969),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1025),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_1039),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1067),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1067),
.B(n_1038),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1025),
.B(n_1033),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_982),
.A2(n_975),
.B(n_979),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1043),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_967),
.B(n_1078),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1032),
.A2(n_1062),
.B1(n_983),
.B2(n_1026),
.Y(n_1151)
);

INVx6_ASAP7_75t_SL g1152 ( 
.A(n_996),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1069),
.A2(n_1070),
.B1(n_1013),
.B2(n_1018),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_1004),
.A2(n_1000),
.B(n_962),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1006),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1045),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_1003),
.B(n_992),
.C(n_1014),
.Y(n_1157)
);

BUFx5_ASAP7_75t_L g1158 ( 
.A(n_1037),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1003),
.A2(n_1035),
.B1(n_1029),
.B2(n_1014),
.Y(n_1159)
);

AOI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_1019),
.A2(n_995),
.B1(n_973),
.B2(n_1040),
.C1(n_1041),
.C2(n_1068),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1034),
.B(n_1051),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1030),
.B(n_1050),
.Y(n_1162)
);

OAI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1019),
.A2(n_1009),
.B(n_1015),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1023),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1050),
.Y(n_1165)
);

OAI31xp33_ASAP7_75t_L g1166 ( 
.A1(n_981),
.A2(n_1050),
.A3(n_1073),
.B(n_1086),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1073),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1088),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1086),
.B(n_1035),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_989),
.B(n_1031),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_989),
.B(n_968),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1027),
.B(n_972),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1001),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1012),
.B(n_1010),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1072),
.B(n_1074),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1077),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1047),
.A2(n_901),
.B1(n_754),
.B2(n_321),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_974),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1077),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_994),
.A2(n_939),
.B(n_917),
.C(n_866),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_967),
.B(n_1078),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_974),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_988),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1077),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1080),
.A2(n_866),
.B1(n_980),
.B2(n_994),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_987),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1080),
.B(n_939),
.C(n_917),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_959),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1077),
.Y(n_1189)
);

AND2x6_ASAP7_75t_L g1190 ( 
.A(n_1044),
.B(n_901),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1057),
.B(n_978),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_965),
.B(n_1057),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1057),
.B(n_978),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1074),
.B(n_966),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_980),
.B(n_978),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1057),
.B(n_978),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1052),
.A2(n_1058),
.B(n_1056),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1052),
.A2(n_1058),
.B(n_1056),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_988),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1047),
.A2(n_985),
.B1(n_1057),
.B2(n_965),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_974),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_966),
.B(n_993),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1042),
.B(n_1044),
.Y(n_1203)
);

NAND2x1_ASAP7_75t_L g1204 ( 
.A(n_967),
.B(n_1078),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_987),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1074),
.B(n_966),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_988),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1098),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1148),
.A2(n_1119),
.B(n_1133),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1109),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1116),
.Y(n_1211)
);

BUFx2_ASAP7_75t_R g1212 ( 
.A(n_1199),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1143),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_SL g1214 ( 
.A(n_1139),
.Y(n_1214)
);

BUFx2_ASAP7_75t_R g1215 ( 
.A(n_1155),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1118),
.A2(n_1198),
.B(n_1197),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1093),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1202),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1121),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1127),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1106),
.B(n_1108),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1129),
.A2(n_1104),
.B1(n_1200),
.B2(n_1192),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1112),
.B(n_1195),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1099),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1115),
.B(n_1123),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1094),
.B(n_1191),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1174),
.A2(n_1172),
.B(n_1185),
.Y(n_1227)
);

AOI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1172),
.A2(n_1185),
.B(n_1161),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1129),
.A2(n_1142),
.B1(n_1196),
.B2(n_1193),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1200),
.A2(n_1112),
.B1(n_1190),
.B2(n_1177),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1147),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1167),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1171),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1190),
.A2(n_1195),
.B1(n_1120),
.B2(n_1100),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1190),
.A2(n_1120),
.B1(n_1091),
.B2(n_1187),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1146),
.B(n_1095),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1122),
.Y(n_1237)
);

CKINVDCx16_ASAP7_75t_R g1238 ( 
.A(n_1103),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1170),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1111),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1184),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1178),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1154),
.A2(n_1157),
.B(n_1169),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1190),
.A2(n_1187),
.B1(n_1134),
.B2(n_1152),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1152),
.A2(n_1090),
.B1(n_1206),
.B2(n_1194),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1182),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1146),
.B(n_1095),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1130),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1159),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1201),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1153),
.A2(n_1125),
.B1(n_1159),
.B2(n_1141),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1125),
.A2(n_1105),
.B1(n_1137),
.B2(n_1203),
.Y(n_1252)
);

CKINVDCx6p67_ASAP7_75t_R g1253 ( 
.A(n_1144),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1175),
.B(n_1156),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1164),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1180),
.A2(n_1131),
.B1(n_1153),
.B2(n_1096),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1183),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1176),
.B(n_1179),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1188),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1186),
.A2(n_1205),
.B1(n_1132),
.B2(n_1136),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1113),
.A2(n_1110),
.B1(n_1101),
.B2(n_1114),
.Y(n_1261)
);

INVxp67_ASAP7_75t_SL g1262 ( 
.A(n_1149),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1138),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1151),
.A2(n_1105),
.B1(n_1138),
.B2(n_1102),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_SL g1265 ( 
.A(n_1189),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1207),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1107),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1154),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1158),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1101),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1158),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1128),
.B(n_1117),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1114),
.A2(n_1150),
.B1(n_1126),
.B2(n_1128),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1158),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1092),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1135),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1166),
.A2(n_1173),
.B(n_1160),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1124),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_SL g1279 ( 
.A(n_1140),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1140),
.Y(n_1280)
);

CKINVDCx6p67_ASAP7_75t_R g1281 ( 
.A(n_1140),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1135),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1181),
.A2(n_1204),
.B(n_1166),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1145),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1158),
.A2(n_1160),
.B1(n_1145),
.B2(n_1173),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1168),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1104),
.A2(n_1047),
.B1(n_901),
.B2(n_985),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1106),
.B(n_1108),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1103),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1144),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1129),
.A2(n_1047),
.B1(n_901),
.B2(n_754),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1167),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1129),
.B(n_1146),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1099),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1148),
.A2(n_1119),
.B(n_1133),
.Y(n_1295)
);

BUFx2_ASAP7_75t_R g1296 ( 
.A(n_1199),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_SL g1297 ( 
.A(n_1144),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1097),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1097),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1129),
.A2(n_1047),
.B1(n_901),
.B2(n_754),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1097),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1097),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1106),
.B(n_1108),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1112),
.B(n_1195),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1129),
.A2(n_1047),
.B1(n_901),
.B2(n_754),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1148),
.A2(n_1119),
.B(n_1133),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1143),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1165),
.Y(n_1308)
);

AO21x1_ASAP7_75t_SL g1309 ( 
.A1(n_1226),
.A2(n_1285),
.B(n_1249),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1228),
.Y(n_1310)
);

INVxp33_ASAP7_75t_L g1311 ( 
.A(n_1265),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1213),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1276),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1308),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1251),
.A2(n_1268),
.B(n_1243),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1276),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1240),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1262),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1233),
.B(n_1223),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1307),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1231),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1233),
.B(n_1269),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1227),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1248),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1239),
.A2(n_1268),
.B(n_1249),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_SL g1326 ( 
.A(n_1257),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1218),
.Y(n_1327)
);

CKINVDCx16_ASAP7_75t_R g1328 ( 
.A(n_1279),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1269),
.B(n_1271),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1223),
.A2(n_1304),
.B(n_1256),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1232),
.B(n_1292),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1221),
.B(n_1225),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1288),
.B(n_1303),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1283),
.A2(n_1216),
.B(n_1306),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1208),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1210),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1258),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1211),
.B(n_1219),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1220),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1255),
.B(n_1237),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1242),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1229),
.A2(n_1222),
.B(n_1261),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1255),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1246),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1250),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1255),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1298),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1299),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1277),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1232),
.B(n_1292),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1277),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1301),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1302),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1263),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1277),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1254),
.B(n_1234),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1293),
.B(n_1276),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1293),
.B(n_1235),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1293),
.B(n_1209),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1278),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1240),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1209),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1216),
.A2(n_1306),
.B(n_1295),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1295),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1224),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1306),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1259),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1287),
.B(n_1247),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1286),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1319),
.B(n_1230),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1319),
.B(n_1282),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1314),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1364),
.A2(n_1300),
.B(n_1291),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1330),
.B(n_1282),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1330),
.B(n_1294),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1330),
.B(n_1260),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1360),
.B(n_1280),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1318),
.Y(n_1379)
);

AND2x2_ASAP7_75t_SL g1380 ( 
.A(n_1360),
.B(n_1305),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1331),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1351),
.Y(n_1382)
);

OAI31xp33_ASAP7_75t_L g1383 ( 
.A1(n_1359),
.A2(n_1244),
.A3(n_1273),
.B(n_1245),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1335),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1335),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1321),
.B(n_1217),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1325),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1336),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1322),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1312),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1315),
.B(n_1247),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1315),
.B(n_1322),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1320),
.B(n_1327),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1322),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1315),
.B(n_1217),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1343),
.B(n_1346),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1315),
.B(n_1236),
.Y(n_1397)
);

OAI211xp5_ASAP7_75t_L g1398 ( 
.A1(n_1342),
.A2(n_1252),
.B(n_1267),
.C(n_1270),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1332),
.A2(n_1272),
.B1(n_1264),
.B2(n_1214),
.C(n_1284),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1363),
.A2(n_1275),
.B(n_1236),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1355),
.B(n_1270),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1338),
.B(n_1281),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1366),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1390),
.B(n_1379),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1398),
.A2(n_1337),
.B(n_1324),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1398),
.A2(n_1333),
.B1(n_1340),
.B2(n_1355),
.C(n_1347),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1377),
.A2(n_1358),
.B1(n_1328),
.B2(n_1359),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1377),
.A2(n_1358),
.B(n_1310),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1383),
.A2(n_1311),
.B(n_1357),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_SL g1411 ( 
.A(n_1379),
.B(n_1316),
.Y(n_1411)
);

OA211x2_ASAP7_75t_L g1412 ( 
.A1(n_1383),
.A2(n_1328),
.B(n_1313),
.C(n_1316),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1380),
.A2(n_1358),
.B1(n_1316),
.B2(n_1313),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1376),
.B(n_1361),
.C(n_1339),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1381),
.B(n_1341),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1381),
.B(n_1341),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1395),
.B(n_1345),
.C(n_1354),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1380),
.A2(n_1309),
.B1(n_1357),
.B2(n_1369),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1382),
.B(n_1344),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1394),
.B(n_1372),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1395),
.B(n_1376),
.C(n_1401),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1395),
.B(n_1348),
.C(n_1354),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1376),
.B(n_1401),
.C(n_1396),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1380),
.A2(n_1386),
.B1(n_1404),
.B2(n_1402),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1394),
.B(n_1349),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_L g1428 ( 
.A(n_1401),
.B(n_1347),
.C(n_1345),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1375),
.A2(n_1392),
.B(n_1371),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1393),
.B(n_1353),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1372),
.B(n_1349),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1387),
.A2(n_1364),
.B(n_1334),
.Y(n_1432)
);

AOI211xp5_ASAP7_75t_L g1433 ( 
.A1(n_1375),
.A2(n_1369),
.B(n_1356),
.C(n_1323),
.Y(n_1433)
);

OAI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1399),
.A2(n_1350),
.B1(n_1352),
.B2(n_1368),
.C(n_1370),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1386),
.B(n_1317),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1378),
.B(n_1392),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1371),
.A2(n_1323),
.B(n_1310),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1374),
.B(n_1367),
.C(n_1370),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1429),
.B(n_1373),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1416),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1432),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1417),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1421),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1420),
.A2(n_1380),
.B1(n_1374),
.B2(n_1309),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1436),
.B(n_1400),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1436),
.B(n_1386),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1425),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1422),
.B(n_1391),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1422),
.B(n_1391),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1415),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1418),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1428),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1424),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1430),
.B(n_1371),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1415),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1423),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1426),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1437),
.B(n_1384),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1414),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1419),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1438),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1441),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1445),
.A2(n_1374),
.B1(n_1407),
.B2(n_1412),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1453),
.B(n_1435),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1449),
.B(n_1431),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1462),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1459),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1462),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1449),
.B(n_1431),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1440),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1441),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1454),
.B(n_1438),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1440),
.Y(n_1476)
);

NOR2xp67_ASAP7_75t_L g1477 ( 
.A(n_1462),
.B(n_1409),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1326),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1454),
.B(n_1385),
.Y(n_1479)
);

INVxp33_ASAP7_75t_L g1480 ( 
.A(n_1448),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1458),
.B(n_1419),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1443),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1458),
.B(n_1427),
.Y(n_1483)
);

AOI211xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1451),
.A2(n_1297),
.B(n_1413),
.C(n_1410),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1443),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1456),
.B(n_1403),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1452),
.B(n_1385),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1452),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1452),
.B(n_1388),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1444),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1488),
.B(n_1456),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_SL g1492 ( 
.A(n_1480),
.B(n_1448),
.C(n_1451),
.Y(n_1492)
);

NOR2x1_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1257),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1479),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1472),
.B(n_1473),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1488),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1463),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1461),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1457),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1480),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1475),
.B(n_1455),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1475),
.B(n_1455),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1478),
.B(n_1238),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1487),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1447),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1467),
.B(n_1457),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1475),
.B(n_1439),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1481),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1489),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1290),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1489),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1478),
.B(n_1362),
.Y(n_1516)
);

OAI31xp33_ASAP7_75t_L g1517 ( 
.A1(n_1484),
.A2(n_1408),
.A3(n_1439),
.B(n_1434),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1471),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1471),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1467),
.B(n_1442),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1476),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1469),
.B(n_1442),
.Y(n_1522)
);

NAND2xp33_ASAP7_75t_L g1523 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1523)
);

OR2x6_ASAP7_75t_L g1524 ( 
.A(n_1468),
.B(n_1290),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1482),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1485),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1485),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1481),
.B(n_1447),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1468),
.B(n_1446),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1503),
.B(n_1469),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1497),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1524),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1518),
.Y(n_1536)
);

AO21x2_ASAP7_75t_L g1537 ( 
.A1(n_1492),
.A2(n_1474),
.B(n_1463),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1531),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1519),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1524),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1495),
.B(n_1483),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1516),
.B(n_1253),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1495),
.B(n_1483),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1521),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1504),
.B(n_1510),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1509),
.B(n_1486),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1493),
.B(n_1496),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1496),
.B(n_1466),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1524),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1517),
.A2(n_1464),
.B1(n_1397),
.B2(n_1374),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1525),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1499),
.B(n_1466),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1526),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1527),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1524),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1512),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1499),
.B(n_1466),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1500),
.B(n_1470),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1502),
.A2(n_1464),
.B1(n_1406),
.B2(n_1412),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1501),
.B(n_1490),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1498),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1494),
.Y(n_1564)
);

AO21x2_ASAP7_75t_L g1565 ( 
.A1(n_1491),
.A2(n_1474),
.B(n_1463),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1502),
.B(n_1490),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1498),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1550),
.A2(n_1511),
.B1(n_1514),
.B2(n_1531),
.Y(n_1568)
);

NAND4xp25_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1484),
.C(n_1505),
.D(n_1516),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_L g1570 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1556),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1561),
.B(n_1511),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1561),
.B(n_1505),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1536),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1537),
.A2(n_1522),
.B1(n_1513),
.B2(n_1507),
.C(n_1515),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1537),
.A2(n_1523),
.B(n_1514),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1537),
.A2(n_1500),
.B1(n_1514),
.B2(n_1531),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1543),
.B(n_1506),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1536),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1542),
.B(n_1253),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1508),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1537),
.A2(n_1523),
.B(n_1514),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1557),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1508),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1556),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1548),
.B(n_1530),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1545),
.B(n_1530),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1539),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1557),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1535),
.B(n_1289),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1556),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1539),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1590),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1574),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1579),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1587),
.B(n_1545),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1552),
.Y(n_1598)
);

NOR2xp67_ASAP7_75t_SL g1599 ( 
.A(n_1572),
.B(n_1538),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1552),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1588),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1592),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1591),
.B(n_1558),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1577),
.B(n_1535),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1583),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1589),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1590),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1570),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1609),
.A2(n_1572),
.B1(n_1573),
.B2(n_1568),
.Y(n_1612)
);

NAND4xp25_ASAP7_75t_L g1613 ( 
.A(n_1598),
.B(n_1573),
.C(n_1575),
.D(n_1569),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1599),
.A2(n_1582),
.B(n_1576),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1608),
.A2(n_1549),
.B1(n_1540),
.B2(n_1534),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1605),
.A2(n_1580),
.B(n_1566),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1593),
.B(n_1580),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1599),
.A2(n_1540),
.B1(n_1549),
.B2(n_1565),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1597),
.Y(n_1619)
);

NOR3x1_ASAP7_75t_L g1620 ( 
.A(n_1602),
.B(n_1533),
.C(n_1532),
.Y(n_1620)
);

NAND4xp25_ASAP7_75t_SL g1621 ( 
.A(n_1597),
.B(n_1559),
.C(n_1532),
.D(n_1533),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1605),
.Y(n_1622)
);

AOI21xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1604),
.A2(n_1538),
.B(n_1534),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1622),
.B(n_1607),
.C(n_1606),
.Y(n_1624)
);

NOR3x1_ASAP7_75t_L g1625 ( 
.A(n_1613),
.B(n_1611),
.C(n_1596),
.Y(n_1625)
);

NOR4xp25_ASAP7_75t_L g1626 ( 
.A(n_1612),
.B(n_1595),
.C(n_1594),
.D(n_1601),
.Y(n_1626)
);

AND5x1_ASAP7_75t_L g1627 ( 
.A(n_1617),
.B(n_1616),
.C(n_1618),
.D(n_1621),
.E(n_1620),
.Y(n_1627)
);

OA22x2_ASAP7_75t_L g1628 ( 
.A1(n_1614),
.A2(n_1611),
.B1(n_1610),
.B2(n_1600),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1623),
.B(n_1596),
.Y(n_1629)
);

NOR3xp33_ASAP7_75t_L g1630 ( 
.A(n_1615),
.B(n_1603),
.C(n_1619),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1619),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1614),
.B(n_1266),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_L g1633 ( 
.A(n_1614),
.B(n_1266),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1626),
.B(n_1538),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1629),
.A2(n_1562),
.B(n_1538),
.C(n_1546),
.Y(n_1635)
);

NAND4xp25_ASAP7_75t_L g1636 ( 
.A(n_1625),
.B(n_1624),
.C(n_1630),
.D(n_1632),
.Y(n_1636)
);

AND4x2_ASAP7_75t_L g1637 ( 
.A(n_1633),
.B(n_1600),
.C(n_1212),
.D(n_1296),
.Y(n_1637)
);

AOI211xp5_ASAP7_75t_L g1638 ( 
.A1(n_1627),
.A2(n_1564),
.B(n_1546),
.C(n_1554),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1631),
.B(n_1534),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1634),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1639),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1638),
.A2(n_1628),
.B1(n_1635),
.B2(n_1564),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1636),
.B(n_1289),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1637),
.A2(n_1565),
.B1(n_1567),
.B2(n_1563),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1636),
.B(n_1544),
.Y(n_1645)
);

AND4x1_ASAP7_75t_L g1646 ( 
.A(n_1643),
.B(n_1215),
.C(n_1551),
.D(n_1560),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1640),
.Y(n_1647)
);

XOR2x1_ASAP7_75t_L g1648 ( 
.A(n_1641),
.B(n_1534),
.Y(n_1648)
);

NOR4xp25_ASAP7_75t_L g1649 ( 
.A(n_1642),
.B(n_1645),
.C(n_1644),
.D(n_1544),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1640),
.B(n_1551),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1648),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1647),
.Y(n_1652)
);

XNOR2xp5_ASAP7_75t_L g1653 ( 
.A(n_1646),
.B(n_1563),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1651),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1654),
.Y(n_1655)
);

OAI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1653),
.B(n_1651),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1655),
.A2(n_1652),
.B1(n_1650),
.B2(n_1649),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1657),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1656),
.Y(n_1659)
);

OR2x6_ASAP7_75t_L g1660 ( 
.A(n_1659),
.B(n_1241),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1658),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1661),
.Y(n_1662)
);

AOI322xp5_ASAP7_75t_L g1663 ( 
.A1(n_1662),
.A2(n_1660),
.A3(n_1567),
.B1(n_1563),
.B2(n_1553),
.C1(n_1554),
.C2(n_1560),
.Y(n_1663)
);

OAI221xp5_ASAP7_75t_R g1664 ( 
.A1(n_1663),
.A2(n_1565),
.B1(n_1553),
.B2(n_1555),
.C(n_1241),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1555),
.B(n_1567),
.C(n_1241),
.Y(n_1665)
);


endmodule