module real_aes_6036_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_13;
wire n_7;
wire n_8;
wire n_12;
wire n_9;
wire n_10;
wire n_11;
NOR2xp33_ASAP7_75t_L g7 ( .A(n_0), .B(n_8), .Y(n_7) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_2), .B(n_13), .Y(n_12) );
BUFx3_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
A2O1A1Ixp33_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_7), .B(n_10), .C(n_12), .Y(n_6) );
NOR2xp33_ASAP7_75t_SL g10 ( .A(n_7), .B(n_11), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_9), .Y(n_8) );
endmodule