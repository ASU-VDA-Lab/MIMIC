module fake_netlist_5_1591_n_2382 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_382, n_554, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2382);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2382;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_832;
wire n_857;
wire n_2305;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_1849;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_602;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_684;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_703;
wire n_1115;
wire n_698;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

INVx3_ASAP7_75t_L g578 ( 
.A(n_515),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_158),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_175),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_349),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_281),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_348),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_190),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_357),
.Y(n_586)
);

NOR2xp67_ASAP7_75t_L g587 ( 
.A(n_183),
.B(n_264),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_397),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_251),
.Y(n_589)
);

INVxp67_ASAP7_75t_SL g590 ( 
.A(n_135),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_284),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_565),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_290),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_233),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_237),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_159),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_74),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_484),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_185),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_170),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_507),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_66),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_45),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_203),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_235),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_361),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_395),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_20),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_76),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_417),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_249),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_33),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_559),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_20),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_424),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_307),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_467),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_287),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_420),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_202),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_491),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_157),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_295),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_494),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_65),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_18),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_222),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_53),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_105),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_473),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_434),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_324),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_350),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_188),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_196),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_166),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_239),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_165),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_499),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_5),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_472),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_471),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_299),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_375),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_122),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_224),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_301),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_528),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_205),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_317),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_452),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_219),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_269),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_382),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_509),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_190),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_226),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_83),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_74),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_94),
.Y(n_661)
);

INVxp33_ASAP7_75t_SL g662 ( 
.A(n_568),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_180),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_148),
.Y(n_664)
);

CKINVDCx14_ASAP7_75t_R g665 ( 
.A(n_356),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_449),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_70),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_319),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_197),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_502),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_192),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_535),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_183),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_203),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_55),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_549),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_112),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_429),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_78),
.Y(n_679)
);

CKINVDCx16_ASAP7_75t_R g680 ( 
.A(n_139),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_119),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_41),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_105),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_182),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_139),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_111),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_1),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_288),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_460),
.Y(n_689)
);

CKINVDCx14_ASAP7_75t_R g690 ( 
.A(n_485),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_506),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_45),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_511),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_441),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_543),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_107),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_279),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_230),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_84),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_182),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_392),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_175),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_305),
.Y(n_703)
);

CKINVDCx14_ASAP7_75t_R g704 ( 
.A(n_273),
.Y(n_704)
);

INVxp33_ASAP7_75t_L g705 ( 
.A(n_118),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_440),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_81),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_163),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_260),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_520),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_521),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_250),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_124),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_205),
.B(n_314),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_176),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_554),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_341),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_3),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_534),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_406),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_75),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_120),
.Y(n_722)
);

CKINVDCx14_ASAP7_75t_R g723 ( 
.A(n_409),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_2),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_450),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_128),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_456),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_178),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_475),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_255),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_570),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_28),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_453),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_390),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_500),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_530),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_318),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_438),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_479),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_546),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_481),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_55),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_268),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_433),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_514),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_285),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_208),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_283),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_517),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_323),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_194),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_418),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_337),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_153),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_165),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_127),
.Y(n_756)
);

BUFx10_ASAP7_75t_L g757 ( 
.A(n_333),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_461),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_282),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_416),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_18),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_212),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_41),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_310),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_498),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_236),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_487),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_223),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_114),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_326),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_60),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_468),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_325),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_322),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_553),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_501),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_27),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_241),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_490),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_199),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_469),
.B(n_504),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_184),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_207),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_370),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_85),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_414),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_311),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_33),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_303),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_88),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_198),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_411),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_206),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_328),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_274),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_122),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_308),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_258),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_186),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_202),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_437),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_84),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_369),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_24),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_388),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_64),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_57),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_480),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_245),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_519),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_257),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_60),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_567),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_91),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_362),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_489),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_387),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_272),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_94),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_85),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_505),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_419),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_291),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_286),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_270),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_169),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_210),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_573),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_422),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_238),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_555),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_342),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_256),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_306),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_133),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_189),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_289),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_410),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_253),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_378),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_338),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_2),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_146),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_336),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_213),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_443),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_483),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_320),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_330),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_82),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_561),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_36),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_510),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_16),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_451),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_201),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_204),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_470),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_114),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_108),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_129),
.Y(n_861)
);

CKINVDCx14_ASAP7_75t_R g862 ( 
.A(n_39),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_566),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_9),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_407),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_262),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_444),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_518),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_93),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_436),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_37),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_347),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_430),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_380),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_244),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_192),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_486),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_508),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_59),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_332),
.Y(n_880)
);

CKINVDCx16_ASAP7_75t_R g881 ( 
.A(n_75),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_386),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_246),
.B(n_389),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_266),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_391),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_22),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_385),
.B(n_297),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_29),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_78),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_503),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_560),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_353),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_177),
.B(n_557),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_196),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_156),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_551),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_179),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_360),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_275),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_454),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_153),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_149),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_191),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_377),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_187),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_545),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_540),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_254),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_145),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_126),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_376),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_529),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_252),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_118),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_136),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_143),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_313),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_125),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_123),
.Y(n_919)
);

BUFx5_ASAP7_75t_L g920 ( 
.A(n_556),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_558),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_372),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_525),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_200),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_44),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_79),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_572),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_496),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_394),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_117),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_280),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_435),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_157),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_62),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_73),
.Y(n_935)
);

CKINVDCx16_ASAP7_75t_R g936 ( 
.A(n_355),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_4),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_526),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_119),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_152),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_53),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_221),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_345),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_466),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_141),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_4),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_50),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_365),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_547),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_189),
.B(n_209),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_160),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_278),
.Y(n_952)
);

BUFx10_ASAP7_75t_L g953 ( 
.A(n_459),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_127),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_159),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_130),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_300),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_552),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_82),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_527),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_50),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_292),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_21),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_393),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_99),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_462),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_140),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_265),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_346),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_533),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_199),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_56),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_193),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_195),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_113),
.Y(n_975)
);

BUFx5_ASAP7_75t_L g976 ( 
.A(n_343),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_201),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_64),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_48),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_37),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_247),
.Y(n_981)
);

BUFx8_ASAP7_75t_SL g982 ( 
.A(n_398),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_335),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_52),
.Y(n_984)
);

CKINVDCx14_ASAP7_75t_R g985 ( 
.A(n_11),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_24),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_181),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_188),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_421),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_351),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_170),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_331),
.Y(n_992)
);

INVxp33_ASAP7_75t_L g993 ( 
.A(n_31),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_187),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_10),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_169),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_476),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_294),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_605),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_625),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_661),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_625),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_708),
.Y(n_1003)
);

AND2x2_ASAP7_75t_R g1004 ( 
.A(n_862),
.B(n_0),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_684),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_661),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_654),
.Y(n_1007)
);

INVx6_ASAP7_75t_L g1008 ( 
.A(n_757),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_621),
.B(n_624),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_860),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_635),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_860),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_757),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_708),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_860),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_837),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_935),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_935),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_935),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_667),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_862),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_680),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_881),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_621),
.B(n_624),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_604),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_920),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_SL g1027 ( 
.A1(n_580),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_706),
.B(n_6),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_706),
.B(n_7),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_614),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_837),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_920),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_724),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_615),
.B(n_8),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_615),
.B(n_646),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_614),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_578),
.A2(n_214),
.B(n_211),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_712),
.B(n_8),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_920),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_751),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_920),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_646),
.B(n_9),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_920),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_712),
.B(n_775),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_579),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_920),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_711),
.B(n_10),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_985),
.B(n_11),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_976),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_751),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_804),
.Y(n_1051)
);

OAI22x1_ASAP7_75t_SL g1052 ( 
.A1(n_602),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_804),
.Y(n_1053)
);

CKINVDCx16_ASAP7_75t_R g1054 ( 
.A(n_588),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_585),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_596),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_619),
.A2(n_216),
.B(n_215),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_597),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_605),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_985),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_941),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_634),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_991),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_991),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_665),
.B(n_15),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_605),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_664),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_665),
.B(n_15),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_651),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_592),
.B(n_16),
.Y(n_1070)
);

OA21x2_ASAP7_75t_L g1071 ( 
.A1(n_737),
.A2(n_17),
.B(n_19),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_651),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_787),
.B(n_17),
.Y(n_1073)
);

BUFx12f_ASAP7_75t_L g1074 ( 
.A(n_634),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_982),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_603),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_612),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_651),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_690),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_950),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_711),
.B(n_26),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_690),
.B(n_27),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_626),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_704),
.A2(n_723),
.B1(n_993),
.B2(n_705),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_636),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_651),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_976),
.Y(n_1087)
);

BUFx8_ASAP7_75t_L g1088 ( 
.A(n_688),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_851),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_704),
.B(n_723),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_976),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_623),
.A2(n_218),
.B(n_217),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_802),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_599),
.Y(n_1094)
);

OA21x2_ASAP7_75t_L g1095 ( 
.A1(n_737),
.A2(n_29),
.B(n_30),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_586),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_976),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_593),
.B(n_30),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_779),
.B(n_31),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_658),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_976),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_953),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_779),
.B(n_795),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_795),
.B(n_32),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_645),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_658),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_826),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_902),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_930),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_951),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_600),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_658),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_956),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_776),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_650),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_953),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_657),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_673),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_677),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_960),
.B(n_34),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_581),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_682),
.Y(n_1122)
);

OAI22x1_ASAP7_75t_SL g1123 ( 
.A1(n_620),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_832),
.B(n_38),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_844),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_666),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_582),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_685),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_844),
.B(n_39),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_666),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_686),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_666),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_666),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_687),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_700),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_702),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_583),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_718),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_721),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_705),
.B(n_40),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_722),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_993),
.B(n_40),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_732),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_608),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_832),
.B(n_42),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_609),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_865),
.B(n_42),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_742),
.Y(n_1148)
);

OAI21xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1035),
.A2(n_1103),
.B(n_1048),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1010),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1012),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1012),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1001),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1090),
.B(n_694),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1006),
.Y(n_1155)
);

OR2x6_ASAP7_75t_L g1156 ( 
.A(n_1144),
.B(n_638),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1008),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1069),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1069),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1018),
.Y(n_1160)
);

INVxp67_ASAP7_75t_R g1161 ( 
.A(n_1065),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1019),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1072),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1062),
.B(n_1074),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1072),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_1140),
.B(n_917),
.C(n_865),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1008),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1121),
.B(n_632),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1078),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1127),
.B(n_734),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1068),
.A2(n_910),
.B1(n_796),
.B2(n_632),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1086),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1015),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1137),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1013),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1112),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1054),
.B(n_870),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1045),
.B(n_917),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_SL g1179 ( 
.A(n_1016),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1015),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1017),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1126),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1009),
.B(n_749),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1017),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1009),
.B(n_874),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_SL g1186 ( 
.A(n_1031),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1030),
.B(n_747),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1024),
.B(n_877),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1024),
.B(n_877),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1082),
.B(n_639),
.Y(n_1190)
);

CKINVDCx6p67_ASAP7_75t_R g1191 ( 
.A(n_1102),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1142),
.A2(n_996),
.B1(n_995),
.B2(n_756),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1055),
.B(n_936),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1040),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_L g1195 ( 
.A(n_1084),
.B(n_987),
.C(n_640),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1044),
.B(n_929),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1040),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1036),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1126),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1125),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1116),
.B(n_587),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1089),
.B(n_714),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1056),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1034),
.B(n_988),
.C(n_628),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1130),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1130),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1050),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1050),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1094),
.B(n_649),
.Y(n_1209)
);

BUFx8_ASAP7_75t_SL g1210 ( 
.A(n_1075),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1132),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1132),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1133),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1000),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1053),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1026),
.A2(n_589),
.B(n_584),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1061),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1117),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1061),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1146),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1064),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1117),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_1096),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1118),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1011),
.B(n_699),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1059),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1118),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1119),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1100),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1111),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1119),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1120),
.B(n_662),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1106),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1115),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1122),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1131),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1135),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1138),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_1022),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1139),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_999),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1014),
.B(n_768),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1093),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_SL g1244 ( 
.A(n_1028),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_L g1245 ( 
.A(n_1042),
.B(n_994),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1028),
.B(n_893),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1141),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1047),
.B(n_730),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1143),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1020),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1076),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_1023),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1077),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1057),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1111),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1085),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1105),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1134),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1081),
.B(n_1099),
.Y(n_1259)
);

NOR3xp33_ASAP7_75t_L g1260 ( 
.A(n_1070),
.B(n_726),
.C(n_590),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1104),
.B(n_1145),
.C(n_1124),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1005),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1063),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1029),
.B(n_810),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1147),
.B(n_818),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1029),
.B(n_890),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1002),
.Y(n_1267)
);

INVx5_ASAP7_75t_L g1268 ( 
.A(n_999),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1098),
.A2(n_607),
.B1(n_611),
.B2(n_594),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1003),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1032),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1039),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1107),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1041),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1038),
.B(n_906),
.Y(n_1275)
);

INVx5_ASAP7_75t_L g1276 ( 
.A(n_999),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1043),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1046),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1108),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1033),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1049),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1051),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1087),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1092),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_1083),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1091),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1128),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1128),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1097),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1148),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1148),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1101),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1136),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_SL g1294 ( 
.A(n_1073),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1058),
.Y(n_1295)
);

BUFx4f_ASAP7_75t_L g1296 ( 
.A(n_1071),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1073),
.B(n_622),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1066),
.B(n_943),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_1129),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1025),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1005),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1025),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1129),
.B(n_629),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1067),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1067),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1021),
.A2(n_946),
.B1(n_959),
.B2(n_876),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1004),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1071),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1109),
.Y(n_1309)
);

INVxp33_ASAP7_75t_L g1310 ( 
.A(n_1109),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1007),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1110),
.B(n_598),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1007),
.B(n_660),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1113),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1095),
.A2(n_979),
.B1(n_771),
.B2(n_800),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1037),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1060),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1114),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1088),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1088),
.B(n_601),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1079),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1027),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1080),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1052),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1123),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1010),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1010),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1121),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1001),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1010),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1054),
.B(n_663),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1001),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1121),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1010),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1011),
.B(n_777),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1008),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_L g1337 ( 
.A(n_1065),
.B(n_669),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1090),
.B(n_606),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1010),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1035),
.B(n_992),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1010),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1054),
.B(n_671),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_1075),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1010),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1054),
.B(n_674),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1010),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1010),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1010),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1001),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1096),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1090),
.B(n_591),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1121),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1008),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1001),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1001),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1010),
.Y(n_1356)
);

NOR2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1116),
.B(n_781),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1010),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1035),
.B(n_643),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1010),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1090),
.B(n_610),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1001),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1001),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1010),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1121),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1137),
.Y(n_1366)
);

AND3x2_ASAP7_75t_L g1367 ( 
.A(n_1048),
.B(n_883),
.C(n_727),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1010),
.Y(n_1368)
);

CKINVDCx6p67_ASAP7_75t_R g1369 ( 
.A(n_1102),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1010),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1001),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1001),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1010),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1010),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1008),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1001),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1090),
.B(n_595),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1010),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1054),
.B(n_675),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1035),
.B(n_698),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1035),
.B(n_766),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1054),
.B(n_679),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1054),
.B(n_681),
.Y(n_1383)
);

CKINVDCx6p67_ASAP7_75t_R g1384 ( 
.A(n_1102),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1001),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_L g1386 ( 
.A(n_1065),
.B(n_683),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1008),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1048),
.B(n_659),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1010),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1001),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1010),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1010),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1001),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1010),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1010),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1037),
.A2(n_616),
.B(n_613),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1010),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1011),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1010),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1054),
.B(n_692),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1010),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1010),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1026),
.A2(n_631),
.B(n_627),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1054),
.B(n_696),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1010),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1001),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1001),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1010),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1121),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1010),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1090),
.B(n_633),
.Y(n_1411)
);

OAI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1318),
.A2(n_713),
.B1(n_728),
.B2(n_715),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1259),
.B(n_617),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1267),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1248),
.B(n_822),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1263),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1265),
.B(n_1232),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1168),
.B(n_830),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1209),
.B(n_707),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1270),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1280),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1351),
.B(n_618),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1282),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1340),
.A2(n_761),
.B1(n_814),
.B2(n_807),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1256),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1225),
.B(n_754),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1377),
.B(n_630),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1199),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1205),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1170),
.B(n_813),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1165),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1239),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1359),
.B(n_969),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1239),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1226),
.B(n_641),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1252),
.Y(n_1436)
);

AND2x2_ASAP7_75t_SL g1437 ( 
.A(n_1269),
.B(n_887),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1438)
);

XNOR2xp5_ASAP7_75t_L g1439 ( 
.A(n_1350),
.B(n_911),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_L g1440 ( 
.A(n_1156),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1233),
.B(n_644),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1233),
.B(n_647),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1190),
.B(n_656),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1190),
.B(n_1154),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1271),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1193),
.B(n_928),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1200),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1214),
.B(n_1338),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1398),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1153),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1155),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1296),
.A2(n_1246),
.B(n_1361),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1272),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1157),
.B(n_755),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1353),
.B(n_763),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1411),
.B(n_691),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1333),
.B(n_769),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1274),
.Y(n_1458)
);

AO221x1_ASAP7_75t_L g1459 ( 
.A1(n_1306),
.A2(n_880),
.B1(n_885),
.B2(n_848),
.C(n_731),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1261),
.B(n_697),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1277),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1203),
.B(n_739),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1165),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1255),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1278),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1281),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1283),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1252),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1188),
.B(n_719),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1286),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1166),
.A2(n_782),
.B1(n_783),
.B2(n_780),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1189),
.B(n_720),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1196),
.B(n_729),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1160),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1174),
.B(n_852),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1365),
.B(n_785),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1289),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1262),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1183),
.B(n_733),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1230),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1292),
.Y(n_1481)
);

AND2x6_ASAP7_75t_SL g1482 ( 
.A(n_1324),
.B(n_859),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1365),
.B(n_788),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1185),
.B(n_735),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1220),
.B(n_738),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1149),
.B(n_790),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1162),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1329),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1171),
.B(n_740),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1301),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1285),
.B(n_791),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1264),
.B(n_1266),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1332),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1335),
.Y(n_1494)
);

OAI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1192),
.A2(n_871),
.B1(n_879),
.B2(n_864),
.C(n_861),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1357),
.B(n_1244),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1161),
.B(n_1178),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1198),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1287),
.Y(n_1499)
);

INVx8_ASAP7_75t_L g1500 ( 
.A(n_1210),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1388),
.A2(n_883),
.B1(n_744),
.B2(n_746),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1164),
.B(n_886),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1275),
.B(n_793),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1323),
.B(n_799),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1175),
.B(n_758),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1229),
.B(n_748),
.Y(n_1506)
);

INVx8_ASAP7_75t_L g1507 ( 
.A(n_1328),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1310),
.B(n_806),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1315),
.A2(n_901),
.B1(n_905),
.B2(n_897),
.Y(n_1509)
);

CKINVDCx16_ASAP7_75t_R g1510 ( 
.A(n_1223),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1352),
.B(n_762),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_L g1512 ( 
.A(n_1308),
.B(n_731),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1409),
.B(n_778),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1299),
.B(n_812),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1331),
.B(n_819),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1366),
.B(n_915),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1349),
.B(n_772),
.Y(n_1517)
);

NOR2xp67_ASAP7_75t_L g1518 ( 
.A(n_1167),
.B(n_774),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_L g1519 ( 
.A(n_1308),
.B(n_731),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1288),
.Y(n_1520)
);

AOI22x1_ASAP7_75t_L g1521 ( 
.A1(n_1316),
.A2(n_642),
.B1(n_648),
.B2(n_637),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1354),
.B(n_784),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1355),
.B(n_786),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1260),
.B(n_986),
.C(n_984),
.Y(n_1524)
);

NOR3xp33_ASAP7_75t_L g1525 ( 
.A(n_1195),
.B(n_926),
.C(n_919),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1215),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1297),
.B(n_820),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1299),
.B(n_803),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1362),
.B(n_789),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1363),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1342),
.B(n_835),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1317),
.A2(n_940),
.B1(n_945),
.B2(n_937),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1345),
.B(n_836),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1371),
.B(n_794),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1379),
.B(n_842),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1382),
.B(n_843),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1367),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1177),
.B(n_808),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1372),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1343),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1245),
.A2(n_798),
.B1(n_801),
.B2(n_797),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1376),
.B(n_816),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1337),
.A2(n_823),
.B1(n_824),
.B2(n_821),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1187),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1303),
.B(n_850),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1386),
.A2(n_653),
.B(n_652),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1383),
.B(n_854),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1290),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1268),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1321),
.A2(n_965),
.B1(n_971),
.B2(n_955),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1291),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1336),
.B(n_1375),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_L g1553 ( 
.A(n_1308),
.B(n_731),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1187),
.Y(n_1554)
);

NOR2xp67_ASAP7_75t_L g1555 ( 
.A(n_1387),
.B(n_825),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_SL g1556 ( 
.A(n_1343),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1213),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1221),
.B(n_973),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1204),
.B(n_827),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1319),
.B(n_828),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1201),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1385),
.B(n_829),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1213),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1400),
.B(n_856),
.Y(n_1564)
);

NOR2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1319),
.B(n_857),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1158),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1316),
.A2(n_668),
.B(n_670),
.C(n_655),
.Y(n_1567)
);

O2A1O1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1218),
.A2(n_975),
.B(n_998),
.C(n_676),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1298),
.A2(n_678),
.B(n_672),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1158),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1404),
.A2(n_833),
.B1(n_838),
.B2(n_831),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1202),
.B(n_997),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1217),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1321),
.A2(n_880),
.B1(n_885),
.B2(n_848),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1159),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1243),
.B(n_1273),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1244),
.B(n_869),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1217),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1390),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1219),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1163),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1294),
.B(n_888),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1393),
.B(n_849),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1320),
.B(n_855),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1311),
.B(n_924),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1294),
.B(n_889),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1313),
.A2(n_872),
.B1(n_878),
.B2(n_867),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1406),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1242),
.B(n_894),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1324),
.B(n_903),
.C(n_895),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1360),
.B(n_882),
.Y(n_1591)
);

NOR3xp33_ASAP7_75t_L g1592 ( 
.A(n_1325),
.B(n_914),
.C(n_909),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1191),
.B(n_961),
.Y(n_1593)
);

AND2x4_ASAP7_75t_SL g1594 ( 
.A(n_1369),
.B(n_974),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1156),
.A2(n_896),
.B1(n_898),
.B2(n_891),
.Y(n_1595)
);

INVx8_ASAP7_75t_L g1596 ( 
.A(n_1164),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1407),
.B(n_900),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1307),
.A2(n_1186),
.B1(n_1179),
.B2(n_1396),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1360),
.B(n_904),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1396),
.A2(n_880),
.B1(n_885),
.B2(n_848),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1322),
.A2(n_693),
.B1(n_695),
.B2(n_689),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1169),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1216),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1173),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1194),
.B(n_701),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1169),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1180),
.B(n_908),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1181),
.B(n_913),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1184),
.B(n_921),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1172),
.B(n_923),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1403),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1176),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1206),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1182),
.B(n_942),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1211),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1384),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1197),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1212),
.B(n_916),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1327),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_L g1620 ( 
.A(n_1268),
.B(n_944),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1234),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1182),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1235),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1273),
.B(n_918),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1236),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1312),
.A2(n_709),
.B(n_703),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_SL g1627 ( 
.A(n_1325),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1250),
.B(n_948),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1334),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1179),
.A2(n_957),
.B1(n_962),
.B2(n_952),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1268),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1251),
.A2(n_933),
.B1(n_934),
.B2(n_925),
.Y(n_1632)
);

INVxp33_ASAP7_75t_L g1633 ( 
.A(n_1207),
.Y(n_1633)
);

NOR2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1208),
.B(n_939),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1241),
.B(n_966),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1237),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1279),
.B(n_968),
.Y(n_1637)
);

AND2x6_ASAP7_75t_SL g1638 ( 
.A(n_1295),
.B(n_710),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1238),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1240),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1247),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1249),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1241),
.B(n_970),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_L g1644 ( 
.A(n_1293),
.B(n_954),
.C(n_947),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_SL g1645 ( 
.A(n_1253),
.B(n_980),
.C(n_977),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1150),
.B(n_1151),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1344),
.B(n_963),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1254),
.A2(n_717),
.B(n_716),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1186),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1346),
.B(n_967),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1257),
.A2(n_983),
.B1(n_989),
.B2(n_981),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1346),
.B(n_725),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1356),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1258),
.B(n_972),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1276),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1150),
.B(n_736),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1417),
.B(n_1284),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1576),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1433),
.B(n_1284),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1438),
.B(n_978),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1512),
.A2(n_1553),
.B(n_1519),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1526),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1437),
.A2(n_743),
.B1(n_745),
.B2(n_741),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1415),
.B(n_750),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1600),
.A2(n_753),
.B1(n_759),
.B2(n_752),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1452),
.A2(n_1302),
.B(n_1300),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1540),
.B(n_1364),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1616),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1413),
.B(n_760),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1448),
.B(n_764),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1497),
.B(n_765),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1464),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1430),
.B(n_767),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1621),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_L g1675 ( 
.A(n_1444),
.B(n_770),
.Y(n_1675)
);

BUFx12f_ASAP7_75t_L g1676 ( 
.A(n_1638),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1449),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1486),
.B(n_1469),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1603),
.A2(n_1222),
.B(n_1218),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1611),
.A2(n_1224),
.B(n_1222),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1472),
.B(n_773),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1499),
.Y(n_1682)
);

AO21x1_ASAP7_75t_L g1683 ( 
.A1(n_1546),
.A2(n_805),
.B(n_792),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1492),
.A2(n_1503),
.B(n_1531),
.C(n_1515),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1473),
.B(n_809),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1520),
.Y(n_1686)
);

AOI21xp33_ASAP7_75t_L g1687 ( 
.A1(n_1533),
.A2(n_815),
.B(n_811),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1601),
.A2(n_1228),
.B(n_1231),
.C(n_1227),
.Y(n_1688)
);

OAI321xp33_ASAP7_75t_L g1689 ( 
.A1(n_1495),
.A2(n_840),
.A3(n_834),
.B1(n_841),
.B2(n_839),
.C(n_817),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1457),
.B(n_845),
.Y(n_1690)
);

AO21x1_ASAP7_75t_L g1691 ( 
.A1(n_1648),
.A2(n_847),
.B(n_846),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1418),
.B(n_853),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1615),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1525),
.A2(n_1504),
.B(n_1460),
.C(n_1567),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1548),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1517),
.A2(n_1305),
.B(n_1304),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1424),
.A2(n_1550),
.B(n_1532),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_SL g1698 ( 
.A(n_1556),
.B(n_858),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1522),
.A2(n_866),
.B(n_863),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1456),
.B(n_868),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1507),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1551),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1459),
.A2(n_1509),
.B1(n_1521),
.B2(n_1535),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1523),
.A2(n_875),
.B(n_873),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1529),
.A2(n_892),
.B(n_884),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1478),
.B(n_899),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1476),
.B(n_1483),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1534),
.A2(n_912),
.B(n_907),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1542),
.A2(n_927),
.B(n_922),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1536),
.A2(n_932),
.B1(n_938),
.B2(n_931),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1547),
.A2(n_958),
.B1(n_964),
.B2(n_949),
.Y(n_1711)
);

OA22x2_ASAP7_75t_L g1712 ( 
.A1(n_1494),
.A2(n_1314),
.B1(n_1309),
.B2(n_990),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1508),
.B(n_1309),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1562),
.A2(n_1276),
.B(n_1152),
.Y(n_1714)
);

OAI321xp33_ASAP7_75t_L g1715 ( 
.A1(n_1412),
.A2(n_1471),
.A3(n_1574),
.B1(n_1501),
.B2(n_1564),
.C(n_1524),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1431),
.Y(n_1716)
);

CKINVDCx6p67_ASAP7_75t_R g1717 ( 
.A(n_1500),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1425),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1490),
.B(n_1364),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1445),
.B(n_1326),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1507),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1623),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1453),
.B(n_1330),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1414),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1625),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1636),
.Y(n_1726)
);

OR2x6_ASAP7_75t_L g1727 ( 
.A(n_1500),
.B(n_1410),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1420),
.Y(n_1728)
);

A2O1A1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1419),
.A2(n_1341),
.B(n_1347),
.C(n_1339),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1421),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1458),
.B(n_1341),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1461),
.B(n_1348),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1583),
.A2(n_1373),
.B(n_1358),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1423),
.A2(n_1373),
.B(n_1374),
.C(n_1358),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1639),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1491),
.B(n_1368),
.Y(n_1736)
);

INVx4_ASAP7_75t_L g1737 ( 
.A(n_1431),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1640),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1597),
.A2(n_1391),
.B(n_1389),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1465),
.B(n_1391),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1641),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1642),
.Y(n_1742)
);

BUFx8_ASAP7_75t_L g1743 ( 
.A(n_1627),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1431),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1443),
.A2(n_1399),
.B1(n_1401),
.B2(n_1394),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1466),
.B(n_1467),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1435),
.A2(n_1442),
.B(n_1441),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1607),
.A2(n_1405),
.B(n_1402),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1480),
.B(n_1370),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1454),
.B(n_1378),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1537),
.A2(n_1410),
.B1(n_1408),
.B2(n_1392),
.Y(n_1751)
);

NAND2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1447),
.B(n_1378),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1432),
.B(n_1392),
.Y(n_1753)
);

CKINVDCx10_ASAP7_75t_R g1754 ( 
.A(n_1627),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1646),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_SL g1756 ( 
.A1(n_1489),
.A2(n_1397),
.B(n_1395),
.C(n_46),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1608),
.A2(n_1397),
.B(n_1395),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1470),
.B(n_220),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1450),
.Y(n_1759)
);

AND2x6_ASAP7_75t_L g1760 ( 
.A(n_1598),
.B(n_225),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1451),
.Y(n_1761)
);

O2A1O1Ixp5_ASAP7_75t_L g1762 ( 
.A1(n_1569),
.A2(n_228),
.B(n_229),
.C(n_227),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1479),
.A2(n_232),
.B(n_231),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1609),
.A2(n_240),
.B(n_234),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1474),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1543),
.B(n_1589),
.Y(n_1766)
);

O2A1O1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1559),
.A2(n_46),
.B(n_43),
.C(n_44),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1455),
.B(n_43),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1422),
.A2(n_243),
.B1(n_248),
.B2(n_242),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1487),
.Y(n_1770)
);

BUFx12f_ASAP7_75t_L g1771 ( 
.A(n_1434),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1568),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1772)
);

BUFx4f_ASAP7_75t_L g1773 ( 
.A(n_1596),
.Y(n_1773)
);

BUFx12f_ASAP7_75t_L g1774 ( 
.A(n_1436),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1624),
.B(n_47),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1477),
.B(n_1481),
.Y(n_1776)
);

OR2x6_ASAP7_75t_SL g1777 ( 
.A(n_1527),
.B(n_49),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1571),
.B(n_51),
.C(n_52),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1484),
.A2(n_261),
.B(n_259),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1427),
.B(n_263),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1463),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1619),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1488),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1506),
.A2(n_271),
.B(n_267),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1619),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_R g1786 ( 
.A(n_1468),
.B(n_54),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1628),
.A2(n_277),
.B(n_276),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1656),
.A2(n_58),
.B(n_54),
.C(n_57),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1426),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1593),
.B(n_58),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1604),
.B(n_293),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1645),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1493),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1561),
.A2(n_65),
.B(n_61),
.C(n_63),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1545),
.B(n_63),
.Y(n_1795)
);

AOI22x1_ASAP7_75t_SL g1796 ( 
.A1(n_1617),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_SL g1797 ( 
.A1(n_1538),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1463),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1626),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1446),
.A2(n_298),
.B1(n_302),
.B2(n_296),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1514),
.B(n_71),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1510),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1463),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1541),
.A2(n_309),
.B1(n_312),
.B2(n_304),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1584),
.A2(n_316),
.B(n_315),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1530),
.B(n_321),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1539),
.B(n_327),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1511),
.B(n_72),
.Y(n_1808)
);

AOI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1610),
.A2(n_334),
.B(n_329),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_L g1810 ( 
.A(n_1462),
.B(n_72),
.C(n_73),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1588),
.B(n_339),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1614),
.A2(n_344),
.B(n_340),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1557),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1644),
.A2(n_354),
.B1(n_358),
.B2(n_352),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1573),
.B(n_359),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1557),
.Y(n_1816)
);

O2A1O1Ixp33_ASAP7_75t_L g1817 ( 
.A1(n_1654),
.A2(n_80),
.B(n_76),
.C(n_77),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1651),
.B(n_77),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1566),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1579),
.Y(n_1820)
);

BUFx12f_ASAP7_75t_L g1821 ( 
.A(n_1565),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1579),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1635),
.A2(n_364),
.B(n_363),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_SL g1824 ( 
.A1(n_1637),
.A2(n_83),
.B(n_80),
.C(n_81),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1570),
.Y(n_1825)
);

NOR2xp67_ASAP7_75t_L g1826 ( 
.A(n_1498),
.B(n_366),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1643),
.A2(n_368),
.B(n_367),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1557),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1575),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1496),
.A2(n_373),
.B1(n_374),
.B2(n_371),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1475),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1578),
.B(n_379),
.Y(n_1832)
);

CKINVDCx8_ASAP7_75t_R g1833 ( 
.A(n_1596),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1544),
.A2(n_383),
.B1(n_384),
.B2(n_381),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1554),
.A2(n_399),
.B1(n_400),
.B2(n_396),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1581),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1563),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1632),
.A2(n_1485),
.B(n_1528),
.C(n_1591),
.Y(n_1838)
);

AO31x2_ASAP7_75t_L g1839 ( 
.A1(n_1683),
.A2(n_1647),
.A3(n_1650),
.B(n_1618),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1684),
.B(n_1687),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1673),
.B(n_1585),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1678),
.A2(n_1595),
.B1(n_1513),
.B2(n_1587),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1661),
.A2(n_1599),
.B(n_1416),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1666),
.A2(n_1680),
.B(n_1679),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1657),
.A2(n_1560),
.B(n_1577),
.Y(n_1845)
);

O2A1O1Ixp5_ASAP7_75t_L g1846 ( 
.A1(n_1659),
.A2(n_1572),
.B(n_1505),
.C(n_1582),
.Y(n_1846)
);

AND2x6_ASAP7_75t_SL g1847 ( 
.A(n_1727),
.B(n_1502),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1682),
.Y(n_1848)
);

AND3x4_ASAP7_75t_L g1849 ( 
.A(n_1810),
.B(n_1592),
.C(n_1590),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1713),
.B(n_1475),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1747),
.A2(n_1613),
.B(n_1633),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1662),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1664),
.A2(n_1634),
.B1(n_1586),
.B2(n_1516),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1707),
.A2(n_1580),
.B(n_1653),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1686),
.Y(n_1855)
);

AO31x2_ASAP7_75t_L g1856 ( 
.A1(n_1665),
.A2(n_1606),
.A3(n_1612),
.B(n_1602),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1672),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1789),
.B(n_1439),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1780),
.A2(n_1429),
.B(n_1428),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1660),
.B(n_1552),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1668),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1694),
.A2(n_1622),
.B(n_1630),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1703),
.A2(n_1605),
.B(n_1652),
.Y(n_1863)
);

O2A1O1Ixp5_ASAP7_75t_L g1864 ( 
.A1(n_1692),
.A2(n_1690),
.B(n_1766),
.C(n_1669),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1695),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1677),
.B(n_1594),
.Y(n_1866)
);

OAI21x1_ASAP7_75t_L g1867 ( 
.A1(n_1696),
.A2(n_1555),
.B(n_1518),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1755),
.B(n_1652),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1674),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1722),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1681),
.A2(n_1629),
.B(n_1620),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1693),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1749),
.Y(n_1873)
);

AO31x2_ASAP7_75t_L g1874 ( 
.A1(n_1691),
.A2(n_1558),
.A3(n_90),
.B(n_87),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1685),
.A2(n_1558),
.B(n_1563),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1715),
.B(n_1440),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1801),
.B(n_1649),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1725),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1716),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1702),
.Y(n_1880)
);

AOI221x1_ASAP7_75t_L g1881 ( 
.A1(n_1763),
.A2(n_497),
.B1(n_402),
.B2(n_403),
.C(n_577),
.Y(n_1881)
);

OAI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1748),
.A2(n_404),
.B(n_401),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1701),
.B(n_1502),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1670),
.B(n_1549),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1718),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1663),
.A2(n_1655),
.B1(n_408),
.B2(n_412),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1700),
.A2(n_413),
.B(n_405),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1779),
.A2(n_423),
.B(n_415),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1768),
.B(n_1482),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1750),
.B(n_89),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1746),
.A2(n_426),
.B(n_425),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1775),
.B(n_89),
.Y(n_1893)
);

OAI21x1_ASAP7_75t_L g1894 ( 
.A1(n_1733),
.A2(n_428),
.B(n_427),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1776),
.A2(n_432),
.B(n_431),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1762),
.A2(n_1697),
.B(n_1724),
.Y(n_1896)
);

AOI21xp33_ASAP7_75t_L g1897 ( 
.A1(n_1808),
.A2(n_90),
.B(n_91),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1736),
.B(n_92),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1838),
.A2(n_92),
.B(n_93),
.C(n_95),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1716),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1671),
.B(n_95),
.Y(n_1901)
);

AO31x2_ASAP7_75t_L g1902 ( 
.A1(n_1729),
.A2(n_96),
.A3(n_97),
.B(n_98),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1728),
.B(n_96),
.Y(n_1903)
);

BUFx4f_ASAP7_75t_L g1904 ( 
.A(n_1717),
.Y(n_1904)
);

AO31x2_ASAP7_75t_L g1905 ( 
.A1(n_1745),
.A2(n_97),
.A3(n_98),
.B(n_99),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1806),
.A2(n_442),
.B(n_439),
.Y(n_1906)
);

OAI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1795),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1771),
.B(n_100),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1739),
.A2(n_1757),
.B(n_1807),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1730),
.B(n_101),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1716),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1811),
.A2(n_446),
.B(n_445),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1819),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1791),
.A2(n_448),
.B(n_447),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1726),
.B(n_102),
.Y(n_1915)
);

A2O1A1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1710),
.A2(n_103),
.B(n_104),
.C(n_106),
.Y(n_1916)
);

NAND2xp33_ASAP7_75t_L g1917 ( 
.A(n_1760),
.B(n_455),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1711),
.A2(n_576),
.B1(n_575),
.B2(n_574),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1744),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1758),
.A2(n_463),
.B(n_457),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1802),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1675),
.A2(n_465),
.B(n_464),
.Y(n_1922)
);

NOR2xp67_ASAP7_75t_SL g1923 ( 
.A(n_1689),
.B(n_103),
.Y(n_1923)
);

OAI21xp33_ASAP7_75t_L g1924 ( 
.A1(n_1790),
.A2(n_109),
.B(n_110),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1825),
.A2(n_477),
.B(n_474),
.Y(n_1925)
);

AO31x2_ASAP7_75t_L g1926 ( 
.A1(n_1799),
.A2(n_109),
.A3(n_111),
.B(n_112),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1809),
.A2(n_482),
.B(n_478),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1829),
.A2(n_492),
.B(n_488),
.Y(n_1928)
);

OR2x6_ASAP7_75t_L g1929 ( 
.A(n_1774),
.B(n_1727),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1836),
.A2(n_571),
.B1(n_569),
.B2(n_564),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1735),
.Y(n_1931)
);

AO21x1_ASAP7_75t_L g1932 ( 
.A1(n_1800),
.A2(n_113),
.B(n_115),
.Y(n_1932)
);

OAI21x1_ASAP7_75t_SL g1933 ( 
.A1(n_1805),
.A2(n_512),
.B(n_495),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1741),
.A2(n_516),
.B(n_513),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1738),
.Y(n_1935)
);

OA21x2_ASAP7_75t_L g1936 ( 
.A1(n_1699),
.A2(n_563),
.B(n_562),
.Y(n_1936)
);

AO31x2_ASAP7_75t_L g1937 ( 
.A1(n_1794),
.A2(n_115),
.A3(n_116),
.B(n_117),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1742),
.B(n_1759),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1761),
.B(n_116),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1765),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1770),
.B(n_120),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1783),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1831),
.A2(n_550),
.B1(n_548),
.B2(n_544),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1782),
.A2(n_542),
.B(n_541),
.Y(n_1944)
);

AOI21xp33_ASAP7_75t_L g1945 ( 
.A1(n_1818),
.A2(n_121),
.B(n_123),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1793),
.B(n_121),
.Y(n_1946)
);

OAI21x1_ASAP7_75t_L g1947 ( 
.A1(n_1785),
.A2(n_539),
.B(n_538),
.Y(n_1947)
);

NOR2x1_ASAP7_75t_SL g1948 ( 
.A(n_1744),
.B(n_522),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1720),
.Y(n_1949)
);

NOR4xp25_ASAP7_75t_L g1950 ( 
.A(n_1792),
.B(n_124),
.C(n_125),
.D(n_126),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1760),
.Y(n_1951)
);

NAND2x1p5_ASAP7_75t_L g1952 ( 
.A(n_1737),
.B(n_523),
.Y(n_1952)
);

OAI21x1_ASAP7_75t_L g1953 ( 
.A1(n_1714),
.A2(n_537),
.B(n_536),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1706),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1820),
.B(n_1822),
.Y(n_1955)
);

AO21x1_ASAP7_75t_L g1956 ( 
.A1(n_1767),
.A2(n_128),
.B(n_129),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1688),
.A2(n_532),
.B(n_531),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1815),
.B(n_1832),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1832),
.B(n_130),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1704),
.B(n_131),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1705),
.B(n_131),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1949),
.B(n_1760),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1850),
.B(n_1712),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1840),
.A2(n_1709),
.B(n_1708),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1869),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1841),
.A2(n_1760),
.B1(n_1778),
.B2(n_1719),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1913),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1860),
.B(n_1777),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1900),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1954),
.B(n_1877),
.Y(n_1970)
);

AND2x2_ASAP7_75t_SL g1971 ( 
.A(n_1917),
.B(n_1698),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1848),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_SL g1973 ( 
.A1(n_1842),
.A2(n_1796),
.B1(n_1753),
.B2(n_1821),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1958),
.B(n_1826),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1876),
.A2(n_1932),
.B1(n_1923),
.B2(n_1945),
.Y(n_1975)
);

A2O1A1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1889),
.A2(n_1864),
.B(n_1863),
.C(n_1862),
.Y(n_1976)
);

NAND2x1p5_ASAP7_75t_L g1977 ( 
.A(n_1900),
.B(n_1773),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1870),
.Y(n_1978)
);

OAI221xp5_ASAP7_75t_SL g1979 ( 
.A1(n_1890),
.A2(n_1817),
.B1(n_1788),
.B2(n_1772),
.C(n_1751),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1857),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1844),
.A2(n_1827),
.B(n_1823),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1868),
.A2(n_1951),
.B1(n_1959),
.B2(n_1865),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1921),
.B(n_1721),
.Y(n_1983)
);

AO32x2_ASAP7_75t_L g1984 ( 
.A1(n_1943),
.A2(n_1835),
.A3(n_1834),
.B1(n_1769),
.B2(n_1804),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1896),
.A2(n_1813),
.B(n_1744),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1855),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1866),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1904),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1880),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1885),
.B(n_1723),
.Y(n_1990)
);

OA21x2_ASAP7_75t_L g1991 ( 
.A1(n_1957),
.A2(n_1734),
.B(n_1740),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1878),
.Y(n_1992)
);

OAI21x1_ASAP7_75t_L g1993 ( 
.A1(n_1909),
.A2(n_1784),
.B(n_1812),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1931),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1858),
.B(n_1667),
.Y(n_1995)
);

NAND2x1_ASAP7_75t_SL g1996 ( 
.A(n_1898),
.B(n_1830),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1849),
.A2(n_1731),
.B1(n_1732),
.B2(n_1814),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1861),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1935),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1940),
.Y(n_2001)
);

OAI21x1_ASAP7_75t_L g2002 ( 
.A1(n_1859),
.A2(n_1787),
.B(n_1764),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1942),
.B(n_1752),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1891),
.B(n_1798),
.Y(n_2004)
);

CKINVDCx6p67_ASAP7_75t_R g2005 ( 
.A(n_1929),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1852),
.B(n_1803),
.Y(n_2006)
);

INVx4_ASAP7_75t_L g2007 ( 
.A(n_1919),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1872),
.B(n_1837),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1853),
.B(n_1901),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1938),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1893),
.B(n_1813),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1919),
.Y(n_2012)
);

BUFx10_ASAP7_75t_L g2013 ( 
.A(n_1883),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1955),
.Y(n_2014)
);

NAND2x1p5_ASAP7_75t_L g2015 ( 
.A(n_1911),
.B(n_1816),
.Y(n_2015)
);

OAI21x1_ASAP7_75t_L g2016 ( 
.A1(n_1944),
.A2(n_1828),
.B(n_1816),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1915),
.Y(n_2017)
);

O2A1O1Ixp33_ASAP7_75t_SL g2018 ( 
.A1(n_1899),
.A2(n_1756),
.B(n_1797),
.C(n_1824),
.Y(n_2018)
);

OR2x6_ASAP7_75t_L g2019 ( 
.A(n_1929),
.B(n_1676),
.Y(n_2019)
);

OAI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1903),
.A2(n_1828),
.B1(n_1816),
.B2(n_1781),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_L g2021 ( 
.A1(n_1947),
.A2(n_1828),
.B(n_524),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1910),
.B(n_132),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1939),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1941),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1851),
.A2(n_1786),
.B1(n_133),
.B2(n_134),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1843),
.A2(n_1884),
.B(n_1875),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1886),
.B(n_132),
.Y(n_2027)
);

NOR2xp67_ASAP7_75t_L g2028 ( 
.A(n_1854),
.B(n_134),
.Y(n_2028)
);

OAI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1927),
.A2(n_136),
.B(n_137),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1845),
.B(n_137),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1856),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1856),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1879),
.B(n_138),
.Y(n_2033)
);

OAI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1846),
.A2(n_138),
.B(n_140),
.Y(n_2034)
);

NOR2x1_ASAP7_75t_SL g2035 ( 
.A(n_1930),
.B(n_141),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1946),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1948),
.B(n_142),
.Y(n_2037)
);

AOI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1881),
.A2(n_142),
.B(n_143),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1937),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1925),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_2040)
);

OAI21x1_ASAP7_75t_L g2041 ( 
.A1(n_1882),
.A2(n_147),
.B(n_148),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1924),
.A2(n_1743),
.B1(n_149),
.B2(n_150),
.Y(n_2042)
);

BUFx12f_ASAP7_75t_L g2043 ( 
.A(n_1847),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1871),
.B(n_147),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1937),
.Y(n_2045)
);

OAI21x1_ASAP7_75t_L g2046 ( 
.A1(n_1894),
.A2(n_150),
.B(n_151),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1867),
.B(n_151),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1960),
.Y(n_2048)
);

AO31x2_ASAP7_75t_L g2049 ( 
.A1(n_1956),
.A2(n_154),
.A3(n_155),
.B(n_158),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1967),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1972),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1963),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2000),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1986),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1989),
.Y(n_2055)
);

BUFx12f_ASAP7_75t_L g2056 ( 
.A(n_2013),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1994),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_2033),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2001),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1980),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1965),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1978),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1992),
.Y(n_2063)
);

INVx4_ASAP7_75t_SL g2064 ( 
.A(n_2049),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_2006),
.B(n_1953),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1976),
.A2(n_1928),
.B(n_1888),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_SL g2067 ( 
.A1(n_1971),
.A2(n_1908),
.B1(n_1950),
.B2(n_1743),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_2009),
.B(n_1907),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2010),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_2040),
.A2(n_1897),
.B1(n_1961),
.B2(n_1918),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2048),
.B(n_2014),
.Y(n_2071)
);

AO21x1_ASAP7_75t_SL g2072 ( 
.A1(n_2034),
.A2(n_1933),
.B(n_1952),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_2033),
.Y(n_2073)
);

CKINVDCx6p67_ASAP7_75t_R g2074 ( 
.A(n_1988),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_2011),
.Y(n_2075)
);

BUFx3_ASAP7_75t_L g2076 ( 
.A(n_1999),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1990),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_2015),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2031),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2032),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2045),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2036),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2023),
.B(n_1839),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1970),
.B(n_1908),
.Y(n_2084)
);

INVx4_ASAP7_75t_SL g2085 ( 
.A(n_2049),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2039),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1969),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2004),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2013),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1969),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2017),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2029),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_2012),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2008),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2003),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2027),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2044),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2030),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2047),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2024),
.B(n_1968),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1995),
.B(n_1916),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1987),
.B(n_1887),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1962),
.B(n_1839),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2022),
.Y(n_2104)
);

OA21x2_ASAP7_75t_L g2105 ( 
.A1(n_1993),
.A2(n_1895),
.B(n_1892),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2028),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1964),
.A2(n_1920),
.B(n_1906),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2047),
.Y(n_2108)
);

CKINVDCx20_ASAP7_75t_R g2109 ( 
.A(n_2005),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_2012),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2049),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2038),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1974),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2038),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2042),
.B(n_1926),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1982),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_2007),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2037),
.Y(n_2118)
);

INVx3_ASAP7_75t_SL g2119 ( 
.A(n_2019),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2037),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1966),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_1977),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2058),
.B(n_2019),
.Y(n_2123)
);

INVx4_ASAP7_75t_L g2124 ( 
.A(n_2117),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_2091),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2077),
.B(n_1997),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2075),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2057),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2053),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2086),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2052),
.B(n_1973),
.Y(n_2131)
);

INVx4_ASAP7_75t_L g2132 ( 
.A(n_2117),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2075),
.B(n_1979),
.Y(n_2133)
);

BUFx2_ASAP7_75t_L g2134 ( 
.A(n_2060),
.Y(n_2134)
);

OR2x6_ASAP7_75t_L g2135 ( 
.A(n_2076),
.B(n_2043),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2052),
.B(n_2025),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2050),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2098),
.B(n_1983),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_2104),
.B(n_1975),
.Y(n_2139)
);

BUFx4f_ASAP7_75t_SL g2140 ( 
.A(n_2074),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2068),
.A2(n_1998),
.B1(n_2020),
.B2(n_1991),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2067),
.A2(n_1991),
.B1(n_1922),
.B2(n_1914),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_2073),
.B(n_2035),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2088),
.B(n_1926),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_2122),
.B(n_2035),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2101),
.B(n_2084),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2096),
.B(n_1905),
.Y(n_2147)
);

BUFx3_ASAP7_75t_L g2148 ( 
.A(n_2076),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2095),
.B(n_1905),
.Y(n_2149)
);

NOR2xp67_ASAP7_75t_L g2150 ( 
.A(n_2122),
.B(n_1985),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2094),
.B(n_1874),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_2090),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2113),
.B(n_1874),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2071),
.B(n_1996),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2071),
.B(n_1902),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_2118),
.B(n_2021),
.Y(n_2156)
);

INVx8_ASAP7_75t_L g2157 ( 
.A(n_2056),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_2087),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2100),
.B(n_1902),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2051),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2120),
.B(n_2016),
.Y(n_2161)
);

INVx5_ASAP7_75t_L g2162 ( 
.A(n_2117),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2079),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2080),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2082),
.B(n_2041),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_2090),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2081),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2112),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2061),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_2087),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2078),
.B(n_2046),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2069),
.B(n_1996),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2097),
.B(n_2018),
.Y(n_2173)
);

BUFx3_ASAP7_75t_L g2174 ( 
.A(n_2093),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2114),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_2109),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2063),
.Y(n_2177)
);

NAND2x1p5_ASAP7_75t_L g2178 ( 
.A(n_2078),
.B(n_2093),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2111),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_2110),
.Y(n_2180)
);

BUFx3_ASAP7_75t_L g2181 ( 
.A(n_2110),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2054),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2055),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_2108),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2059),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2062),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2067),
.B(n_1984),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2102),
.B(n_1984),
.Y(n_2188)
);

AOI21xp33_ASAP7_75t_L g2189 ( 
.A1(n_2070),
.A2(n_2026),
.B(n_2002),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2121),
.B(n_1912),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2102),
.B(n_1936),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2083),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2116),
.B(n_1934),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2115),
.B(n_155),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2099),
.B(n_160),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2127),
.B(n_2133),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2130),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2126),
.B(n_2106),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2168),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2139),
.B(n_2083),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2130),
.Y(n_2201)
);

BUFx2_ASAP7_75t_L g2202 ( 
.A(n_2134),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2168),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2175),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_2179),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_2161),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2179),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2146),
.B(n_2065),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2137),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_2148),
.Y(n_2210)
);

BUFx3_ASAP7_75t_L g2211 ( 
.A(n_2152),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2131),
.B(n_2103),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2187),
.B(n_2064),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2160),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_2192),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2183),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_2161),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_2166),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2182),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2185),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2194),
.B(n_2103),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2138),
.B(n_2119),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2195),
.B(n_2064),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_2143),
.B(n_2064),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_2143),
.B(n_2085),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2154),
.B(n_2070),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_2156),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2136),
.B(n_2085),
.Y(n_2228)
);

OR2x2_ASAP7_75t_L g2229 ( 
.A(n_2147),
.B(n_2119),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2144),
.B(n_2085),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2163),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2163),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2164),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2164),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2159),
.B(n_2089),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2149),
.B(n_2072),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2155),
.B(n_2092),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2167),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_2172),
.B(n_2066),
.Y(n_2239)
);

NOR2xp67_ASAP7_75t_L g2240 ( 
.A(n_2162),
.B(n_2124),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2162),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_2192),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2221),
.B(n_2212),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2207),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2199),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2197),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_2210),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2206),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2201),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2235),
.B(n_2188),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2236),
.B(n_2151),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2213),
.B(n_2191),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2213),
.B(n_2153),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2196),
.B(n_2158),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2237),
.B(n_2170),
.Y(n_2255)
);

AND2x4_ASAP7_75t_SL g2256 ( 
.A(n_2224),
.B(n_2145),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2205),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2226),
.B(n_2186),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2198),
.B(n_2200),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2205),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2239),
.B(n_2165),
.Y(n_2261)
);

NOR2xp67_ASAP7_75t_L g2262 ( 
.A(n_2222),
.B(n_2124),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2203),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_2215),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2228),
.B(n_2123),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2239),
.B(n_2128),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2204),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2215),
.Y(n_2268)
);

BUFx2_ASAP7_75t_L g2269 ( 
.A(n_2202),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2230),
.B(n_2167),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2242),
.Y(n_2271)
);

NOR2x1p5_ASAP7_75t_L g2272 ( 
.A(n_2229),
.B(n_2176),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2242),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2209),
.Y(n_2274)
);

AND2x2_ASAP7_75t_SL g2275 ( 
.A(n_2230),
.B(n_2142),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2248),
.B(n_2257),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2256),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2274),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2267),
.Y(n_2279)
);

NOR2x1_ASAP7_75t_SL g2280 ( 
.A(n_2268),
.B(n_2214),
.Y(n_2280)
);

OAI31xp33_ASAP7_75t_L g2281 ( 
.A1(n_2272),
.A2(n_2141),
.A3(n_2222),
.B(n_2145),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2267),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2250),
.B(n_2227),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2248),
.B(n_2206),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2260),
.B(n_2206),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2244),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2262),
.B(n_2208),
.Y(n_2287)
);

INVxp67_ASAP7_75t_L g2288 ( 
.A(n_2269),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_2256),
.Y(n_2289)
);

NAND3xp33_ASAP7_75t_SL g2290 ( 
.A(n_2247),
.B(n_2066),
.C(n_2109),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2246),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2249),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2259),
.B(n_2261),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2266),
.B(n_2211),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_L g2295 ( 
.A(n_2254),
.B(n_2211),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2261),
.B(n_2216),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2270),
.B(n_2217),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2245),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2263),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2243),
.B(n_2219),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_2264),
.B(n_2227),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2252),
.B(n_2227),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2264),
.B(n_2255),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2285),
.B(n_2270),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2279),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2297),
.B(n_2302),
.Y(n_2306)
);

INVx2_ASAP7_75t_SL g2307 ( 
.A(n_2303),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_2293),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2282),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_2296),
.Y(n_2310)
);

OAI221xp5_ASAP7_75t_L g2311 ( 
.A1(n_2281),
.A2(n_2258),
.B1(n_2135),
.B2(n_2218),
.C(n_2220),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2300),
.B(n_2252),
.Y(n_2312)
);

AOI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2290),
.A2(n_2275),
.B1(n_2224),
.B2(n_2225),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2286),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2294),
.A2(n_2275),
.B1(n_2224),
.B2(n_2225),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2288),
.B(n_2253),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2301),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2305),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2311),
.A2(n_2295),
.B1(n_2278),
.B2(n_2299),
.C(n_2292),
.Y(n_2319)
);

NOR3xp33_ASAP7_75t_L g2320 ( 
.A(n_2313),
.B(n_2287),
.C(n_2123),
.Y(n_2320)
);

A2O1A1Ixp33_ASAP7_75t_L g2321 ( 
.A1(n_2315),
.A2(n_2277),
.B(n_2289),
.C(n_2218),
.Y(n_2321)
);

OR2x2_ASAP7_75t_L g2322 ( 
.A(n_2307),
.B(n_2283),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2309),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2314),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2317),
.Y(n_2325)
);

AOI221xp5_ASAP7_75t_L g2326 ( 
.A1(n_2319),
.A2(n_2310),
.B1(n_2308),
.B2(n_2316),
.C(n_2312),
.Y(n_2326)
);

OAI211xp5_ASAP7_75t_L g2327 ( 
.A1(n_2321),
.A2(n_2291),
.B(n_2273),
.C(n_2271),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2320),
.A2(n_2304),
.B1(n_2297),
.B2(n_2225),
.Y(n_2328)
);

AOI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2325),
.A2(n_2304),
.B1(n_2253),
.B2(n_2251),
.Y(n_2329)
);

AOI211xp5_ASAP7_75t_SL g2330 ( 
.A1(n_2318),
.A2(n_2240),
.B(n_2289),
.C(n_2277),
.Y(n_2330)
);

INVxp67_ASAP7_75t_L g2331 ( 
.A(n_2324),
.Y(n_2331)
);

INVx5_ASAP7_75t_SL g2332 ( 
.A(n_2322),
.Y(n_2332)
);

NAND4xp25_ASAP7_75t_L g2333 ( 
.A(n_2323),
.B(n_2181),
.C(n_2174),
.D(n_2265),
.Y(n_2333)
);

AOI221xp5_ASAP7_75t_L g2334 ( 
.A1(n_2326),
.A2(n_2331),
.B1(n_2327),
.B2(n_2333),
.C(n_2328),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2332),
.B(n_2306),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2330),
.B(n_2276),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2329),
.A2(n_2135),
.B(n_2157),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2327),
.A2(n_2285),
.B1(n_2217),
.B2(n_2223),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2326),
.B(n_2280),
.Y(n_2339)
);

NOR3x1_ASAP7_75t_L g2340 ( 
.A(n_2327),
.B(n_2241),
.C(n_1754),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2335),
.B(n_2276),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2334),
.B(n_2298),
.Y(n_2342)
);

NAND3xp33_ASAP7_75t_L g2343 ( 
.A(n_2339),
.B(n_2162),
.C(n_2238),
.Y(n_2343)
);

OAI322xp33_ASAP7_75t_L g2344 ( 
.A1(n_2342),
.A2(n_2337),
.A3(n_2338),
.B1(n_2336),
.B2(n_2340),
.C1(n_2233),
.C2(n_2173),
.Y(n_2344)
);

NOR2x1_ASAP7_75t_L g2345 ( 
.A(n_2343),
.B(n_2341),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2342),
.B(n_2157),
.Y(n_2346)
);

NOR2xp67_ASAP7_75t_L g2347 ( 
.A(n_2343),
.B(n_161),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2347),
.Y(n_2348)
);

NAND4xp75_ASAP7_75t_L g2349 ( 
.A(n_2345),
.B(n_2241),
.C(n_2140),
.D(n_2150),
.Y(n_2349)
);

AOI31xp33_ASAP7_75t_L g2350 ( 
.A1(n_2346),
.A2(n_2178),
.A3(n_2132),
.B(n_2190),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2344),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2345),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2345),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_SL g2354 ( 
.A(n_2352),
.B(n_2193),
.C(n_2107),
.Y(n_2354)
);

AND2x2_ASAP7_75t_SL g2355 ( 
.A(n_2348),
.B(n_2132),
.Y(n_2355)
);

AO22x2_ASAP7_75t_L g2356 ( 
.A1(n_2353),
.A2(n_2125),
.B1(n_2284),
.B2(n_2129),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2351),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2349),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2350),
.B(n_2180),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2358),
.B(n_2357),
.Y(n_2360)
);

INVx2_ASAP7_75t_SL g2361 ( 
.A(n_2355),
.Y(n_2361)
);

OA22x2_ASAP7_75t_L g2362 ( 
.A1(n_2359),
.A2(n_2284),
.B1(n_2125),
.B2(n_2231),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_SL g2363 ( 
.A1(n_2354),
.A2(n_2180),
.B1(n_162),
.B2(n_163),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2356),
.B(n_2180),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2360),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2363),
.A2(n_2361),
.B(n_2364),
.Y(n_2366)
);

OA22x2_ASAP7_75t_L g2367 ( 
.A1(n_2362),
.A2(n_2169),
.B1(n_2177),
.B2(n_2184),
.Y(n_2367)
);

OA21x2_ASAP7_75t_L g2368 ( 
.A1(n_2360),
.A2(n_2107),
.B(n_1981),
.Y(n_2368)
);

AOI221xp5_ASAP7_75t_L g2369 ( 
.A1(n_2363),
.A2(n_2189),
.B1(n_162),
.B2(n_164),
.C(n_166),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_2363),
.A2(n_2156),
.B(n_2171),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2365),
.B(n_161),
.Y(n_2371)
);

AOI22xp33_ASAP7_75t_L g2372 ( 
.A1(n_2366),
.A2(n_2217),
.B1(n_2232),
.B2(n_2234),
.Y(n_2372)
);

AOI21xp33_ASAP7_75t_SL g2373 ( 
.A1(n_2367),
.A2(n_164),
.B(n_167),
.Y(n_2373)
);

OAI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2369),
.A2(n_2184),
.B(n_168),
.Y(n_2374)
);

XNOR2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2370),
.B(n_167),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2373),
.B(n_2368),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_SL g2377 ( 
.A1(n_2371),
.A2(n_2374),
.B1(n_2372),
.B2(n_2375),
.Y(n_2377)
);

AOI21xp5_ASAP7_75t_L g2378 ( 
.A1(n_2371),
.A2(n_2105),
.B(n_171),
.Y(n_2378)
);

OAI222xp33_ASAP7_75t_L g2379 ( 
.A1(n_2375),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.C1(n_173),
.C2(n_174),
.Y(n_2379)
);

OA21x2_ASAP7_75t_L g2380 ( 
.A1(n_2379),
.A2(n_172),
.B(n_173),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_SL g2381 ( 
.A1(n_2380),
.A2(n_2377),
.B1(n_2376),
.B2(n_2378),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2381),
.A2(n_2171),
.B1(n_2231),
.B2(n_2232),
.Y(n_2382)
);


endmodule