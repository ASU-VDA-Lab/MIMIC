module fake_jpeg_29225_n_345 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_28),
.Y(n_57)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_52),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_36),
.B1(n_34),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_68),
.B1(n_52),
.B2(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_69),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_20),
.B1(n_37),
.B2(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_44),
.B1(n_20),
.B2(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_36),
.B1(n_38),
.B2(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_43),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_76),
.B1(n_92),
.B2(n_106),
.Y(n_118)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_25),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_44),
.B1(n_51),
.B2(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_43),
.C(n_50),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_50),
.C(n_31),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_47),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_23),
.B1(n_20),
.B2(n_38),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_33),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_26),
.B1(n_31),
.B2(n_35),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_35),
.B(n_26),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_23),
.B1(n_20),
.B2(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_114),
.B(n_21),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_44),
.B1(n_49),
.B2(n_46),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_138),
.B1(n_71),
.B2(n_67),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_23),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_132),
.C(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_66),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_92),
.Y(n_146)
);

NOR2x1_ASAP7_75t_R g130 ( 
.A(n_95),
.B(n_22),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_80),
.B(n_22),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_32),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_32),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_123),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_76),
.A2(n_49),
.B1(n_45),
.B2(n_46),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_101),
.B1(n_90),
.B2(n_77),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_146),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_92),
.B(n_83),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_117),
.A3(n_140),
.B1(n_125),
.B2(n_136),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_155),
.B1(n_158),
.B2(n_140),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_154),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_127),
.C(n_130),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_153),
.C(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_159),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_78),
.B(n_94),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_151),
.A2(n_107),
.B(n_108),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_97),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_103),
.C(n_100),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_46),
.B1(n_45),
.B2(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_91),
.C(n_81),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_45),
.B1(n_46),
.B2(n_81),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_94),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_112),
.C(n_119),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_116),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_177),
.B1(n_182),
.B2(n_192),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_120),
.B1(n_110),
.B2(n_113),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_142),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_186),
.C(n_187),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_113),
.B1(n_126),
.B2(n_108),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_146),
.B1(n_154),
.B2(n_147),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_128),
.B1(n_135),
.B2(n_139),
.Y(n_222)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_107),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_162),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_191),
.B(n_122),
.Y(n_218)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_125),
.B1(n_45),
.B2(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_200),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_162),
.B1(n_150),
.B2(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_190),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_109),
.B1(n_135),
.B2(n_117),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_213),
.B1(n_88),
.B2(n_79),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_162),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_192),
.B1(n_172),
.B2(n_171),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_216),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_24),
.B1(n_38),
.B2(n_27),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_176),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_217)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_224),
.B(n_71),
.Y(n_244)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_136),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_186),
.B1(n_99),
.B2(n_86),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_183),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_225),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_170),
.A2(n_128),
.B1(n_139),
.B2(n_122),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_21),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_227),
.A2(n_238),
.B1(n_239),
.B2(n_245),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_170),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_234),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_244),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_219),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_190),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_180),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_222),
.B1(n_205),
.B2(n_204),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_74),
.C(n_71),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_246),
.C(n_250),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_41),
.C(n_40),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_28),
.B(n_25),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_218),
.C(n_208),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_208),
.B1(n_206),
.B2(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_227),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_262),
.B1(n_263),
.B2(n_0),
.Y(n_284)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_199),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_269),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_250),
.A2(n_205),
.B1(n_204),
.B2(n_203),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_203),
.C(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_264),
.C(n_241),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_206),
.C(n_200),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_226),
.B(n_245),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_220),
.B1(n_210),
.B2(n_39),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_210),
.B1(n_37),
.B2(n_12),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_210),
.C(n_37),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_8),
.B(n_9),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_243),
.B(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_7),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_8),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_19),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_19),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_248),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_287),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_281),
.B1(n_270),
.B2(n_285),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_286),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_238),
.C(n_239),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_283),
.C(n_251),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_25),
.B(n_8),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_279),
.B(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_7),
.C(n_16),
.Y(n_283)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_259),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_17),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_260),
.B(n_17),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_13),
.Y(n_299)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_265),
.B1(n_270),
.B2(n_263),
.C(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_295),
.A2(n_6),
.B(n_1),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_288),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_9),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_1),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_251),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_280),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_253),
.C(n_264),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_283),
.C(n_255),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_278),
.B1(n_255),
.B2(n_286),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_309),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_287),
.B(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_312),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_316),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_275),
.B1(n_262),
.B2(n_256),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_9),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_0),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_302),
.C(n_298),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_2),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_296),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_5),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_301),
.B(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

AO221x1_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_303),
.B1(n_294),
.B2(n_316),
.C(n_317),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_1),
.B(n_2),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_304),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_327),
.A2(n_331),
.B(n_333),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_330),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_2),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_334),
.B(n_4),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_3),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_4),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_322),
.B1(n_324),
.B2(n_323),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_336),
.B(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_4),
.C(n_5),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_338),
.B(n_337),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_340),
.C(n_5),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_5),
.Y(n_345)
);


endmodule