module fake_jpeg_5163_n_71 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_4),
.B1(n_21),
.B2(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_6),
.B(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_3),
.C(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_18),
.B(n_0),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_0),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_52),
.C(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_49),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_10),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_29),
.A2(n_34),
.B1(n_38),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_30),
.B1(n_43),
.B2(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_45),
.B1(n_37),
.B2(n_25),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_56),
.B1(n_54),
.B2(n_46),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_40),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_23),
.B1(n_36),
.B2(n_24),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.C(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_49),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_56),
.B1(n_55),
.B2(n_50),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.C(n_68),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_68),
.B(n_61),
.C(n_60),
.Y(n_71)
);


endmodule