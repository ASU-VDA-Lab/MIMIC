module fake_jpeg_2617_n_559 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_559);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_559;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_6),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_78),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_64),
.Y(n_139)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_118),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_70),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_0),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_71),
.B(n_110),
.Y(n_158)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_72),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_0),
.C(n_1),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_114),
.C(n_35),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_13),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_35),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_88),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

CKINVDCx6p67_ASAP7_75t_R g190 ( 
.A(n_91),
.Y(n_190)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_104),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_33),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_117),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_44),
.B(n_2),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_35),
.B(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_19),
.B(n_3),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_119),
.B(n_121),
.Y(n_191)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_57),
.Y(n_138)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_26),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_122),
.B(n_106),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_126),
.Y(n_200)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_129),
.B(n_161),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_138),
.B(n_163),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_35),
.B(n_25),
.C(n_53),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_141),
.A2(n_173),
.B(n_170),
.C(n_152),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_71),
.A2(n_24),
.B1(n_32),
.B2(n_53),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_145),
.A2(n_155),
.B1(n_169),
.B2(n_175),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_64),
.A2(n_29),
.B1(n_51),
.B2(n_49),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_146),
.A2(n_157),
.B1(n_167),
.B2(n_181),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_60),
.A2(n_24),
.B1(n_32),
.B2(n_25),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_30),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_156),
.B(n_160),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_97),
.A2(n_31),
.B1(n_51),
.B2(n_49),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_30),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_57),
.C(n_55),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_69),
.B(n_19),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_48),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_164),
.B(n_166),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_68),
.B(n_48),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_76),
.A2(n_31),
.B1(n_29),
.B2(n_51),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_84),
.A2(n_28),
.B1(n_55),
.B2(n_45),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_45),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_172),
.B(n_178),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_58),
.A2(n_29),
.B1(n_49),
.B2(n_34),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_89),
.A2(n_34),
.B1(n_31),
.B2(n_42),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_184),
.B1(n_82),
.B2(n_79),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_92),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_34),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_179),
.B(n_195),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_113),
.A2(n_95),
.B1(n_91),
.B2(n_42),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_7),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_3),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_7),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_196),
.A2(n_211),
.B(n_13),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_59),
.A2(n_42),
.B1(n_56),
.B2(n_46),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_197),
.A2(n_198),
.B1(n_154),
.B2(n_170),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_100),
.A2(n_42),
.B1(n_36),
.B2(n_46),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_101),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_74),
.B(n_7),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_62),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_213),
.B(n_215),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_214),
.A2(n_234),
.B1(n_237),
.B2(n_263),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_63),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_216),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_142),
.A2(n_56),
.B1(n_67),
.B2(n_116),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_217),
.Y(n_323)
);

OA22x2_ASAP7_75t_SL g218 ( 
.A1(n_158),
.A2(n_83),
.B1(n_56),
.B2(n_42),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_218),
.A2(n_275),
.B(n_185),
.C(n_152),
.Y(n_316)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_139),
.Y(n_221)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_227),
.Y(n_288)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_132),
.A2(n_177),
.B1(n_127),
.B2(n_182),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_231),
.Y(n_328)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_42),
.B1(n_36),
.B2(n_43),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_240),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_36),
.B1(n_43),
.B2(n_11),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_245),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_241),
.B(n_242),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_43),
.B1(n_9),
.B2(n_11),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_243),
.A2(n_247),
.B1(n_256),
.B2(n_262),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_194),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_244),
.B(n_248),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_149),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_252),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_188),
.A2(n_43),
.B1(n_9),
.B2(n_12),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_173),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_165),
.Y(n_249)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_250),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_141),
.B(n_8),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_271),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_127),
.B(n_8),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_130),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_258),
.B(n_269),
.Y(n_337)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_157),
.A2(n_146),
.B(n_167),
.C(n_144),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_281),
.B(n_162),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_212),
.A2(n_201),
.B1(n_168),
.B2(n_137),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_131),
.A2(n_143),
.B1(n_182),
.B2(n_134),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_165),
.A2(n_187),
.B1(n_207),
.B2(n_168),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_264),
.A2(n_252),
.B1(n_239),
.B2(n_218),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_265),
.A2(n_278),
.B1(n_136),
.B2(n_153),
.Y(n_314)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_136),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_140),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_276),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_134),
.A2(n_193),
.B1(n_174),
.B2(n_135),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_277),
.A2(n_284),
.B1(n_185),
.B2(n_159),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_128),
.A2(n_162),
.B1(n_189),
.B2(n_147),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_173),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_282),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_137),
.A2(n_192),
.B(n_187),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_135),
.A2(n_193),
.B1(n_174),
.B2(n_148),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_128),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_133),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_233),
.B(n_154),
.C(n_159),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_293),
.B(n_271),
.C(n_276),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_302),
.B(n_322),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_238),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_303),
.B(n_309),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_222),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_223),
.A2(n_189),
.B1(n_147),
.B2(n_148),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_310),
.A2(n_340),
.B1(n_278),
.B2(n_240),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_339),
.B1(n_253),
.B2(n_250),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_335),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_215),
.B(n_153),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_318),
.B(n_319),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_213),
.B(n_180),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_245),
.B1(n_246),
.B2(n_249),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_233),
.B(n_159),
.CI(n_133),
.CON(n_321),
.SN(n_321)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_321),
.Y(n_348)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_283),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_327),
.B(n_279),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_236),
.B(n_226),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_266),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_228),
.A2(n_255),
.B1(n_214),
.B2(n_236),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_260),
.A2(n_251),
.B1(n_218),
.B2(n_233),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_261),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_342),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_267),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_302),
.A2(n_275),
.B(n_224),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_316),
.A2(n_281),
.B(n_273),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_345),
.A2(n_349),
.B(n_343),
.Y(n_400)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_296),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_371),
.Y(n_385)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_365),
.Y(n_415)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_355),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_356),
.A2(n_359),
.B1(n_364),
.B2(n_373),
.Y(n_394)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_360),
.B(n_367),
.Y(n_396)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_305),
.Y(n_361)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_247),
.B1(n_273),
.B2(n_256),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_308),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_R g366 ( 
.A(n_289),
.B(n_253),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_380),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_333),
.B(n_229),
.Y(n_367)
);

AO22x1_ASAP7_75t_SL g368 ( 
.A1(n_340),
.A2(n_273),
.B1(n_225),
.B2(n_219),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_370),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_286),
.A2(n_273),
.B1(n_270),
.B2(n_268),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_369),
.A2(n_376),
.B1(n_323),
.B2(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_290),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_290),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_372),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_286),
.A2(n_272),
.B1(n_285),
.B2(n_230),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_288),
.B(n_235),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_379),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_318),
.Y(n_391)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_378),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_297),
.B(n_232),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_254),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_298),
.B(n_257),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_293),
.C(n_336),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_297),
.A2(n_282),
.B1(n_220),
.B2(n_221),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_382),
.A2(n_314),
.B1(n_291),
.B2(n_329),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_400),
.B(n_376),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_397),
.Y(n_417)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_348),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_393),
.Y(n_420)
);

AO22x1_ASAP7_75t_L g397 ( 
.A1(n_349),
.A2(n_291),
.B1(n_310),
.B2(n_328),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_319),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_405),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_407),
.C(n_416),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_375),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_307),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_351),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_411),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_317),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_307),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_357),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_349),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_416),
.B(n_368),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_423),
.C(n_436),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_385),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_422),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_389),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_368),
.C(n_380),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_387),
.A2(n_345),
.B1(n_364),
.B2(n_354),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_424),
.A2(n_425),
.B1(n_431),
.B2(n_446),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_376),
.B1(n_369),
.B2(n_335),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_426),
.A2(n_427),
.B(n_439),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_400),
.A2(n_376),
.B(n_328),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_404),
.A2(n_323),
.B1(n_380),
.B2(n_366),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_436),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_415),
.A2(n_304),
.B1(n_355),
.B2(n_346),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_442),
.Y(n_455)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_306),
.Y(n_435)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_321),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_388),
.A2(n_304),
.B1(n_382),
.B2(n_352),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_394),
.B1(n_397),
.B2(n_398),
.Y(n_447)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_404),
.A2(n_324),
.B(n_300),
.Y(n_439)
);

OAI21xp33_ASAP7_75t_L g440 ( 
.A1(n_410),
.A2(n_321),
.B(n_298),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_440),
.B(n_443),
.Y(n_450)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_415),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_410),
.A2(n_317),
.B(n_350),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_389),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_399),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_363),
.B1(n_358),
.B2(n_361),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_447),
.A2(n_458),
.B1(n_422),
.B2(n_444),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_407),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_454),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_456),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_445),
.A2(n_397),
.B1(n_405),
.B2(n_391),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_414),
.C(n_413),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_462),
.C(n_463),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_414),
.C(n_413),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_408),
.C(n_395),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_396),
.B1(n_386),
.B2(n_408),
.Y(n_464)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_435),
.B(n_396),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_465),
.B(n_421),
.Y(n_490)
);

AO21x1_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_470),
.B(n_441),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_433),
.A2(n_395),
.B1(n_392),
.B2(n_402),
.Y(n_468)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_468),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_419),
.B(n_392),
.C(n_402),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_439),
.C(n_417),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_424),
.A2(n_383),
.B1(n_403),
.B2(n_365),
.Y(n_470)
);

OAI22x1_ASAP7_75t_SL g472 ( 
.A1(n_425),
.A2(n_383),
.B1(n_377),
.B2(n_370),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_446),
.B1(n_442),
.B2(n_445),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_298),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_443),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_475),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_476),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_467),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_479),
.A2(n_458),
.B1(n_447),
.B2(n_472),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_483),
.Y(n_497)
);

MAJx2_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_426),
.C(n_430),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_462),
.C(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_460),
.C(n_463),
.Y(n_498)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_487),
.Y(n_504)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_452),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_454),
.B(n_429),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_491),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_427),
.B(n_431),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_489),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_492),
.Y(n_506)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_457),
.A2(n_437),
.B1(n_430),
.B2(n_432),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_455),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_502),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_499),
.B(n_505),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_480),
.C(n_477),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_508),
.C(n_510),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_501),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_479),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_486),
.A2(n_467),
.B1(n_450),
.B2(n_466),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_507),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_470),
.C(n_473),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_482),
.A2(n_453),
.B(n_471),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_509),
.A2(n_491),
.B(n_476),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_449),
.Y(n_510)
);

OAI322xp33_ASAP7_75t_L g513 ( 
.A1(n_506),
.A2(n_474),
.A3(n_483),
.B1(n_485),
.B2(n_495),
.C1(n_488),
.C2(n_481),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_513),
.A2(n_497),
.B(n_499),
.Y(n_526)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_504),
.Y(n_514)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_516),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_489),
.C(n_478),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_503),
.C(n_508),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_517),
.Y(n_534)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_521),
.Y(n_525)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_494),
.C(n_428),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_524),
.C(n_511),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_526),
.A2(n_530),
.B(n_531),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_519),
.A2(n_507),
.B1(n_511),
.B2(n_505),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_529),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_523),
.A2(n_497),
.B(n_448),
.Y(n_530)
);

XOR2x2_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_459),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_523),
.A2(n_520),
.B1(n_522),
.B2(n_519),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_524),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_517),
.A2(n_438),
.B(n_434),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_315),
.B(n_338),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_537),
.A2(n_542),
.B1(n_543),
.B2(n_544),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_512),
.C(n_371),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_540),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_512),
.C(n_353),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_372),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_541),
.B(n_531),
.Y(n_546)
);

OAI221xp5_ASAP7_75t_L g542 ( 
.A1(n_525),
.A2(n_315),
.B1(n_329),
.B2(n_334),
.C(n_338),
.Y(n_542)
);

AOI322xp5_ASAP7_75t_L g544 ( 
.A1(n_530),
.A2(n_372),
.A3(n_332),
.B1(n_420),
.B2(n_326),
.C1(n_312),
.C2(n_334),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_546),
.B(n_550),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_529),
.Y(n_548)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_548),
.A2(n_331),
.B(n_292),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_538),
.A2(n_528),
.B(n_311),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_549),
.A2(n_311),
.B1(n_274),
.B2(n_259),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_536),
.B(n_332),
.C(n_331),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_551),
.A2(n_553),
.B(n_554),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_548),
.A2(n_301),
.B(n_295),
.Y(n_554)
);

AOI321xp33_ASAP7_75t_L g556 ( 
.A1(n_552),
.A2(n_547),
.A3(n_545),
.B1(n_550),
.B2(n_295),
.C(n_301),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_292),
.C(n_216),
.Y(n_557)
);

AO21x1_ASAP7_75t_L g558 ( 
.A1(n_557),
.A2(n_555),
.B(n_326),
.Y(n_558)
);

BUFx24_ASAP7_75t_SL g559 ( 
.A(n_558),
.Y(n_559)
);


endmodule