module fake_jpeg_1891_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_0),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_55),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_51),
.B1(n_56),
.B2(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_56),
.B1(n_55),
.B2(n_57),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_69),
.B1(n_70),
.B2(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_47),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_52),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_72),
.B1(n_58),
.B2(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_73),
.B1(n_72),
.B2(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_47),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_71),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_53),
.B(n_64),
.Y(n_123)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_68),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_49),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_52),
.C(n_50),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_112),
.C(n_3),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_65),
.B1(n_70),
.B2(n_60),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_119),
.B(n_8),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_29),
.B1(n_39),
.B2(n_38),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_63),
.C(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_76),
.B(n_66),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_96),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_24),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_100),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_126),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_105),
.B1(n_108),
.B2(n_117),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_23),
.B1(n_44),
.B2(n_41),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_133),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_140),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_27),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_116),
.C(n_110),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_10),
.B(n_11),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_11),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_25),
.B1(n_37),
.B2(n_35),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_46),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_154),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_112),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_131),
.C(n_28),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_12),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_127),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_161),
.B1(n_143),
.B2(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_167),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_170),
.B1(n_150),
.B2(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_154),
.C(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_176),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_159),
.B1(n_156),
.B2(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_166),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_171),
.C(n_169),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_148),
.Y(n_183)
);

NAND4xp25_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.C(n_178),
.D(n_147),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_178),
.B(n_177),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_170),
.C(n_150),
.Y(n_187)
);

NAND4xp25_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_181),
.C(n_161),
.D(n_180),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_179),
.C(n_31),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_33),
.C(n_15),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_16),
.Y(n_191)
);


endmodule