module real_jpeg_31485_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_366;
wire n_149;
wire n_332;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_653;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_0),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_1),
.A2(n_358),
.B1(n_359),
.B2(n_362),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_1),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_1),
.A2(n_358),
.B1(n_422),
.B2(n_427),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_1),
.A2(n_358),
.B1(n_547),
.B2(n_550),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_1),
.A2(n_358),
.B1(n_587),
.B2(n_593),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_3),
.A2(n_153),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_3),
.A2(n_269),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_3),
.A2(n_190),
.B1(n_269),
.B2(n_526),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_3),
.A2(n_269),
.B1(n_568),
.B2(n_573),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_61),
.B1(n_110),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_61),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_5),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_5),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_5),
.A2(n_199),
.B1(n_240),
.B2(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_5),
.A2(n_240),
.B1(n_408),
.B2(n_410),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_5),
.A2(n_240),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_6),
.B(n_347),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_6),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_6),
.B(n_146),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g499 ( 
.A1(n_6),
.A2(n_500),
.A3(n_502),
.B1(n_506),
.B2(n_512),
.Y(n_499)
);

OAI32xp33_ASAP7_75t_L g544 ( 
.A1(n_6),
.A2(n_500),
.A3(n_502),
.B1(n_506),
.B2(n_512),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_6),
.A2(n_419),
.B1(n_553),
.B2(n_554),
.Y(n_552)
);

OAI21xp33_ASAP7_75t_L g632 ( 
.A1(n_6),
.A2(n_209),
.B(n_578),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_7),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_7),
.A2(n_115),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_7),
.A2(n_115),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_7),
.A2(n_115),
.B1(n_444),
.B2(n_448),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_8),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_8),
.A2(n_151),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_8),
.A2(n_151),
.B1(n_295),
.B2(n_300),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_8),
.A2(n_151),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_11),
.Y(n_286)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_11),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_14),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_14),
.B(n_251),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_15),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_15),
.A2(n_109),
.B1(n_190),
.B2(n_194),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_15),
.A2(n_109),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_16),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_17),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_18),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_18),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_18),
.A2(n_101),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_18),
.A2(n_101),
.B1(n_226),
.B2(n_229),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_18),
.A2(n_101),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_253),
.B(n_655),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_250),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_21),
.B(n_251),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_246),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_180),
.C(n_244),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_24),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_159),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_65),
.C(n_112),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_27),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_27),
.A2(n_65),
.B1(n_66),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_27),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_44),
.B(n_59),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_28),
.A2(n_44),
.B1(n_59),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_28),
.A2(n_44),
.B1(n_407),
.B2(n_412),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_28),
.B(n_407),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_28),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

OAI22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_37),
.B2(n_41),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_36),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_36),
.Y(n_290)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_36),
.Y(n_323)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_36),
.Y(n_336)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_36),
.Y(n_447)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_37),
.Y(n_611)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_40),
.Y(n_220)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_40),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_42),
.Y(n_603)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_43),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_44),
.B(n_622),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_45),
.A2(n_189),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_45),
.A2(n_224),
.B1(n_225),
.B2(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_45),
.A2(n_224),
.B1(n_294),
.B2(n_383),
.Y(n_382)
);

OAI21xp33_ASAP7_75t_SL g524 ( 
.A1(n_45),
.A2(n_525),
.B(n_529),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_45),
.A2(n_224),
.B1(n_525),
.B2(n_546),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_45),
.A2(n_546),
.B1(n_562),
.B2(n_563),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_49),
.Y(n_517)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_56),
.Y(n_409)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_58),
.Y(n_196)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_58),
.Y(n_299)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_64),
.Y(n_228)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_95),
.B1(n_105),
.B2(n_107),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_67),
.A2(n_105),
.B1(n_421),
.B2(n_430),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_68),
.A2(n_105),
.B1(n_107),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_68),
.A2(n_95),
.B1(n_105),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_68),
.A2(n_106),
.B1(n_198),
.B2(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_68),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_68),
.B(n_372),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_82),
.Y(n_68)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_76),
.B2(n_80),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_74),
.Y(n_302)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_75),
.Y(n_505)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_79),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_90),
.B2(n_93),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_85),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_125),
.B1(n_128),
.B2(n_131),
.Y(n_124)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_94),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_100),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_100),
.Y(n_426)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_104),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_106),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_106),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_111),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_183),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_122),
.B1(n_145),
.B2(n_147),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_114),
.B(n_146),
.Y(n_243)
);

BUFx4f_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_123),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_123),
.B(n_268),
.Y(n_267)
);

AO22x1_ASAP7_75t_L g394 ( 
.A1(n_123),
.A2(n_146),
.B1(n_268),
.B2(n_357),
.Y(n_394)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_123),
.A2(n_346),
.B(n_415),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_135),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_128),
.Y(n_341)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_130),
.Y(n_354)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2x1_ASAP7_75t_SL g266 ( 
.A(n_146),
.B(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_146),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_149),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_150),
.Y(n_345)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_156),
.Y(n_347)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_158),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_167),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_179),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_175),
.Y(n_361)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_245),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B(n_206),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_182),
.B(n_185),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_182),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_186),
.A2(n_187),
.B(n_197),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_186),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_192),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_196),
.Y(n_384)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_206),
.B(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_222),
.B(n_233),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_207),
.A2(n_208),
.B1(n_233),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_207),
.A2(n_208),
.B1(n_223),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_216),
.B(n_218),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_209),
.A2(n_218),
.B1(n_283),
.B2(n_291),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_209),
.A2(n_283),
.B1(n_378),
.B2(n_381),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_209),
.A2(n_316),
.B1(n_443),
.B2(n_449),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_209),
.A2(n_567),
.B(n_578),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_210),
.A2(n_315),
.B1(n_324),
.B2(n_330),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_210),
.B(n_520),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_210),
.A2(n_585),
.B1(n_596),
.B2(n_598),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_212),
.Y(n_332)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_216),
.A2(n_443),
.B(n_519),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_216),
.A2(n_519),
.B(n_586),
.Y(n_630)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_223),
.Y(n_477)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_232),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_232),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_232),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_232),
.Y(n_616)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_243),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_234),
.B(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_253),
.A2(n_656),
.B(n_657),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_306),
.B(n_653),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_303),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_256),
.B(n_303),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_257),
.B(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_261),
.B(n_263),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_272),
.C(n_281),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_265),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_265),
.B(n_275),
.Y(n_470)
);

NAND2x1_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_266),
.B(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_273),
.A2(n_468),
.B(n_470),
.Y(n_467)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_276),
.Y(n_392)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_279),
.Y(n_373)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_281),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_293),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_282),
.Y(n_396)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_286),
.Y(n_572)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_290),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_293),
.Y(n_397)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_299),
.Y(n_609)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_489),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_458),
.B(n_483),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_398),
.C(n_431),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_310),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_374),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_311),
.B(n_375),
.C(n_395),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_355),
.C(n_363),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_313),
.B(n_401),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_337),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_314),
.B(n_337),
.Y(n_435)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_322),
.Y(n_448)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_324),
.B(n_520),
.Y(n_578)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_329),
.Y(n_451)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_332),
.Y(n_522)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_335),
.Y(n_521)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI32xp33_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_341),
.A3(n_342),
.B1(n_346),
.B2(n_348),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_SL g351 ( 
.A(n_340),
.Y(n_351)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_351),
.Y(n_507)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_363),
.Y(n_401)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_365),
.B(n_371),
.Y(n_363)
);

OAI22x1_ASAP7_75t_L g390 ( 
.A1(n_364),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_364),
.A2(n_371),
.B(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_365),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_395),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_389),
.Y(n_375)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_382),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_382),
.Y(n_403)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_383),
.Y(n_412)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_393),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_393),
.B(n_419),
.Y(n_565)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_394),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_398),
.Y(n_492)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.C(n_404),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_399),
.A2(n_400),
.B1(n_455),
.B2(n_457),
.Y(n_454)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_402),
.A2(n_403),
.B1(n_405),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_405),
.Y(n_456)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.C(n_420),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_420),
.Y(n_434)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_407),
.Y(n_563)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_419),
.B(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_419),
.B(n_606),
.Y(n_605)
);

OAI21xp33_ASAP7_75t_SL g622 ( 
.A1(n_419),
.A2(n_605),
.B(n_623),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_419),
.B(n_562),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_419),
.B(n_635),
.Y(n_634)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_454),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_432),
.B(n_454),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_436),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_433),
.B(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_435),
.B(n_437),
.Y(n_535)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_442),
.C(n_452),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_438),
.B(n_532),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_440),
.B(n_441),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_442),
.A2(n_452),
.B1(n_453),
.B2(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_442),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx12f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_455),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_491),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_460),
.A2(n_463),
.B(n_478),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_463),
.Y(n_488)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_464),
.Y(n_487)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_472),
.C(n_476),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2x1_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_481),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.C(n_475),
.Y(n_472)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_476),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_479),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_482),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_484),
.A2(n_487),
.B(n_488),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_494),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_536),
.B(n_651),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_534),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_497),
.B(n_652),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_523),
.C(n_530),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_498),
.A2(n_523),
.B1(n_524),
.B2(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_498),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_518),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_501),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_516),
.Y(n_625)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_527),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_529),
.B(n_621),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_534),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_579),
.B(n_650),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_557),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_542),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_539),
.B(n_542),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_545),
.C(n_551),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_559),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_551),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_548),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_560),
.Y(n_557)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_558),
.Y(n_648)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_564),
.C(n_566),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_561),
.B(n_565),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_566),
.B(n_643),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_569),
.B(n_602),
.Y(n_601)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_572),
.Y(n_577)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_646),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_641),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_582),
.A2(n_626),
.B(n_640),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_599),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_584),
.B(n_599),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_597),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_620),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_600),
.B(n_620),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_601),
.A2(n_604),
.B1(n_610),
.B2(n_612),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_603),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_617),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_628),
.A2(n_631),
.B(n_639),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_629),
.B(n_630),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_629),
.B(n_630),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_632),
.B(n_633),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_634),
.B(n_636),
.Y(n_633)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_642),
.B(n_644),
.Y(n_641)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_642),
.Y(n_649)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_647),
.B1(n_648),
.B2(n_649),
.Y(n_646)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);


endmodule