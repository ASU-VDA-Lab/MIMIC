module fake_jpeg_6968_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_21),
.B1(n_33),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_55),
.B1(n_61),
.B2(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_21),
.B1(n_29),
.B2(n_37),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_31),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_65),
.Y(n_94)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_33),
.B1(n_20),
.B2(n_30),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_30),
.B1(n_17),
.B2(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_74),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_42),
.C(n_39),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_89),
.C(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_77),
.B1(n_85),
.B2(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_45),
.B1(n_50),
.B2(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_42),
.B1(n_39),
.B2(n_37),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_22),
.B1(n_35),
.B2(n_18),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_35),
.C(n_18),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_45),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_22),
.B1(n_35),
.B2(n_18),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_53),
.B1(n_51),
.B2(n_27),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_66),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_35),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_35),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_108),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_53),
.Y(n_108)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_85),
.B1(n_92),
.B2(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_116),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_84),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_53),
.B1(n_51),
.B2(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_86),
.B1(n_72),
.B2(n_70),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_51),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_74),
.B(n_82),
.C(n_75),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_118),
.B(n_86),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_19),
.B(n_18),
.C(n_32),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_126),
.B(n_128),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_132),
.B1(n_134),
.B2(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_137),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_117),
.B1(n_79),
.B2(n_115),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_77),
.B1(n_71),
.B2(n_68),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_106),
.B(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_149),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_89),
.B1(n_69),
.B2(n_73),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_72),
.B1(n_70),
.B2(n_83),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_146),
.B(n_148),
.Y(n_168)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_90),
.C(n_13),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_114),
.B1(n_111),
.B2(n_109),
.C(n_13),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_18),
.B(n_19),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_11),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_19),
.B(n_34),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_70),
.B1(n_72),
.B2(n_64),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_120),
.B1(n_109),
.B2(n_19),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_97),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_156),
.B(n_141),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_114),
.B1(n_119),
.B2(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_131),
.B1(n_128),
.B2(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_167),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_106),
.B(n_116),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_161),
.B(n_162),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_136),
.C(n_138),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_179),
.C(n_123),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_104),
.B(n_95),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_114),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_174),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_114),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_0),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_34),
.B2(n_1),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_129),
.B(n_146),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_0),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_121),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_124),
.C(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_10),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_156),
.B(n_173),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_196),
.C(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_185),
.B(n_189),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_171),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_205),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_194),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_121),
.C(n_101),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_199),
.B1(n_175),
.B2(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_121),
.B1(n_101),
.B2(n_2),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_8),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_8),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_9),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_214),
.C(n_227),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_155),
.C(n_151),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_223),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_202),
.Y(n_233)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_169),
.B1(n_188),
.B2(n_177),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_178),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_228),
.B(n_181),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_204),
.CI(n_195),
.CON(n_244),
.SN(n_244)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_158),
.B1(n_151),
.B2(n_164),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_225),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_168),
.C(n_163),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_163),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_154),
.B1(n_152),
.B2(n_157),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_230),
.B(n_238),
.CI(n_228),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_191),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_234),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_202),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_196),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_239),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_205),
.C(n_192),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_176),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_246),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_211),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_204),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_7),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_0),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_223),
.B(n_207),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_256),
.B(n_235),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_259),
.B(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_225),
.B1(n_208),
.B2(n_216),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_257),
.B1(n_238),
.B2(n_11),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_241),
.B1(n_223),
.B2(n_226),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_241),
.A2(n_212),
.B(n_224),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_228),
.B1(n_215),
.B2(n_217),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_233),
.Y(n_265)
);

FAx1_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_0),
.CI(n_1),
.CON(n_262),
.SN(n_262)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_260),
.Y(n_264)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_11),
.B(n_15),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_266),
.C(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_236),
.C(n_240),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_240),
.C(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_239),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_274),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_261),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_10),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_256),
.B1(n_255),
.B2(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_277),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_254),
.C(n_262),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_258),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_16),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_6),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_284),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_290),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_265),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_276),
.C(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_6),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_1),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_278),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_3),
.C2(n_2),
.Y(n_293)
);

NOR4xp25_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_296),
.C(n_288),
.D(n_3),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_16),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_287),
.B(n_298),
.C(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_293),
.Y(n_301)
);


endmodule