module fake_aes_10235_n_559 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_559);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_559;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g71 ( .A(n_30), .Y(n_71) );
INVx1_ASAP7_75t_SL g72 ( .A(n_3), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_22), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_4), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_23), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_37), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_5), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_58), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_42), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_19), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_60), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_11), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_36), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_2), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_1), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_61), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_57), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_18), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_46), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_35), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_28), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_47), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_68), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_6), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_4), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_63), .B(n_51), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_45), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_26), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_24), .Y(n_110) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_25), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_53), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_7), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
NOR2xp33_ASAP7_75t_R g117 ( .A(n_83), .B(n_33), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_99), .B(n_0), .Y(n_119) );
INVxp33_ASAP7_75t_SL g120 ( .A(n_99), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_80), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_96), .B(n_0), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_83), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_105), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_89), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_89), .B(n_2), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_75), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
NOR2xp33_ASAP7_75t_R g132 ( .A(n_98), .B(n_34), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_115), .Y(n_133) );
INVxp67_ASAP7_75t_SL g134 ( .A(n_79), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_98), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_87), .B(n_3), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_82), .B(n_5), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_94), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
INVxp33_ASAP7_75t_SL g146 ( .A(n_72), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_85), .A2(n_88), .B1(n_113), .B2(n_87), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_102), .B(n_6), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_102), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_86), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_90), .Y(n_153) );
NOR2xp67_ASAP7_75t_L g154 ( .A(n_90), .B(n_8), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_111), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_122), .Y(n_157) );
OR2x6_ASAP7_75t_L g158 ( .A(n_119), .B(n_88), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_126), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_122), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_135), .B(n_107), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_118), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_124), .B(n_91), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_126), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_135), .B(n_74), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_121), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_120), .B(n_71), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_139), .Y(n_171) );
AO22x2_ASAP7_75t_L g172 ( .A1(n_119), .A2(n_110), .B1(n_114), .B2(n_104), .Y(n_172) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_150), .A2(n_114), .B(n_92), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_127), .B(n_116), .Y(n_175) );
OAI22xp33_ASAP7_75t_SL g176 ( .A1(n_138), .A2(n_113), .B1(n_108), .B2(n_110), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_127), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_144), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_128), .B(n_112), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
AND2x4_ASAP7_75t_SL g182 ( .A(n_129), .B(n_108), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_134), .B(n_139), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
INVx5_ASAP7_75t_L g185 ( .A(n_126), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_130), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_134), .B(n_74), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_137), .B(n_100), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
NAND2x1p5_ASAP7_75t_L g191 ( .A(n_141), .B(n_112), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_142), .B(n_77), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_142), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_129), .B(n_77), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_147), .B(n_104), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_125), .B(n_71), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_153), .B(n_103), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
AOI22x1_ASAP7_75t_L g204 ( .A1(n_155), .A2(n_100), .B1(n_95), .B2(n_76), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_123), .B(n_101), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_154), .B(n_80), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_183), .B(n_103), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_167), .A2(n_190), .B(n_177), .C(n_186), .Y(n_208) );
NOR3xp33_ASAP7_75t_SL g209 ( .A(n_178), .B(n_136), .C(n_156), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_158), .B(n_123), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_206), .Y(n_211) );
AND2x6_ASAP7_75t_L g212 ( .A(n_183), .B(n_76), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_162), .B(n_132), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_158), .B(n_149), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_206), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_206), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_161), .B(n_152), .Y(n_219) );
CKINVDCx8_ASAP7_75t_R g220 ( .A(n_158), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_161), .B(n_117), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_171), .B(n_146), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_162), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_171), .B(n_200), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_200), .B(n_84), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_206), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_172), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_193), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_170), .B(n_97), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_205), .B(n_133), .Y(n_232) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_182), .B(n_80), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_172), .A2(n_80), .B1(n_95), .B2(n_106), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_172), .Y(n_236) );
INVxp67_ASAP7_75t_SL g237 ( .A(n_203), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g238 ( .A1(n_172), .A2(n_80), .B1(n_102), .B2(n_109), .Y(n_238) );
AND3x1_ASAP7_75t_L g239 ( .A(n_196), .B(n_151), .C(n_148), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_193), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_191), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_203), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_191), .B(n_106), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_188), .B(n_109), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_196), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_193), .Y(n_247) );
CKINVDCx8_ASAP7_75t_R g248 ( .A(n_188), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_168), .Y(n_249) );
INVxp67_ASAP7_75t_SL g250 ( .A(n_197), .Y(n_250) );
BUFx12f_ASAP7_75t_L g251 ( .A(n_188), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_168), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_167), .B(n_109), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_188), .B(n_109), .Y(n_254) );
BUFx12f_ASAP7_75t_L g255 ( .A(n_197), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_202), .B(n_109), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_197), .B(n_109), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_179), .B(n_102), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_202), .B(n_102), .Y(n_259) );
NOR2xp33_ASAP7_75t_R g260 ( .A(n_169), .B(n_9), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_257), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_255), .Y(n_263) );
AOI21xp33_ASAP7_75t_L g264 ( .A1(n_219), .A2(n_164), .B(n_176), .Y(n_264) );
INVx6_ASAP7_75t_SL g265 ( .A(n_214), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_224), .A2(n_190), .B(n_199), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_250), .A2(n_197), .B1(n_199), .B2(n_169), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_250), .A2(n_186), .B1(n_177), .B2(n_195), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_252), .B(n_194), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_229), .B(n_194), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g272 ( .A(n_218), .B(n_195), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_224), .A2(n_192), .B(n_184), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_241), .B(n_192), .Y(n_274) );
NOR2xp33_ASAP7_75t_R g275 ( .A(n_220), .B(n_184), .Y(n_275) );
O2A1O1Ixp5_ASAP7_75t_SL g276 ( .A1(n_243), .A2(n_166), .B(n_189), .C(n_175), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_233), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_251), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_230), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_223), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_228), .A2(n_204), .B1(n_173), .B2(n_163), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_230), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_210), .B(n_173), .Y(n_286) );
OR2x6_ASAP7_75t_L g287 ( .A(n_216), .B(n_160), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_240), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_233), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_216), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_244), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_208), .A2(n_140), .B(n_143), .C(n_151), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_225), .B(n_173), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_225), .B(n_204), .Y(n_294) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_214), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_236), .B(n_10), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_247), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_237), .A2(n_160), .B(n_163), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_237), .A2(n_174), .B(n_198), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_212), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_249), .B(n_10), .Y(n_302) );
OR2x6_ASAP7_75t_L g303 ( .A(n_232), .B(n_143), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_272), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_297), .A2(n_212), .B1(n_238), .B2(n_207), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_302), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_301), .B(n_239), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_264), .A2(n_246), .B1(n_222), .B2(n_226), .C(n_221), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_301), .B(n_215), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_275), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_301), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_290), .B(n_212), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_272), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_294), .A2(n_254), .B(n_234), .C(n_238), .Y(n_317) );
AOI221x1_ASAP7_75t_L g318 ( .A1(n_292), .A2(n_259), .B1(n_256), .B2(n_254), .C(n_245), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_297), .A2(n_212), .B1(n_207), .B2(n_226), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_297), .B(n_227), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_291), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_270), .Y(n_322) );
OR2x2_ASAP7_75t_SL g323 ( .A(n_280), .B(n_209), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_282), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_270), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_292), .A2(n_253), .B(n_213), .C(n_145), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_270), .Y(n_327) );
AOI211xp5_ASAP7_75t_L g328 ( .A1(n_311), .A2(n_275), .B(n_260), .C(n_289), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_320), .B(n_274), .Y(n_329) );
INVx4_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_306), .A2(n_267), .B1(n_268), .B2(n_248), .Y(n_332) );
OA21x2_ASAP7_75t_L g333 ( .A1(n_318), .A2(n_283), .B(n_293), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_307), .A2(n_276), .B(n_273), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_306), .A2(n_289), .B1(n_287), .B2(n_278), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_326), .A2(n_286), .B(n_283), .Y(n_336) );
OAI21x1_ASAP7_75t_SL g337 ( .A1(n_319), .A2(n_266), .B(n_261), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_321), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_304), .B(n_303), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_308), .A2(n_231), .B1(n_263), .B2(n_217), .C(n_211), .Y(n_341) );
AOI221x1_ASAP7_75t_L g342 ( .A1(n_317), .A2(n_143), .B1(n_145), .B2(n_148), .C(n_151), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_324), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_319), .A2(n_212), .B1(n_295), .B2(n_207), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_324), .A2(n_300), .B(n_261), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_322), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_317), .A2(n_145), .B(n_148), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_325), .Y(n_349) );
NAND3xp33_ASAP7_75t_L g350 ( .A(n_326), .B(n_213), .C(n_282), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_327), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_332), .A2(n_309), .B1(n_316), .B2(n_304), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_336), .A2(n_310), .B(n_315), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_343), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_332), .A2(n_295), .B1(n_265), .B2(n_207), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_328), .A2(n_316), .B1(n_287), .B2(n_310), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_329), .B(n_274), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_329), .B(n_312), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_341), .A2(n_263), .B1(n_258), .B2(n_288), .C(n_285), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_347), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_347), .B(n_274), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_339), .B(n_290), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_335), .B(n_314), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_347), .Y(n_366) );
AO21x2_ASAP7_75t_L g367 ( .A1(n_350), .A2(n_253), .B(n_299), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_341), .A2(n_258), .B1(n_284), .B2(n_281), .C(n_313), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_339), .B(n_323), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_340), .A2(n_313), .B1(n_298), .B2(n_312), .C(n_277), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_331), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_351), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_340), .B(n_338), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_331), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
OAI22xp33_ASAP7_75t_SL g378 ( .A1(n_335), .A2(n_314), .B1(n_277), .B2(n_262), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_338), .B(n_207), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_328), .B(n_312), .C(n_262), .Y(n_380) );
BUFx4f_ASAP7_75t_SL g381 ( .A(n_330), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_344), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_375), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_362), .B(n_348), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_360), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_362), .B(n_348), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_378), .A2(n_352), .B(n_348), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_366), .B(n_348), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_364), .B(n_351), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_360), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_364), .B(n_363), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_356), .A2(n_345), .B(n_352), .C(n_330), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_365), .B(n_344), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_373), .B(n_349), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_374), .B(n_349), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_355), .B(n_333), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_369), .A2(n_337), .B1(n_298), .B2(n_350), .C(n_344), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_363), .B(n_333), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_381), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
NAND2xp33_ASAP7_75t_R g405 ( .A(n_365), .B(n_377), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_365), .B(n_342), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_357), .A2(n_333), .B1(n_314), .B2(n_296), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_365), .A2(n_265), .B1(n_333), .B2(n_279), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_372), .B(n_342), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_370), .B(n_334), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_376), .B(n_282), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_370), .B(n_334), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_358), .B(n_12), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_353), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_404), .B(n_354), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_383), .B(n_371), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
NOR2xp33_ASAP7_75t_R g425 ( .A(n_402), .B(n_13), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_392), .B(n_15), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_390), .B(n_16), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_399), .B(n_367), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_396), .B(n_368), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_417), .B(n_16), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_384), .B(n_367), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_396), .B(n_361), .Y(n_432) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_405), .B(n_367), .Y(n_433) );
NAND2xp33_ASAP7_75t_R g434 ( .A(n_406), .B(n_346), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
OAI31xp33_ASAP7_75t_SL g437 ( .A1(n_385), .A2(n_265), .A3(n_271), .B(n_296), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_398), .B(n_279), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_387), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_403), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_403), .B(n_20), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_407), .B(n_27), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_391), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_416), .B(n_31), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_400), .B(n_165), .C(n_201), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_411), .B(n_32), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_386), .B(n_38), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_389), .B(n_39), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_389), .B(n_40), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_412), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_401), .B(n_41), .Y(n_452) );
NAND4xp75_ASAP7_75t_L g453 ( .A(n_408), .B(n_43), .C(n_44), .D(n_48), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_411), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_407), .B(n_174), .Y(n_455) );
NAND2xp33_ASAP7_75t_SL g456 ( .A(n_405), .B(n_49), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_414), .B(n_55), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_418), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_406), .B(n_242), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_420), .B(n_56), .Y(n_461) );
INVx6_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_424), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_446), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_458), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_443), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_460), .A2(n_419), .B1(n_420), .B2(n_406), .Y(n_468) );
AND3x2_ASAP7_75t_L g469 ( .A(n_437), .B(n_394), .C(n_410), .Y(n_469) );
OAI21xp33_ASAP7_75t_SL g470 ( .A1(n_454), .A2(n_388), .B(n_409), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_460), .B(n_419), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_456), .A2(n_393), .B(n_410), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_456), .B(n_410), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_425), .A2(n_413), .B1(n_421), .B2(n_415), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_440), .Y(n_475) );
INVxp67_ASAP7_75t_L g476 ( .A(n_454), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_425), .A2(n_415), .B(n_413), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_435), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_426), .B(n_59), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_430), .B(n_62), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_451), .B(n_64), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_422), .B(n_66), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_460), .A2(n_67), .B1(n_181), .B2(n_180), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_422), .B(n_157), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_441), .B(n_159), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_423), .A2(n_159), .B1(n_165), .B2(n_187), .C(n_201), .Y(n_487) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_459), .A2(n_159), .B(n_165), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_460), .A2(n_185), .B1(n_165), .B2(n_159), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_442), .A2(n_166), .B(n_185), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_431), .B(n_165), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_429), .A2(n_187), .B1(n_201), .B2(n_166), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_432), .A2(n_166), .B1(n_185), .B2(n_187), .C1(n_201), .C2(n_461), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_427), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_428), .B(n_187), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_459), .B(n_185), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_495), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_472), .A2(n_434), .B1(n_462), .B2(n_445), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_465), .B(n_462), .Y(n_501) );
NAND2xp33_ASAP7_75t_SL g502 ( .A(n_473), .B(n_434), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_496), .B(n_452), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_464), .Y(n_505) );
XOR2x2_ASAP7_75t_L g506 ( .A(n_469), .B(n_447), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_467), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_472), .B(n_433), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_470), .B(n_449), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_476), .B(n_444), .Y(n_510) );
NAND2xp33_ASAP7_75t_SL g511 ( .A(n_468), .B(n_450), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_477), .B(n_453), .C(n_455), .Y(n_512) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_485), .B(n_457), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_490), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_471), .B(n_448), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_475), .B(n_185), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_474), .B(n_489), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_486), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_507), .B(n_478), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_508), .B(n_483), .C(n_482), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_509), .A2(n_494), .B(n_479), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_509), .A2(n_483), .B(n_491), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_500), .B(n_491), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_504), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_502), .B(n_489), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_499), .B(n_480), .Y(n_527) );
AOI211xp5_ASAP7_75t_L g528 ( .A1(n_500), .A2(n_487), .B(n_484), .C(n_481), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_508), .A2(n_494), .B1(n_492), .B2(n_497), .C(n_493), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_505), .Y(n_531) );
BUFx4f_ASAP7_75t_SL g532 ( .A(n_518), .Y(n_532) );
NAND3xp33_ASAP7_75t_SL g533 ( .A(n_518), .B(n_488), .C(n_498), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_501), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_514), .B(n_488), .Y(n_535) );
XOR2xp5_ASAP7_75t_L g536 ( .A(n_506), .B(n_516), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_511), .A2(n_512), .B1(n_503), .B2(n_510), .Y(n_537) );
XNOR2xp5_ASAP7_75t_L g538 ( .A(n_536), .B(n_516), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_525), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_537), .B(n_519), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_531), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_524), .B(n_513), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_534), .B(n_515), .Y(n_543) );
OAI321xp33_ASAP7_75t_L g544 ( .A1(n_522), .A2(n_517), .A3(n_526), .B1(n_523), .B2(n_529), .C(n_528), .Y(n_544) );
NAND3x1_ASAP7_75t_SL g545 ( .A(n_521), .B(n_527), .C(n_535), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_520), .A2(n_527), .B1(n_530), .B2(n_537), .C(n_533), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_532), .A2(n_537), .B1(n_536), .B2(n_509), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_523), .A2(n_522), .B(n_537), .C(n_524), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_538), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_543), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_548), .B(n_540), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_551), .B(n_547), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g553 ( .A(n_550), .B(n_544), .Y(n_553) );
AO22x2_ASAP7_75t_L g554 ( .A1(n_549), .A2(n_545), .B1(n_539), .B2(n_541), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_553), .B(n_550), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_552), .Y(n_556) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_556), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_557), .A2(n_555), .B1(n_554), .B2(n_546), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_558), .A2(n_555), .B(n_542), .Y(n_559) );
endmodule