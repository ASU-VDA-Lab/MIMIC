module fake_jpeg_8569_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_31),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.C(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_17),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_32),
.B1(n_20),
.B2(n_39),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_52),
.B1(n_57),
.B2(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_45),
.B(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_25),
.B1(n_17),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_36),
.B1(n_28),
.B2(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_37),
.B1(n_19),
.B2(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_31),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_56),
.B1(n_50),
.B2(n_47),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_70),
.B1(n_75),
.B2(n_47),
.Y(n_87)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_24),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_46),
.B1(n_49),
.B2(n_23),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_77),
.C(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_13),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_18),
.B1(n_31),
.B2(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_42),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_42),
.A3(n_33),
.B1(n_23),
.B2(n_4),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_48),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_87),
.B1(n_77),
.B2(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_9),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_63),
.Y(n_105)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_66),
.C(n_79),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_115),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_88),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_73),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_81),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_62),
.B(n_68),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_106),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_120),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_91),
.B1(n_96),
.B2(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_91),
.B1(n_86),
.B2(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_134),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_103),
.C(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_141),
.B1(n_5),
.B2(n_6),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_116),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_137),
.A2(n_116),
.B(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_5),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_108),
.B1(n_100),
.B2(n_109),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_99),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_14),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_129),
.B1(n_127),
.B2(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_148),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_132),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_152),
.B(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_92),
.B1(n_120),
.B2(n_7),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_134),
.C(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_154),
.B(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_135),
.C(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_144),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_164),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_149),
.B1(n_145),
.B2(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_162),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_164),
.B(n_131),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_158),
.B(n_159),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_165),
.B(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_163),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_169),
.C(n_10),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_14),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_174),
.Y(n_177)
);


endmodule