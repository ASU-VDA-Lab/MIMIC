module real_jpeg_33058_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_0),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_147),
.B1(n_151),
.B2(n_156),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_1),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_1),
.A2(n_156),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_4),
.Y(n_102)
);

OAI22x1_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_102),
.B1(n_159),
.B2(n_166),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_4),
.A2(n_102),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_8),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_8),
.A2(n_173),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_8),
.A2(n_34),
.B(n_251),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_12),
.A2(n_86),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_12),
.A2(n_92),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_12),
.A2(n_92),
.B1(n_260),
.B2(n_264),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_225),
.Y(n_13)
);

NAND2xp33_ASAP7_75t_R g14 ( 
.A(n_15),
.B(n_223),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_201),
.Y(n_16)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_17),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_117),
.B2(n_118),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_68),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

OAI22x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B1(n_41),
.B2(n_49),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_22),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_27),
.Y(n_194)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_27),
.Y(n_309)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_28),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_30),
.Y(n_264)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_33),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_34),
.A2(n_245),
.B(n_251),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_35),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_35),
.A2(n_258),
.B1(n_265),
.B2(n_268),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_37),
.Y(n_190)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_37),
.Y(n_253)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_38),
.Y(n_248)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_61),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_84),
.B(n_96),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_69),
.B(n_173),
.Y(n_242)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_70),
.B(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx5_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_90),
.Y(n_218)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_106),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_170),
.B1(n_199),
.B2(n_200),
.Y(n_118)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_146),
.B(n_157),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_120),
.A2(n_146),
.B1(n_205),
.B2(n_213),
.Y(n_204)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_120),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_132),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_136),
.B1(n_139),
.B2(n_142),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_135),
.Y(n_289)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_138),
.Y(n_300)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_153),
.Y(n_279)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_157),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_158),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_189),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_189),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_176),
.B1(n_180),
.B2(n_184),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_173),
.B(n_291),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g297 ( 
.A1(n_173),
.A2(n_290),
.B(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_173),
.B(n_253),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_173),
.B(n_213),
.Y(n_311)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_185),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_191),
.A2(n_259),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.C(n_214),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_230),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B(n_222),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_254),
.B(n_326),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_231),
.B(n_233),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_229),
.B(n_232),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_233),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.C(n_243),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_236),
.B(n_242),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_297),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_243),
.A2(n_244),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_320),
.B(n_325),
.Y(n_254)
);

AO21x1_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_301),
.B(n_319),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_269),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_269),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_295),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_R g321 ( 
.A(n_270),
.B(n_295),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_277),
.B(n_285),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_288),
.B(n_290),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx4f_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_310),
.B(n_318),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_312),
.Y(n_318)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);


endmodule