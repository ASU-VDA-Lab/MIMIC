module real_jpeg_18342_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_92),
.B1(n_97),
.B2(n_101),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_0),
.A2(n_70),
.B1(n_101),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_2),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_3),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_3),
.A2(n_208),
.B1(n_536),
.B2(n_540),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_4),
.A2(n_135),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_4),
.A2(n_135),
.B1(n_336),
.B2(n_339),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_4),
.A2(n_135),
.B1(n_431),
.B2(n_434),
.Y(n_430)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_5),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_6),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_6),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_76),
.B1(n_80),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_7),
.A2(n_82),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_7),
.A2(n_82),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_8),
.A2(n_126),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_8),
.A2(n_126),
.B1(n_381),
.B2(n_384),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_8),
.A2(n_126),
.B1(n_446),
.B2(n_449),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_9),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_9),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_9),
.A2(n_263),
.B(n_325),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g346 ( 
.A1(n_9),
.A2(n_338),
.A3(n_347),
.B1(n_351),
.B2(n_353),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_9),
.A2(n_311),
.B1(n_393),
.B2(n_397),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_9),
.B(n_249),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_9),
.A2(n_83),
.B1(n_470),
.B2(n_478),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_10),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_10),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_10),
.A2(n_279),
.B1(n_290),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_10),
.A2(n_70),
.B1(n_279),
.B2(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_10),
.A2(n_279),
.B1(n_471),
.B2(n_474),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_11),
.A2(n_69),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_11),
.A2(n_69),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_12),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_12),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_14),
.A2(n_58),
.B1(n_175),
.B2(n_180),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_14),
.A2(n_58),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_14),
.A2(n_58),
.B1(n_128),
.B2(n_549),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_16),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_16),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_16),
.A2(n_145),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_16),
.A2(n_145),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_16),
.A2(n_145),
.B1(n_357),
.B2(n_361),
.Y(n_356)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_17),
.Y(n_125)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_17),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_517),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_280),
.B(n_514),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_235),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_22),
.B(n_235),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_184),
.Y(n_22)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_23),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_105),
.C(n_139),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_25),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_74),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_26),
.A2(n_27),
.B1(n_74),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_27)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_28),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_28),
.B(n_64),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_28),
.A2(n_62),
.B1(n_335),
.B2(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_28),
.A2(n_62),
.B1(n_421),
.B2(n_425),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_28),
.A2(n_62),
.B1(n_380),
.B2(n_425),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_28),
.A2(n_62),
.B1(n_534),
.B2(n_535),
.Y(n_533)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_34),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_34),
.Y(n_207)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_34),
.Y(n_271)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_34),
.Y(n_309)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_34),
.Y(n_418)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_35),
.Y(n_363)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_36),
.Y(n_464)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_37),
.Y(n_408)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_37),
.Y(n_473)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_51),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_42),
.Y(n_168)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_43),
.Y(n_383)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_49),
.Y(n_410)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_52),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_55),
.Y(n_352)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_57),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_57),
.Y(n_427)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_62),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_63),
.A2(n_187),
.B1(n_188),
.B2(n_196),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_63),
.A2(n_187),
.B1(n_315),
.B2(n_320),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_63),
.A2(n_187),
.B1(n_315),
.B2(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_63),
.B(n_311),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_68),
.Y(n_317)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_74),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_83),
.B1(n_91),
.B2(n_102),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_75),
.A2(n_83),
.B1(n_202),
.B2(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_78),
.Y(n_307)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_78),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_83),
.A2(n_202),
.B(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_83),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_83),
.A2(n_230),
.B1(n_430),
.B2(n_435),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_83),
.A2(n_445),
.B1(n_470),
.B2(n_482),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_84),
.A2(n_227),
.B1(n_268),
.B2(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_84),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_86),
.Y(n_484)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_87),
.Y(n_231)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_90),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_91),
.Y(n_228)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_96),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_99),
.Y(n_477)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_100),
.Y(n_433)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_105),
.B(n_140),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_123),
.B1(n_132),
.B2(n_138),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_106),
.A2(n_132),
.B1(n_138),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_106),
.A2(n_123),
.B1(n_138),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_106),
.A2(n_138),
.B1(n_275),
.B2(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_106),
.A2(n_138),
.B1(n_213),
.B2(n_548),
.Y(n_547)
);

AO21x2_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_116),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_107),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_108),
.Y(n_327)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_120),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_120),
.Y(n_262)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_121),
.Y(n_295)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_130),
.Y(n_277)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_130),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_134),
.Y(n_278)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_138),
.B(n_311),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_149),
.B1(n_173),
.B2(n_174),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_142),
.A2(n_150),
.B1(n_242),
.B2(n_249),
.Y(n_241)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

OAI22x1_ASAP7_75t_SL g217 ( 
.A1(n_149),
.A2(n_173),
.B1(n_174),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_149),
.A2(n_173),
.B1(n_289),
.B2(n_296),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_149),
.A2(n_173),
.B1(n_296),
.B2(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_149),
.A2(n_173),
.B1(n_289),
.B2(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_150),
.A2(n_249),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_158),
.B(n_164),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_157),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_158),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_162),
.Y(n_302)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_163),
.Y(n_293)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_163),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_163),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_169),
.B2(n_172),
.Y(n_164)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_171),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g424 ( 
.A(n_171),
.Y(n_424)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_171),
.Y(n_539)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_179),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_180),
.Y(n_297)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_210),
.B1(n_233),
.B2(n_234),
.Y(n_184)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_185),
.B(n_234),
.C(n_520),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_200),
.B1(n_201),
.B2(n_209),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_186),
.B(n_201),
.Y(n_543)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_195),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_196),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_200),
.A2(n_201),
.B1(n_546),
.B2(n_547),
.Y(n_545)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_204),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_222),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_212),
.B(n_217),
.C(n_222),
.Y(n_522)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_218),
.Y(n_526)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B(n_226),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_232),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_227),
.A2(n_305),
.B1(n_356),
.B2(n_364),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_227),
.A2(n_444),
.B1(n_453),
.B2(n_454),
.Y(n_443)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_236),
.B(n_238),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_240),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_250),
.C(n_273),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_241),
.A2(n_273),
.B1(n_274),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_241),
.Y(n_503)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

INVx8_ASAP7_75t_L g529 ( 
.A(n_243),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_250),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_266),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_266),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_263),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_271),
.Y(n_452)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_497),
.B(n_511),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_370),
.B(n_496),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_328),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_284),
.B(n_328),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_312),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_286),
.B(n_287),
.C(n_312),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_303),
.C(n_310),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_288),
.B(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_303),
.A2(n_304),
.B1(n_310),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_311),
.B(n_412),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_SL g421 ( 
.A1(n_311),
.A2(n_411),
.B(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_311),
.B(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_323),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_321),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g506 ( 
.A(n_314),
.B(n_321),
.C(n_323),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_319),
.Y(n_540)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.C(n_344),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_330),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_333),
.A2(n_344),
.B1(n_345),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_354),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_354),
.B1(n_355),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_400),
.B(n_495),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_376),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_372),
.B(n_376),
.Y(n_495)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.C(n_390),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_377),
.B(n_492),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_379),
.A2(n_390),
.B1(n_391),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx8_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI21x1_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_489),
.B(n_494),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_441),
.B(n_488),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_428),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_403),
.B(n_428),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_419),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_404),
.A2(n_419),
.B1(n_420),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

OAI32xp33_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_407),
.A3(n_409),
.B1(n_411),
.B2(n_413),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_409),
.Y(n_414)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_436),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_429),
.B(n_438),
.C(n_440),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_430),
.Y(n_454)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_436)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_437),
.Y(n_440)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_457),
.B(n_487),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_455),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_455),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_480),
.B(n_486),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_469),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_465),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_485),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_485),
.Y(n_486)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_SL g494 ( 
.A(n_490),
.B(n_491),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_500),
.B(n_507),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_500),
.C(n_513),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.C(n_506),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_501),
.B(n_509),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_506),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_510),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_552),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_519),
.B(n_521),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_542),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_525),
.A2(n_533),
.B(n_541),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_533),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_543),
.A2(n_544),
.B1(n_545),
.B2(n_551),
.Y(n_542)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_543),
.Y(n_551)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);


endmodule