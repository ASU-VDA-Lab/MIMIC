module real_jpeg_9338_n_11 (n_239, n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_239;
input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_8),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_0),
.A2(n_1),
.B1(n_21),
.B2(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_10),
.B1(n_21),
.B2(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_31),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_35),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_2),
.B(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_4),
.A2(n_9),
.B(n_51),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_5),
.A2(n_6),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_21),
.B(n_24),
.C(n_28),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g28 ( 
.A(n_5),
.B(n_21),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_6),
.A3(n_21),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_49),
.B(n_52),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_6),
.B(n_52),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_8),
.B1(n_20),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_9),
.B1(n_26),
.B2(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_32),
.B(n_52),
.C(n_124),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_10),
.B1(n_26),
.B2(n_40),
.Y(n_201)
);

HAxp5_ASAP7_75t_SL g31 ( 
.A(n_7),
.B(n_32),
.CON(n_31),
.SN(n_31)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_10),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_20),
.B1(n_50),
.B2(n_51),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_21),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_32),
.B1(n_50),
.B2(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_9),
.B(n_41),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_9),
.B(n_24),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_71),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_70),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_57),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_15),
.B(n_57),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_56),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_29),
.B2(n_30),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_24),
.B1(n_27),
.B2(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_38),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_23),
.B(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_24),
.A2(n_27),
.B1(n_47),
.B2(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_25),
.B(n_26),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_39),
.B2(n_41),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_32),
.B(n_49),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_32),
.B(n_91),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.C(n_48),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_83),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_60),
.B1(n_83),
.B2(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_44),
.A2(n_60),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_44),
.B(n_83),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_44),
.A2(n_60),
.B1(n_196),
.B2(n_197),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_44),
.A2(n_60),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_44),
.A2(n_197),
.B(n_213),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_44),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_48),
.A2(n_64),
.B1(n_66),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_53),
.B(n_55),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_53),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_49),
.A2(n_53),
.B1(n_81),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_50),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_65),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_64),
.C(n_66),
.Y(n_65)
);

AOI211xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_80),
.B(n_82),
.C(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_65),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_66),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_69),
.Y(n_146)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_221),
.A3(n_231),
.B1(n_236),
.B2(n_237),
.C(n_239),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_207),
.B(n_220),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_188),
.B(n_206),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_116),
.B(n_172),
.C(n_187),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_104),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_76),
.B(n_104),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_95),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_88),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_78),
.B(n_88),
.C(n_95),
.Y(n_173)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_85),
.B1(n_89),
.B2(n_94),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_85),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_85),
.B1(n_123),
.B2(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_102),
.C(n_127),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_80),
.A2(n_85),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_155),
.C(n_161),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_80),
.A2(n_85),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_80),
.B(n_89),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_80),
.B(n_178),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_83),
.A2(n_85),
.B(n_149),
.C(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_83),
.A2(n_84),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_102),
.C(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_84),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_84),
.B(n_216),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_86),
.A2(n_103),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_86),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_179),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_103),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_96),
.A2(n_97),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_96),
.A2(n_97),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_102),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_111),
.B1(n_126),
.B2(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_111),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_102),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_145),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_113),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_106),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_108),
.B1(n_144),
.B2(n_149),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_138),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_171),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_164),
.B(n_170),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_151),
.B(n_163),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_141),
.B(n_150),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_130),
.B(n_140),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_143),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_173),
.B(n_174),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_185),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_184),
.C(n_185),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_190),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_203),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_195),
.C(n_203),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_193),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_204),
.B(n_205),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_202),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_200),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_209),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_218),
.B2(n_219),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_215),
.C(n_219),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_223),
.C(n_227),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_229),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_227),
.A2(n_228),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);


endmodule