module fake_jpeg_30917_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_4),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_59),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_1),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_64),
.Y(n_72)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_19),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_54),
.C(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_2),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_48),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_77),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_56),
.B1(n_46),
.B2(n_45),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_56),
.B1(n_46),
.B2(n_42),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_55),
.B1(n_52),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_43),
.B1(n_55),
.B2(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_54),
.B1(n_51),
.B2(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_49),
.C(n_3),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_21),
.B1(n_40),
.B2(n_39),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_18),
.C(n_38),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_83),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_66),
.B(n_77),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_102),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_101),
.B1(n_11),
.B2(n_16),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_37),
.B(n_27),
.C(n_28),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_104),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_9),
.B(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_109),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_30),
.C(n_35),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_117),
.C(n_92),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_115),
.B1(n_97),
.B2(n_102),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_31),
.C(n_14),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_25),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_107),
.B1(n_116),
.B2(n_92),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_102),
.B(n_106),
.C(n_36),
.D(n_32),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_125),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_126),
.Y(n_127)
);

AOI21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_122),
.B(n_118),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_124),
.B(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_125),
.C(n_114),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_33),
.Y(n_131)
);


endmodule