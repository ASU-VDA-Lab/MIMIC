module fake_jpeg_3412_n_226 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_27),
.B(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_22),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_2),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_3),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_51),
.Y(n_96)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_69),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_89),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_96),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_78),
.B(n_74),
.C(n_61),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_98),
.B(n_60),
.C(n_54),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_54),
.B(n_60),
.C(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_112),
.Y(n_131)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_82),
.B1(n_89),
.B2(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_65),
.B1(n_68),
.B2(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_66),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_59),
.B1(n_70),
.B2(n_63),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_70),
.B1(n_63),
.B2(n_57),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_100),
.C(n_104),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_26),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_129),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_59),
.B(n_65),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_29),
.B(n_48),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_125),
.B1(n_68),
.B2(n_28),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_114),
.B1(n_104),
.B2(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_133),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_65),
.B1(n_62),
.B2(n_71),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_24),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_62),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_124),
.B1(n_129),
.B2(n_117),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_122),
.B1(n_32),
.B2(n_33),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_147),
.B1(n_151),
.B2(n_14),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_4),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_136),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_4),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_148),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_6),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_15),
.B(n_16),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_7),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_35),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_34),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_175),
.Y(n_186)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_41),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_18),
.B(n_20),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_179),
.B(n_163),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_141),
.B1(n_155),
.B2(n_21),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_190),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_171),
.B(n_161),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_178),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_38),
.B(n_40),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_170),
.B(n_162),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_177),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_202),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_187),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_160),
.B(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_192),
.C(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_195),
.B1(n_191),
.B2(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_197),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_216),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_212),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_208),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_218),
.C(n_195),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_215),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_222),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_214),
.C(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_206),
.B(n_47),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_43),
.Y(n_226)
);


endmodule