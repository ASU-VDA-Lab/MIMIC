module fake_jpeg_28670_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_58),
.B1(n_42),
.B2(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_60),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_6),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_72),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_10),
.B(n_11),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_47),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_8),
.Y(n_88)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_49),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_6),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_48),
.B1(n_42),
.B2(n_44),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_89),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_45),
.B(n_50),
.C(n_8),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_92),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_50),
.B(n_53),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_73),
.C(n_14),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_43),
.B1(n_20),
.B2(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_84),
.B1(n_25),
.B2(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_7),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_7),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_91),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_10),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_23),
.B(n_32),
.C(n_12),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_77),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_13),
.B(n_15),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_106),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_18),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_78),
.B1(n_76),
.B2(n_31),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_96),
.B1(n_94),
.B2(n_99),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_101),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.C(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_96),
.C(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_113),
.B1(n_95),
.B2(n_99),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.Y(n_120)
);

AOI31xp67_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_112),
.A3(n_97),
.B(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_28),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_29),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_109),
.Y(n_124)
);


endmodule