module fake_netlist_1_6210_n_743 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_743);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_743;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_22), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_11), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_63), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_3), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_66), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_8), .Y(n_91) );
BUFx10_ASAP7_75t_L g92 ( .A(n_80), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_3), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_24), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_44), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_39), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_27), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_75), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_65), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_28), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_34), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_30), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_7), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_36), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_41), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_33), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_11), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_42), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_55), .Y(n_110) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_60), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_68), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_9), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_54), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
BUFx10_ASAP7_75t_L g118 ( .A(n_21), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_40), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_46), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_52), .Y(n_121) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_31), .B(n_71), .Y(n_122) );
INVx2_ASAP7_75t_SL g123 ( .A(n_49), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_56), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_76), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_5), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_10), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_23), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_127), .B(n_0), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_86), .B(n_0), .Y(n_136) );
CKINVDCx6p67_ASAP7_75t_R g137 ( .A(n_87), .Y(n_137) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_89), .A2(n_38), .B(n_79), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_109), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_123), .B(n_1), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_123), .B(n_1), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_84), .B(n_2), .Y(n_146) );
INVx1_ASAP7_75t_SL g147 ( .A(n_119), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_86), .B(n_2), .Y(n_148) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_94), .A2(n_43), .B(n_78), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_115), .B(n_4), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_82), .B(n_4), .Y(n_154) );
BUFx8_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_95), .Y(n_156) );
BUFx8_ASAP7_75t_L g157 ( .A(n_97), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_97), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_85), .B(n_5), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_130), .B(n_6), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_98), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_98), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_99), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_92), .B(n_9), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_101), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_102), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_115), .B(n_10), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_85), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_102), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_103), .Y(n_172) );
NOR3xp33_ASAP7_75t_L g173 ( .A(n_91), .B(n_12), .C(n_13), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_91), .B(n_12), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_92), .B(n_13), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_103), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_165), .B(n_129), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_170), .B(n_88), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_137), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_170), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_132), .B(n_108), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_137), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_167), .B(n_131), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_132), .B(n_108), .Y(n_192) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_148), .B(n_131), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_138), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_148), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_152), .B(n_129), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_152), .B(n_104), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_152), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_135), .B(n_112), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_169), .B(n_104), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_135), .B(n_110), .Y(n_208) );
NOR2x1p5_ASAP7_75t_L g209 ( .A(n_137), .B(n_113), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_169), .B(n_125), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_147), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_141), .B(n_128), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_141), .B(n_96), .Y(n_214) );
OAI221xp5_ASAP7_75t_L g215 ( .A1(n_150), .A2(n_93), .B1(n_125), .B2(n_107), .C(n_117), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_169), .B(n_128), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_143), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_143), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_156), .B(n_100), .Y(n_223) );
NAND3x1_ASAP7_75t_L g224 ( .A(n_173), .B(n_126), .C(n_121), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_165), .B(n_126), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_156), .B(n_117), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_145), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_145), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_167), .B(n_171), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_155), .A2(n_111), .B1(n_105), .B2(n_121), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_160), .B(n_92), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_142), .Y(n_233) );
NAND3xp33_ASAP7_75t_L g234 ( .A(n_155), .B(n_120), .C(n_116), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_160), .B(n_118), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_175), .B(n_120), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_151), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_167), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_151), .Y(n_239) );
AND2x6_ASAP7_75t_L g240 ( .A(n_171), .B(n_116), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_142), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_166), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_158), .B(n_106), .Y(n_243) );
AO22x2_ASAP7_75t_L g244 ( .A1(n_173), .A2(n_176), .B1(n_161), .B2(n_162), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_221), .B(n_155), .Y(n_245) );
INVx5_ASAP7_75t_L g246 ( .A(n_240), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_233), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_181), .Y(n_249) );
NAND2x1_ASAP7_75t_L g250 ( .A(n_240), .B(n_149), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_241), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_187), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_240), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_227), .A2(n_149), .B(n_158), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_240), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_193), .A2(n_157), .B1(n_155), .B2(n_171), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_228), .B(n_134), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_210), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_179), .B(n_157), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_177), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_183), .B(n_134), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_225), .B(n_157), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_183), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_180), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_183), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_240), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_192), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_225), .B(n_157), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_193), .A2(n_147), .B1(n_174), .B2(n_159), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_210), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_225), .B(n_176), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_210), .Y(n_275) );
OR2x6_ASAP7_75t_L g276 ( .A(n_178), .B(n_174), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_244), .A2(n_162), .B1(n_168), .B2(n_161), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_199), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_178), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_192), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_180), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_232), .B(n_168), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_190), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_192), .B(n_163), .Y(n_286) );
INVxp67_ASAP7_75t_SL g287 ( .A(n_238), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_200), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_190), .Y(n_289) );
OR2x6_ASAP7_75t_L g290 ( .A(n_209), .B(n_159), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_200), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_187), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_200), .B(n_154), .Y(n_293) );
INVx2_ASAP7_75t_SL g294 ( .A(n_218), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_205), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_207), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_185), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_207), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_235), .B(n_163), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_206), .B(n_172), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_191), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_214), .B(n_172), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_231), .A2(n_146), .B1(n_154), .B2(n_164), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_218), .Y(n_304) );
OR2x4_ASAP7_75t_L g305 ( .A(n_208), .B(n_166), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_223), .B(n_172), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_205), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
INVxp33_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_215), .B(n_118), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_182), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_177), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_229), .Y(n_314) );
NOR2xp33_ASAP7_75t_R g315 ( .A(n_184), .B(n_118), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_188), .B(n_164), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_177), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_263), .A2(n_244), .B1(n_195), .B2(n_197), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_307), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_262), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_317), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_247), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_276), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_280), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_266), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_266), .Y(n_329) );
BUFx12f_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_254), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_255), .Y(n_333) );
BUFx4f_ASAP7_75t_SL g334 ( .A(n_281), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_268), .B(n_234), .Y(n_335) );
AOI21xp5_ASAP7_75t_SL g336 ( .A1(n_255), .A2(n_149), .B(n_186), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_264), .A2(n_236), .B1(n_198), .B2(n_201), .Y(n_337) );
BUFx4f_ASAP7_75t_L g338 ( .A(n_276), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_247), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_309), .B(n_236), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_263), .A2(n_244), .B1(n_217), .B2(n_189), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_259), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_251), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_262), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_268), .B(n_186), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_262), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_257), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_282), .A2(n_213), .B(n_243), .C(n_226), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_309), .B(n_213), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_270), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_251), .Y(n_352) );
CKINVDCx11_ASAP7_75t_R g353 ( .A(n_281), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_280), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_262), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_262), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_270), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_246), .B(n_177), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_257), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_312), .Y(n_361) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_283), .B(n_186), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_252), .A2(n_189), .B(n_229), .C(n_142), .Y(n_363) );
CKINVDCx6p67_ASAP7_75t_R g364 ( .A(n_276), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_278), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_279), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_259), .B(n_224), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_299), .B(n_164), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_269), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_284), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_279), .B(n_186), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_313), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_299), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_322), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_342), .A2(n_374), .B1(n_334), .B2(n_368), .C1(n_349), .C2(n_353), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_322), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_369), .B(n_293), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_330), .A2(n_267), .B1(n_315), .B2(n_272), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_336), .A2(n_250), .B(n_256), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_368), .A2(n_248), .B1(n_249), .B2(n_290), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_354), .A2(n_290), .B1(n_310), .B2(n_293), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_345), .A2(n_245), .B(n_317), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_324), .A2(n_290), .B1(n_293), .B2(n_298), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_322), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_323), .Y(n_387) );
BUFx8_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
AOI21xp5_ASAP7_75t_SL g389 ( .A1(n_322), .A2(n_317), .B(n_312), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_327), .A2(n_290), .B1(n_298), .B2(n_313), .Y(n_390) );
BUFx10_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_364), .B(n_286), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_327), .B(n_294), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_331), .A2(n_303), .B(n_277), .C(n_274), .Y(n_394) );
CKINVDCx6p67_ASAP7_75t_R g395 ( .A(n_364), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_332), .B(n_267), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_338), .A2(n_258), .B1(n_294), .B2(n_304), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_338), .A2(n_304), .B1(n_265), .B2(n_271), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_369), .B(n_285), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_338), .B(n_288), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_336), .A2(n_317), .B(n_312), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g403 ( .A1(n_363), .A2(n_302), .B(n_300), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_338), .A2(n_291), .B1(n_296), .B2(n_308), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_367), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_318), .A2(n_305), .B1(n_260), .B2(n_273), .Y(n_406) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_326), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_325), .A2(n_289), .B1(n_283), .B2(n_295), .Y(n_408) );
BUFx4f_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_380), .A2(n_339), .B(n_346), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_376), .A2(n_330), .B1(n_340), .B2(n_325), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_376), .A2(n_330), .B1(n_261), .B2(n_373), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_401), .A2(n_322), .B(n_355), .Y(n_413) );
NOR2x1_ASAP7_75t_SL g414 ( .A(n_407), .B(n_339), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
AOI222xp33_ASAP7_75t_L g416 ( .A1(n_378), .A2(n_365), .B1(n_366), .B2(n_371), .C1(n_275), .C2(n_348), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_386), .B(n_343), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_365), .B1(n_337), .B2(n_341), .C(n_366), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
BUFx4f_ASAP7_75t_SL g422 ( .A(n_395), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_387), .A2(n_343), .B1(n_352), .B2(n_305), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_395), .A2(n_305), .B1(n_358), .B2(n_352), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_379), .A2(n_373), .B1(n_351), .B2(n_328), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_396), .A2(n_328), .B1(n_329), .B2(n_351), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_397), .A2(n_398), .B1(n_382), .B2(n_378), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_381), .A2(n_371), .B1(n_306), .B2(n_153), .C(n_316), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_399), .B(n_372), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_406), .A2(n_153), .B1(n_287), .B2(n_335), .C(n_140), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_393), .A2(n_329), .B1(n_372), .B2(n_319), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_399), .Y(n_435) );
OAI222xp33_ASAP7_75t_L g436 ( .A1(n_384), .A2(n_392), .B1(n_390), .B2(n_405), .C1(n_393), .C2(n_400), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_393), .A2(n_319), .B1(n_320), .B2(n_350), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_409), .A2(n_153), .B1(n_196), .B2(n_355), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_411), .A2(n_393), .B1(n_388), .B2(n_400), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_412), .A2(n_404), .B1(n_408), .B2(n_409), .C(n_133), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_430), .A2(n_409), .B1(n_407), .B2(n_350), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_418), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_416), .A2(n_409), .B1(n_320), .B2(n_319), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_420), .A2(n_380), .B(n_250), .C(n_105), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_435), .B(n_391), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_439), .A2(n_389), .B(n_355), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_435), .B(n_391), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_432), .B(n_391), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_438), .A2(n_383), .B(n_385), .Y(n_451) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_426), .A2(n_122), .B(n_140), .C(n_133), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_439), .A2(n_389), .B(n_355), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_416), .B(n_166), .C(n_140), .Y(n_454) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_436), .B(n_106), .C(n_359), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_427), .A2(n_124), .B(n_133), .C(n_139), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_420), .A2(n_139), .B1(n_319), .B2(n_350), .C(n_320), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_415), .A2(n_350), .B1(n_320), .B2(n_391), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_415), .B(n_139), .C(n_204), .D(n_203), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_333), .B1(n_166), .B2(n_347), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_438), .A2(n_402), .B(n_385), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_417), .A2(n_166), .B(n_151), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_414), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_414), .B(n_377), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_424), .A2(n_333), .B1(n_166), .B2(n_347), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_433), .B(n_151), .C(n_149), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_429), .A2(n_375), .B1(n_402), .B2(n_377), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_432), .B(n_149), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_431), .A2(n_423), .B(n_425), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_421), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_410), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_429), .B(n_377), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_422), .A2(n_196), .B1(n_375), .B2(n_385), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_475), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_444), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_444), .B(n_410), .Y(n_479) );
OAI31xp33_ASAP7_75t_SL g480 ( .A1(n_465), .A2(n_423), .A3(n_431), .B(n_428), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_467), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_473), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_473), .B(n_410), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_463), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_462), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_462), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_472), .A2(n_410), .B1(n_428), .B2(n_375), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_443), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_452), .B(n_437), .C(n_434), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_466), .Y(n_490) );
OAI31xp33_ASAP7_75t_L g491 ( .A1(n_456), .A2(n_295), .A3(n_283), .B(n_289), .Y(n_491) );
NOR2x1_ASAP7_75t_L g492 ( .A(n_467), .B(n_428), .Y(n_492) );
NAND2x1p5_ASAP7_75t_SL g493 ( .A(n_471), .B(n_402), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_466), .B(n_14), .Y(n_494) );
OAI21x1_ASAP7_75t_L g495 ( .A1(n_448), .A2(n_413), .B(n_362), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_463), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_474), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_467), .B(n_375), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_14), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_457), .B(n_15), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_440), .B(n_16), .C(n_17), .D(n_18), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_474), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_463), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_451), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_455), .B(n_219), .C(n_239), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_475), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_457), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_447), .Y(n_509) );
NAND3xp33_ASAP7_75t_SL g510 ( .A(n_445), .B(n_16), .C(n_17), .Y(n_510) );
AND2x2_ASAP7_75t_SL g511 ( .A(n_471), .B(n_375), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_449), .B(n_18), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_451), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_450), .B(n_19), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_453), .B(n_321), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_450), .B(n_454), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_451), .B(n_20), .Y(n_517) );
OAI33xp33_ASAP7_75t_L g518 ( .A1(n_442), .A2(n_20), .A3(n_216), .B1(n_237), .B2(n_191), .B3(n_194), .Y(n_518) );
OAI33xp33_ASAP7_75t_L g519 ( .A1(n_460), .A2(n_237), .A3(n_194), .B1(n_202), .B2(n_216), .B3(n_211), .Y(n_519) );
OAI221xp5_ASAP7_75t_SL g520 ( .A1(n_441), .A2(n_314), .B1(n_289), .B2(n_295), .C(n_211), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_446), .A2(n_269), .A3(n_347), .B(n_360), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_459), .B(n_333), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_446), .B(n_344), .Y(n_523) );
OAI33xp33_ASAP7_75t_L g524 ( .A1(n_470), .A2(n_204), .A3(n_203), .B1(n_202), .B2(n_253), .B3(n_301), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_476), .B(n_196), .Y(n_525) );
OAI33xp33_ASAP7_75t_L g526 ( .A1(n_464), .A2(n_253), .A3(n_292), .B1(n_301), .B2(n_37), .B3(n_45), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_461), .B(n_196), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_479), .B(n_230), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_506), .B(n_458), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_484), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_479), .B(n_239), .Y(n_532) );
AOI221xp5_ASAP7_75t_L g533 ( .A1(n_501), .A2(n_468), .B1(n_239), .B2(n_230), .C(n_219), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_483), .B(n_239), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_477), .B(n_219), .Y(n_535) );
OAI21xp33_ASAP7_75t_SL g536 ( .A1(n_480), .A2(n_333), .B(n_361), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_510), .B(n_220), .C(n_242), .D(n_292), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_483), .B(n_230), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_478), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_507), .B(n_230), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_481), .Y(n_542) );
NAND5xp2_ASAP7_75t_L g543 ( .A(n_491), .B(n_25), .C(n_26), .D(n_29), .E(n_48), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_478), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_482), .B(n_219), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_482), .B(n_50), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_497), .B(n_51), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_497), .B(n_53), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_502), .B(n_362), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_508), .B(n_346), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_506), .A2(n_346), .B1(n_361), .B2(n_357), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_485), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_502), .B(n_481), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_514), .B(n_58), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_496), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_486), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_490), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_488), .B(n_59), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_508), .B(n_344), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_481), .B(n_61), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_481), .B(n_62), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_517), .B(n_312), .C(n_361), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_511), .B(n_64), .Y(n_567) );
OAI31xp33_ASAP7_75t_L g568 ( .A1(n_514), .A2(n_370), .A3(n_360), .B(n_242), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_494), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_493), .B(n_509), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_511), .B(n_67), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_493), .B(n_69), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g573 ( .A(n_489), .B(n_220), .C(n_370), .D(n_360), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_503), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_494), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_511), .B(n_70), .Y(n_576) );
INVx5_ASAP7_75t_L g577 ( .A(n_517), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_499), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_500), .B(n_356), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_503), .B(n_73), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_504), .B(n_74), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_493), .B(n_81), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_499), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_321), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_509), .B(n_321), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_500), .B(n_356), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_512), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_512), .B(n_370), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_492), .B(n_356), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_587), .B(n_492), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_555), .B(n_548), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
OAI21xp33_ASAP7_75t_L g593 ( .A1(n_536), .A2(n_487), .B(n_489), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_543), .B(n_518), .C(n_519), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_578), .B(n_523), .Y(n_595) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_556), .A2(n_521), .B(n_491), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_570), .B(n_498), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_555), .B(n_513), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_544), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_548), .B(n_513), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_548), .B(n_505), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_515), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_563), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_531), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_560), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_572), .A2(n_522), .B(n_516), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_577), .B(n_525), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_550), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_542), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_558), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_559), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g615 ( .A(n_533), .B(n_521), .C(n_520), .D(n_527), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_529), .B(n_515), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_564), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_573), .B(n_526), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_532), .B(n_515), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_583), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_553), .A2(n_524), .B(n_525), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_569), .B(n_515), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_498), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_541), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_575), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_551), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_534), .B(n_523), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_530), .A2(n_527), .B(n_495), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_531), .B(n_498), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_534), .B(n_498), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_540), .B(n_523), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_540), .B(n_523), .Y(n_632) );
NOR2xp67_ASAP7_75t_SL g633 ( .A(n_561), .B(n_528), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_551), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_538), .B(n_495), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_538), .B(n_528), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_557), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_557), .B(n_357), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_574), .B(n_357), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_542), .B(n_312), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_577), .B(n_355), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_577), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_577), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_626), .B(n_574), .Y(n_644) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_596), .B(n_568), .C(n_576), .D(n_567), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_620), .B(n_572), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_634), .B(n_545), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_625), .B(n_545), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_594), .A2(n_537), .B(n_566), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_595), .B(n_535), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_591), .B(n_577), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_592), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_612), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_591), .B(n_584), .Y(n_654) );
OAI321xp33_ASAP7_75t_L g655 ( .A1(n_628), .A2(n_567), .A3(n_571), .B1(n_576), .B2(n_582), .C(n_565), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_597), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_599), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_610), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_611), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_609), .A2(n_582), .B(n_571), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_613), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_614), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_590), .B(n_588), .Y(n_663) );
AO22x1_ASAP7_75t_L g664 ( .A1(n_642), .A2(n_563), .B1(n_565), .B2(n_547), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_602), .B(n_584), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_608), .B(n_547), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_602), .B(n_616), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_605), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_624), .B(n_549), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_622), .B(n_546), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_618), .A2(n_561), .B(n_546), .C(n_549), .Y(n_671) );
NOR2xp67_ASAP7_75t_L g672 ( .A(n_642), .B(n_581), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_598), .B(n_585), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_627), .B(n_586), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_637), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_617), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_622), .B(n_579), .Y(n_677) );
AND2x2_ASAP7_75t_SL g678 ( .A(n_609), .B(n_581), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_604), .B(n_580), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_606), .B(n_580), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_641), .A2(n_562), .B(n_552), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_637), .Y(n_682) );
AO22x1_ASAP7_75t_L g683 ( .A1(n_643), .A2(n_589), .B1(n_326), .B2(n_360), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_600), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_618), .A2(n_589), .B1(n_370), .B2(n_355), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_600), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_601), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_601), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_631), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_632), .Y(n_690) );
XNOR2x2_ASAP7_75t_L g691 ( .A(n_615), .B(n_589), .Y(n_691) );
XNOR2x1_ASAP7_75t_L g692 ( .A(n_603), .B(n_326), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_593), .B(n_326), .C(n_246), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_629), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_607), .A2(n_246), .B1(n_326), .B2(n_633), .C(n_635), .Y(n_695) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_641), .B(n_326), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_623), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_616), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_619), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_619), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_623), .B(n_246), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_621), .A2(n_636), .B1(n_635), .B2(n_630), .C(n_640), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_630), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_620), .B(n_625), .Y(n_704) );
CKINVDCx16_ASAP7_75t_R g705 ( .A(n_656), .Y(n_705) );
AOI22xp5_ASAP7_75t_SL g706 ( .A1(n_664), .A2(n_660), .B1(n_697), .B2(n_653), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_645), .A2(n_702), .B1(n_663), .B2(n_703), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_663), .A2(n_703), .B1(n_649), .B2(n_670), .Y(n_708) );
NOR2xp33_ASAP7_75t_R g709 ( .A(n_678), .B(n_691), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_657), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_686), .B(n_668), .Y(n_711) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_693), .B(n_671), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_671), .A2(n_653), .B1(n_695), .B2(n_668), .C(n_677), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_704), .B(n_698), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_694), .B(n_667), .Y(n_715) );
INVxp33_ASAP7_75t_SL g716 ( .A(n_694), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_686), .B(n_700), .Y(n_717) );
XNOR2xp5_ASAP7_75t_L g718 ( .A(n_692), .B(n_678), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g719 ( .A1(n_692), .A2(n_670), .B(n_685), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_713), .B(n_655), .C(n_683), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_707), .A2(n_704), .B1(n_646), .B2(n_676), .C(n_662), .Y(n_721) );
XNOR2xp5_ASAP7_75t_L g722 ( .A(n_706), .B(n_659), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_711), .Y(n_723) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_709), .A2(n_646), .B(n_689), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_716), .A2(n_658), .B1(n_661), .B2(n_652), .C(n_690), .Y(n_725) );
OAI211xp5_ASAP7_75t_SL g726 ( .A1(n_708), .A2(n_669), .B(n_666), .C(n_699), .Y(n_726) );
NAND4xp75_ASAP7_75t_L g727 ( .A(n_712), .B(n_672), .C(n_651), .D(n_701), .Y(n_727) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_719), .B(n_681), .C(n_673), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_705), .B1(n_719), .B2(n_710), .C(n_714), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g730 ( .A1(n_720), .A2(n_718), .B(n_715), .Y(n_730) );
OAI22x1_ASAP7_75t_L g731 ( .A1(n_722), .A2(n_717), .B1(n_687), .B2(n_688), .Y(n_731) );
AOI211xp5_ASAP7_75t_L g732 ( .A1(n_724), .A2(n_650), .B(n_674), .C(n_648), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_721), .A2(n_684), .B1(n_687), .B2(n_647), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_733), .B(n_723), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_732), .Y(n_735) );
NOR3xp33_ASAP7_75t_L g736 ( .A(n_729), .B(n_730), .C(n_727), .Y(n_736) );
OR3x1_ASAP7_75t_L g737 ( .A(n_735), .B(n_726), .C(n_731), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_734), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_738), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_737), .B(n_736), .Y(n_740) );
AOI222xp33_ASAP7_75t_L g741 ( .A1(n_739), .A2(n_725), .B1(n_696), .B2(n_682), .C1(n_675), .C2(n_644), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_741), .B(n_740), .C(n_680), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_742), .A2(n_675), .B1(n_679), .B2(n_654), .C(n_665), .Y(n_743) );
endmodule