module fake_jpeg_16259_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

AND2x4_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_42),
.B1(n_20),
.B2(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_35),
.B1(n_27),
.B2(n_18),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_28),
.B(n_19),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_35),
.B1(n_27),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_56),
.B1(n_68),
.B2(n_74),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_71),
.Y(n_109)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_35),
.B1(n_24),
.B2(n_22),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_21),
.B(n_31),
.C(n_32),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_20),
.B(n_23),
.Y(n_104)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_51),
.B1(n_21),
.B2(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_83),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_79),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_47),
.B1(n_51),
.B2(n_48),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_62),
.B1(n_45),
.B2(n_26),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_39),
.B(n_50),
.C(n_38),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_82),
.B(n_85),
.C(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_89),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_37),
.C(n_40),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_96),
.B1(n_98),
.B2(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_39),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_91),
.B(n_84),
.Y(n_140)
);

OAI211xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_42),
.B(n_29),
.C(n_30),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_42),
.B1(n_32),
.B2(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_62),
.B1(n_12),
.B2(n_13),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_61),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_48),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_1),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_2),
.Y(n_115)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_19),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_48),
.B(n_45),
.C(n_23),
.Y(n_117)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_75),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_138),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_121),
.B1(n_133),
.B2(n_96),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_129),
.B1(n_81),
.B2(n_78),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_69),
.B1(n_73),
.B2(n_62),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_72),
.B1(n_63),
.B2(n_53),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_137),
.B1(n_81),
.B2(n_107),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_51),
.B(n_48),
.C(n_45),
.Y(n_128)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_44),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_76),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_140),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_136),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_26),
.B1(n_44),
.B2(n_28),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_19),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_108),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_99),
.C(n_80),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_152),
.C(n_162),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

AOI31xp33_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_82),
.A3(n_104),
.B(n_101),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_130),
.B(n_122),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_149),
.B(n_168),
.Y(n_182)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_148),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_90),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_108),
.B1(n_95),
.B2(n_103),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_95),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_106),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_97),
.B1(n_77),
.B2(n_102),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_87),
.B1(n_86),
.B2(n_44),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_86),
.B1(n_15),
.B2(n_13),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_165),
.B1(n_168),
.B2(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_19),
.C(n_28),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_28),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_139),
.C(n_136),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_138),
.B1(n_125),
.B2(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_117),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_19),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_132),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_36),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_174),
.B(n_191),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_117),
.B1(n_115),
.B2(n_127),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_176),
.B1(n_186),
.B2(n_187),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_117),
.B1(n_115),
.B2(n_128),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_177),
.B(n_179),
.C(n_181),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_137),
.C(n_119),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_135),
.C(n_129),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_7),
.B(n_8),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_185),
.B(n_9),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_164),
.B1(n_146),
.B2(n_149),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_117),
.B1(n_124),
.B2(n_114),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_124),
.B(n_114),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_195),
.B(n_7),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_112),
.B1(n_113),
.B2(n_122),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_207),
.B1(n_176),
.B2(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_26),
.B1(n_79),
.B2(n_25),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_205),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_26),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_145),
.A2(n_156),
.B(n_161),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_201),
.B(n_204),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_79),
.B(n_25),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_172),
.A2(n_25),
.B(n_36),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_36),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_216),
.B(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_144),
.B1(n_160),
.B2(n_153),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_235),
.B1(n_175),
.B2(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_221),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_188),
.B1(n_184),
.B2(n_185),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_173),
.B(n_162),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_189),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_226),
.B(n_188),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_195),
.A2(n_7),
.B(n_8),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_230),
.B1(n_198),
.B2(n_192),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_234),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_10),
.B1(n_11),
.B2(n_181),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_173),
.C(n_177),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_251),
.C(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_250),
.B(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_258),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_214),
.A2(n_182),
.B1(n_194),
.B2(n_184),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_179),
.C(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_223),
.Y(n_280)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_200),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_211),
.A2(n_194),
.B1(n_174),
.B2(n_178),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_205),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_201),
.B1(n_196),
.B2(n_204),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_10),
.C(n_11),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_231),
.C(n_233),
.Y(n_285)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_209),
.B1(n_228),
.B2(n_210),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_228),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_222),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_270),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_222),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_262),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_240),
.B(n_241),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_284),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_225),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_258),
.B(n_239),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_223),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_220),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_248),
.C(n_252),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_242),
.B(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_285),
.B(n_260),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_287),
.B(n_221),
.Y(n_316)
);

OAI321xp33_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_249),
.A3(n_252),
.B1(n_244),
.B2(n_238),
.C(n_248),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_299),
.B(n_224),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_294),
.C(n_301),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_253),
.C(n_247),
.Y(n_294)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_303),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_238),
.B1(n_247),
.B2(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_271),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_273),
.A2(n_208),
.B(n_216),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_269),
.A2(n_274),
.B(n_282),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_267),
.B(n_285),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_227),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_230),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_280),
.B(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_264),
.C(n_283),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_315),
.C(n_289),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_308),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_317),
.B1(n_292),
.B2(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_290),
.B(n_229),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_288),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_284),
.B(n_277),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_316),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_224),
.B(n_234),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_321),
.B(n_322),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_234),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_289),
.C(n_288),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_327),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_325),
.B(n_326),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_286),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_312),
.B(n_286),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_311),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_319),
.B(n_324),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_331),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_338),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_319),
.B(n_316),
.Y(n_336)
);

AOI31xp33_ASAP7_75t_L g341 ( 
.A1(n_336),
.A2(n_328),
.A3(n_306),
.B(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_305),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_314),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_339),
.B(n_321),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_341),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_334),
.A2(n_306),
.B(n_323),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_342),
.A2(n_337),
.B(n_336),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_345),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_332),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_340),
.B(n_343),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_347),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_346),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_335),
.Y(n_353)
);


endmodule