module fake_ariane_706_n_551 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_551);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_551;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_261;
wire n_220;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_528;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_518;
wire n_439;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_511;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_451;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_234;
wire n_492;
wire n_280;
wire n_252;
wire n_215;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_540;
wire n_216;
wire n_544;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_509;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_506;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_531;

INVx1_ASAP7_75t_L g157 ( 
.A(n_31),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_26),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_141),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_20),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_37),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_54),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_50),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_3),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_90),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_14),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_11),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_35),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_4),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_58),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_122),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_45),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_124),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_92),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_13),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_49),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_64),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_80),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_133),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_8),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_18),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_10),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_39),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_139),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_129),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_113),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_93),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_38),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_72),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_33),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_99),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_118),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_108),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_21),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_96),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_94),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_114),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_24),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_30),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

BUFx8_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_219),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_169),
.B(n_221),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_162),
.B(n_0),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g254 ( 
.A1(n_157),
.A2(n_0),
.B(n_2),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_158),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_165),
.B(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_166),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_171),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_172),
.B(n_5),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_187),
.B(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_6),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_182),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_163),
.B(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_227),
.Y(n_274)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_12),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_189),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_180),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

AO21x2_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_207),
.B(n_161),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_192),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_180),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_206),
.C(n_228),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_265),
.B(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_252),
.B(n_233),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_159),
.B1(n_183),
.B2(n_185),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_252),
.B(n_194),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_273),
.B(n_213),
.Y(n_302)
);

AND2x6_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_195),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

NOR2x1p5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_161),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_258),
.A2(n_190),
.B1(n_185),
.B2(n_201),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_212),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_190),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_237),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_196),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_260),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_264),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_264),
.C(n_268),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_268),
.B1(n_254),
.B2(n_248),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_241),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_303),
.A2(n_248),
.B1(n_276),
.B2(n_197),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_275),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_197),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_288),
.B(n_167),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_199),
.Y(n_334)
);

NAND2x1p5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_201),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_202),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_316),
.B(n_170),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_303),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_207),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_236),
.B(n_234),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_275),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_276),
.B1(n_238),
.B2(n_232),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_275),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_275),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_285),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_231),
.B(n_230),
.C(n_226),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_286),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_203),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_289),
.A2(n_214),
.B(n_225),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

OR2x6_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_280),
.Y(n_365)
);

O2A1O1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_358),
.A2(n_291),
.B(n_302),
.C(n_223),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_354),
.A2(n_363),
.B(n_360),
.C(n_322),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_336),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_323),
.B(n_304),
.Y(n_374)
);

NOR2x1p5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_175),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_312),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_7),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_319),
.A2(n_215),
.B(n_208),
.C(n_209),
.Y(n_379)
);

BUFx4f_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_349),
.A2(n_222),
.B1(n_224),
.B2(n_229),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_181),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_344),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_321),
.A2(n_220),
.B(n_216),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

O2A1O1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_355),
.A2(n_331),
.B(n_330),
.C(n_362),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

BUFx2_ASAP7_75t_SL g390 ( 
.A(n_332),
.Y(n_390)
);

OR2x6_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_298),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_198),
.B(n_210),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_298),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_191),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_342),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_339),
.B(n_200),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

O2A1O1Ixp5_ASAP7_75t_SL g399 ( 
.A1(n_343),
.A2(n_298),
.B(n_9),
.C(n_8),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_9),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_326),
.B(n_15),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_335),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_16),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_338),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_399),
.A2(n_347),
.B(n_342),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_388),
.A2(n_324),
.B(n_350),
.C(n_351),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_370),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_392),
.A2(n_351),
.B(n_348),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_364),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_329),
.B(n_359),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

NAND2x1p5_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_359),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_393),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

OAI221xp5_ASAP7_75t_L g421 ( 
.A1(n_381),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.C(n_32),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_404),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_42),
.B(n_43),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_379),
.A2(n_44),
.B(n_46),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_382),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_373),
.A2(n_47),
.B(n_51),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_365),
.B(n_52),
.Y(n_427)
);

AO21x2_ASAP7_75t_L g428 ( 
.A1(n_396),
.A2(n_406),
.B(n_394),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_397),
.B(n_386),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_53),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_378),
.B(n_55),
.Y(n_431)
);

AOI222xp33_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.C1(n_61),
.C2(n_62),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_366),
.A2(n_63),
.B(n_66),
.C(n_67),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_68),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_383),
.A2(n_374),
.B(n_376),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_391),
.B1(n_400),
.B2(n_403),
.Y(n_440)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_414),
.A2(n_384),
.B(n_387),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_377),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_376),
.Y(n_443)
);

OAI221xp5_ASAP7_75t_SL g444 ( 
.A1(n_432),
.A2(n_390),
.B1(n_398),
.B2(n_371),
.C(n_389),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_424),
.A2(n_390),
.B(n_398),
.C(n_389),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_71),
.B(n_73),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_74),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_75),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_435),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_411),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_85),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_432),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_426),
.A2(n_91),
.B(n_97),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_98),
.C(n_101),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_L g455 ( 
.A1(n_421),
.A2(n_425),
.B1(n_437),
.B2(n_436),
.Y(n_455)
);

OAI211xp5_ASAP7_75t_SL g456 ( 
.A1(n_420),
.A2(n_102),
.B(n_103),
.C(n_104),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_105),
.B1(n_106),
.B2(n_111),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_423),
.A2(n_112),
.B(n_120),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_434),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_434),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_415),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_412),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_459),
.Y(n_466)
);

BUFx2_ASAP7_75t_SL g467 ( 
.A(n_450),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_451),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_408),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_412),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_438),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_R g474 ( 
.A(n_460),
.B(n_415),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_417),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_417),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_430),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_429),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_465),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_463),
.Y(n_482)
);

OAI211xp5_ASAP7_75t_L g483 ( 
.A1(n_470),
.A2(n_444),
.B(n_468),
.C(n_421),
.Y(n_483)
);

OAI31xp33_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_454),
.A3(n_456),
.B(n_422),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_419),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_419),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_470),
.A2(n_428),
.B(n_429),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_419),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_430),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_438),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_407),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_473),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_407),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_428),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_476),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_474),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_484),
.B(n_433),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_446),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_458),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_453),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_127),
.Y(n_507)
);

BUFx12f_ASAP7_75t_L g508 ( 
.A(n_479),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_131),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_135),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_138),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_491),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_140),
.Y(n_513)
);

AOI211x1_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_456),
.B(n_144),
.C(n_150),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_503),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_503),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_490),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_479),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_512),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_480),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_504),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_516),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_517),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_525),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_523),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_524),
.B(n_522),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_522),
.Y(n_530)
);

NOR4xp25_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_483),
.C(n_518),
.D(n_510),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_532),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_521),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_530),
.A2(n_501),
.B(n_519),
.C(n_507),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_506),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_534),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_535),
.Y(n_538)
);

OR4x2_ASAP7_75t_L g539 ( 
.A(n_537),
.B(n_538),
.C(n_536),
.D(n_501),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_536),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_540),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_539),
.A2(n_511),
.B1(n_490),
.B2(n_526),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_540),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_541),
.A2(n_504),
.B(n_502),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_543),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_542),
.B1(n_514),
.B2(n_502),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_544),
.A2(n_506),
.B1(n_508),
.B2(n_509),
.Y(n_547)
);

OAI221xp5_ASAP7_75t_L g548 ( 
.A1(n_546),
.A2(n_488),
.B1(n_480),
.B2(n_509),
.C(n_482),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_547),
.A2(n_482),
.B1(n_488),
.B2(n_153),
.Y(n_549)
);

NAND2x1_ASAP7_75t_SL g550 ( 
.A(n_549),
.B(n_142),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_548),
.B1(n_155),
.B2(n_156),
.Y(n_551)
);


endmodule