module fake_jpeg_2183_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_63),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_65),
.B(n_66),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_32),
.B(n_15),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g204 ( 
.A(n_67),
.Y(n_204)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_76),
.Y(n_158)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_90),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_89),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_94),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_29),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_96),
.Y(n_170)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_100),
.Y(n_150)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_101),
.Y(n_215)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_27),
.B(n_1),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_23),
.B(n_1),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_118),
.Y(n_173)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_27),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

BUFx12f_ASAP7_75t_SL g123 ( 
.A(n_31),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_52),
.B(n_48),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_124),
.B(n_125),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_30),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_59),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_35),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_26),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_33),
.B(n_14),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_48),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_133),
.Y(n_243)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_59),
.B1(n_56),
.B2(n_55),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_151),
.A2(n_189),
.B1(n_6),
.B2(n_10),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_153),
.A2(n_206),
.B(n_53),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_166),
.B(n_172),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_96),
.B(n_52),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_180),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_41),
.Y(n_182)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_81),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_117),
.A2(n_35),
.B1(n_56),
.B2(n_55),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_100),
.B(n_41),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_60),
.C(n_72),
.Y(n_228)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_61),
.B(n_43),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_42),
.Y(n_238)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_77),
.Y(n_205)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_84),
.A2(n_56),
.B1(n_55),
.B2(n_49),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_62),
.Y(n_207)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_70),
.Y(n_208)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_83),
.B(n_58),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_213),
.B(n_217),
.Y(n_274)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_93),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_219),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_79),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_222),
.B(n_223),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_43),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_224),
.A2(n_232),
.B1(n_233),
.B2(n_255),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_173),
.A2(n_126),
.B1(n_122),
.B2(n_113),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_226),
.A2(n_231),
.B1(n_266),
.B2(n_206),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_228),
.B(n_218),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_164),
.A2(n_111),
.B1(n_98),
.B2(n_104),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_49),
.B1(n_53),
.B2(n_50),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_49),
.B1(n_50),
.B2(n_42),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_155),
.B(n_39),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_234),
.B(n_237),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_235),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_155),
.B(n_39),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_238),
.B(n_247),
.Y(n_319)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_171),
.Y(n_239)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_131),
.Y(n_241)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_150),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_242),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_133),
.B(n_82),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_245),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_158),
.B(n_139),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_248),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_68),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_250),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_158),
.B(n_121),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_251),
.B(n_267),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_144),
.B(n_33),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_258),
.Y(n_326)
);

CKINVDCx9p33_ASAP7_75t_R g254 ( 
.A(n_204),
.Y(n_254)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_38),
.B1(n_58),
.B2(n_99),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_256),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_145),
.B(n_121),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_160),
.B(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_259),
.B(n_263),
.Y(n_342)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_260),
.Y(n_352)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_163),
.B(n_3),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_156),
.B(n_101),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_162),
.Y(n_265)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_151),
.A2(n_97),
.B1(n_69),
.B2(n_115),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_138),
.B(n_4),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_175),
.A2(n_89),
.B1(n_103),
.B2(n_99),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_268),
.A2(n_269),
.B1(n_292),
.B2(n_156),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_167),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_184),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_270),
.A2(n_291),
.B1(n_181),
.B2(n_171),
.Y(n_337)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_272),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_162),
.Y(n_275)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_146),
.Y(n_281)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_169),
.Y(n_282)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

CKINVDCx9p33_ASAP7_75t_R g283 ( 
.A(n_204),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_137),
.Y(n_285)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_165),
.Y(n_287)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

BUFx12_ASAP7_75t_L g288 ( 
.A(n_152),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_288),
.Y(n_299)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_159),
.Y(n_289)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_132),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_165),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_293),
.B(n_141),
.Y(n_345)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_170),
.Y(n_294)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_169),
.Y(n_295)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_303),
.Y(n_363)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_219),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_300),
.B(n_322),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_225),
.B(n_154),
.C(n_135),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_301),
.B(n_318),
.C(n_331),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_286),
.A2(n_193),
.B1(n_161),
.B2(n_179),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_149),
.B1(n_253),
.B2(n_242),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_305),
.A2(n_316),
.B1(n_324),
.B2(n_353),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_266),
.A2(n_147),
.B1(n_190),
.B2(n_186),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_148),
.C(n_140),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_218),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_245),
.A2(n_218),
.B1(n_178),
.B2(n_137),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_244),
.B(n_141),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_344),
.Y(n_376)
);

OA22x2_ASAP7_75t_L g330 ( 
.A1(n_270),
.A2(n_210),
.B1(n_181),
.B2(n_196),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_337),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_249),
.B(n_211),
.C(n_185),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_251),
.A2(n_291),
.B1(n_210),
.B2(n_196),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_239),
.B1(n_240),
.B2(n_275),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_271),
.B(n_141),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_345),
.B(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_280),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_262),
.A2(n_186),
.B1(n_176),
.B2(n_183),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_347),
.Y(n_355)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_229),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_362),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_326),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_394),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_268),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_358),
.B(n_398),
.Y(n_411)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_347),
.Y(n_359)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_349),
.B(n_318),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_360),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_221),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_366),
.A2(n_378),
.B1(n_383),
.B2(n_391),
.Y(n_407)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_368),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_183),
.B1(n_279),
.B2(n_176),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_370),
.A2(n_392),
.B1(n_395),
.B2(n_307),
.Y(n_432)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_312),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_371),
.Y(n_423)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_385),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_298),
.A2(n_256),
.B1(n_282),
.B2(n_295),
.Y(n_378)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_297),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_379),
.Y(n_404)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_315),
.A2(n_235),
.B1(n_250),
.B2(n_265),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_310),
.B(n_277),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_384),
.B(n_393),
.Y(n_427)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_220),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_346),
.Y(n_429)
);

OR2x2_ASAP7_75t_SL g387 ( 
.A(n_331),
.B(n_272),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_387),
.A2(n_304),
.B(n_152),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_264),
.C(n_257),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_389),
.C(n_390),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_241),
.C(n_280),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_320),
.B(n_284),
.C(n_261),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_309),
.A2(n_269),
.B1(n_209),
.B2(n_134),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_330),
.A2(n_260),
.B1(n_253),
.B2(n_191),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_319),
.B(n_313),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_306),
.B(n_299),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_330),
.A2(n_294),
.B1(n_236),
.B2(n_281),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_323),
.B(n_273),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_400),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_325),
.B(n_273),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_325),
.B(n_311),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_346),
.C(n_308),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_248),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_363),
.A2(n_341),
.B(n_350),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_402),
.A2(n_406),
.B(n_418),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_SL g406 ( 
.A1(n_363),
.A2(n_341),
.B(n_330),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_329),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_413),
.B(n_420),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_363),
.A2(n_340),
.B1(n_332),
.B2(n_317),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_414),
.A2(n_419),
.B1(n_432),
.B2(n_395),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_381),
.A2(n_350),
.B(n_338),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_374),
.A2(n_340),
.B1(n_332),
.B2(n_317),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_329),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_365),
.Y(n_422)
);

INVx13_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_358),
.A2(n_308),
.B(n_352),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_424),
.A2(n_391),
.B(n_390),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_386),
.B(n_352),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_429),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_439),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_362),
.B(n_307),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_433),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_296),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_374),
.A2(n_296),
.B1(n_314),
.B2(n_321),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_370),
.B1(n_361),
.B2(n_377),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_382),
.B(n_321),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_437),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_373),
.B(n_285),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_373),
.C(n_387),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_447),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_436),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_445),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_436),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_436),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_465),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_360),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_449),
.A2(n_439),
.B(n_421),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_360),
.C(n_388),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_455),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_424),
.A2(n_374),
.B1(n_366),
.B2(n_392),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_451),
.A2(n_453),
.B1(n_459),
.B2(n_469),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_375),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_454),
.B(n_460),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_356),
.Y(n_455)
);

INVx13_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_457),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_458),
.A2(n_473),
.B1(n_419),
.B2(n_428),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_378),
.B1(n_383),
.B2(n_389),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_376),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_412),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_461),
.B(n_464),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_430),
.C(n_433),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_402),
.Y(n_500)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_401),
.B(n_364),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_413),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_407),
.A2(n_380),
.B1(n_371),
.B2(n_314),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_359),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_471),
.B(n_474),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_420),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_429),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_407),
.A2(n_367),
.B1(n_372),
.B2(n_355),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_418),
.B(n_227),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_409),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_476),
.B(n_505),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_478),
.A2(n_501),
.B1(n_468),
.B2(n_425),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_452),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_479),
.B(n_481),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_480),
.A2(n_416),
.B(n_410),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_440),
.Y(n_481)
);

AO22x1_ASAP7_75t_SL g487 ( 
.A1(n_451),
.A2(n_414),
.B1(n_411),
.B2(n_423),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_444),
.Y(n_522)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_489),
.Y(n_514)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_457),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_490),
.B(n_503),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_447),
.B(n_441),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_492),
.B(n_494),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_450),
.B(n_405),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_463),
.Y(n_495)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_448),
.Y(n_499)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_499),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_416),
.C(n_410),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_449),
.A2(n_411),
.B1(n_405),
.B2(n_434),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_442),
.B(n_431),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_SL g533 ( 
.A(n_502),
.B(n_456),
.C(n_426),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_453),
.A2(n_459),
.B1(n_469),
.B2(n_472),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_442),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_504),
.B(n_445),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_409),
.Y(n_505)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_508),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_477),
.A2(n_488),
.B(n_502),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_509),
.A2(n_526),
.B(n_491),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_523),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_496),
.Y(n_511)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_511),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_484),
.Y(n_513)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_513),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_493),
.A2(n_443),
.B1(n_446),
.B2(n_458),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_515),
.A2(n_518),
.B1(n_522),
.B2(n_501),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_517),
.A2(n_507),
.B1(n_489),
.B2(n_491),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_488),
.A2(n_473),
.B1(n_468),
.B2(n_444),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_462),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_531),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_483),
.B(n_423),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_529),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_475),
.B(n_404),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_527),
.B(n_534),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_483),
.B(n_408),
.C(n_422),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_524),
.C(n_521),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_435),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_477),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_408),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_537),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_542),
.B(n_555),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_531),
.B(n_492),
.C(n_500),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_550),
.C(n_554),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_536),
.B(n_480),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_SL g572 ( 
.A(n_546),
.B(n_551),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_508),
.C(n_482),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_536),
.B(n_499),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_511),
.A2(n_497),
.B1(n_478),
.B2(n_495),
.Y(n_553)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_553),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_523),
.B(n_482),
.C(n_487),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_487),
.Y(n_555)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_556),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_562),
.Y(n_577)
);

INVx13_ASAP7_75t_L g558 ( 
.A(n_519),
.Y(n_558)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_522),
.B(n_486),
.C(n_403),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_563),
.C(n_519),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_525),
.A2(n_538),
.B1(n_515),
.B2(n_532),
.Y(n_560)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_560),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_517),
.A2(n_486),
.B1(n_485),
.B2(n_456),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_518),
.B(n_470),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_561),
.A2(n_509),
.B(n_526),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_564),
.A2(n_567),
.B(n_576),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_552),
.B(n_512),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_566),
.B(n_571),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_557),
.A2(n_535),
.B(n_537),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_569),
.B(n_563),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_513),
.C(n_530),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_514),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_573),
.B(n_583),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_545),
.B(n_516),
.C(n_520),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_574),
.B(n_581),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_541),
.A2(n_533),
.B(n_485),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_539),
.B(n_466),
.Y(n_579)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_579),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_547),
.C(n_544),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_548),
.B(n_415),
.Y(n_582)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_582),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_559),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_540),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_591),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_594),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_570),
.A2(n_562),
.B1(n_543),
.B2(n_555),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_588),
.A2(n_592),
.B1(n_597),
.B2(n_598),
.Y(n_616)
);

AOI21xp33_ASAP7_75t_L g591 ( 
.A1(n_564),
.A2(n_558),
.B(n_551),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_576),
.A2(n_554),
.B1(n_540),
.B2(n_547),
.Y(n_592)
);

HB1xp67_ASAP7_75t_SL g593 ( 
.A(n_574),
.Y(n_593)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_593),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_565),
.B(n_546),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_415),
.C(n_466),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_596),
.B(n_601),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_570),
.A2(n_379),
.B1(n_227),
.B2(n_246),
.Y(n_597)
);

AOI211xp5_ASAP7_75t_L g598 ( 
.A1(n_567),
.A2(n_304),
.B(n_397),
.C(n_157),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_246),
.C(n_288),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_578),
.B(n_288),
.C(n_152),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_581),
.Y(n_610)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_586),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_608),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g605 ( 
.A1(n_600),
.A2(n_573),
.B(n_577),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_605),
.A2(n_615),
.B(n_579),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_587),
.B(n_573),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_611),
.Y(n_619)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_586),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_610),
.B(n_594),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_569),
.Y(n_611)
);

BUFx24_ASAP7_75t_SL g612 ( 
.A(n_599),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_596),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_585),
.B(n_584),
.C(n_568),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_614),
.B(n_606),
.C(n_609),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_595),
.A2(n_577),
.B(n_575),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_603),
.A2(n_588),
.B(n_580),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_620),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_614),
.A2(n_590),
.B1(n_589),
.B2(n_611),
.Y(n_620)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_621),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_622),
.B(n_625),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_624),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_613),
.B(n_597),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_601),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_627),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_572),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_625),
.B(n_622),
.C(n_619),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_11),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_619),
.B(n_606),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_630),
.B(n_635),
.Y(n_638)
);

MAJx2_ASAP7_75t_L g635 ( 
.A(n_618),
.B(n_572),
.C(n_602),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_634),
.A2(n_617),
.B(n_598),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_636),
.A2(n_637),
.B1(n_639),
.B2(n_631),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_629),
.B(n_10),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_632),
.A2(n_157),
.B(n_11),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_640),
.B(n_633),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_641),
.B(n_642),
.C(n_631),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_643),
.A2(n_638),
.B(n_157),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_11),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_645),
.A2(n_13),
.B1(n_491),
.B2(n_283),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_13),
.Y(n_647)
);


endmodule