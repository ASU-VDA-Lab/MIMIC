module fake_netlist_6_259_n_1724 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1724);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1724;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_47),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_21),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_37),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_106),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_88),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_13),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_5),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_8),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_82),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_79),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_60),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_49),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_4),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_20),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_77),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_16),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_55),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_23),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_34),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_7),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_27),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_30),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_18),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_26),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_121),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_34),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_10),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_94),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_124),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_46),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_65),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_85),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_73),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_2),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_16),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_63),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_62),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_33),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_54),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_120),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_81),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_59),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_51),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_13),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_7),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_80),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_40),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_30),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_115),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_17),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_56),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_126),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_96),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_143),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_66),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_24),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_122),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_57),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_53),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_22),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_125),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_152),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_58),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_76),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_103),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_129),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_42),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_9),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_3),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_10),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_17),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_97),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_155),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_133),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_24),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_109),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_50),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_40),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_15),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_49),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_100),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_153),
.Y(n_283)
);

BUFx8_ASAP7_75t_SL g284 ( 
.A(n_86),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_14),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_68),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_150),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_64),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_114),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_78),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_43),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_39),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_42),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_95),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_127),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_32),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_33),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_11),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_29),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_36),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_138),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_99),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_50),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_36),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_45),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_145),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_14),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_44),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_71),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_167),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_173),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_157),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_189),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_223),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_245),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_241),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_284),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_240),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_174),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_274),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_160),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_166),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_168),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_175),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_240),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_180),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_181),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_182),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_185),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_202),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_253),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_203),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_205),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_204),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_204),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_207),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_208),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_209),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_201),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_212),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_178),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_178),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_214),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_193),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_219),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_227),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_193),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_228),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_242),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_243),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_194),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_172),
.B(n_0),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_246),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_194),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_252),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_196),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_258),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_259),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_260),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_261),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_196),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_299),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_263),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_271),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_215),
.B(n_0),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_275),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_215),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_229),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_229),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_158),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_231),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_231),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_282),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_233),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_315),
.B(n_170),
.Y(n_391)
);

AND3x1_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_279),
.C(n_232),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

CKINVDCx11_ASAP7_75t_R g395 ( 
.A(n_320),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_324),
.B(n_172),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

NAND2x1p5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_233),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_346),
.B(n_186),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_283),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_331),
.B(n_170),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_186),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_226),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_323),
.B(n_267),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_R g424 ( 
.A(n_384),
.B(n_161),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_367),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_312),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_367),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_369),
.B(n_226),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_165),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_313),
.B(n_316),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_382),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_165),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_333),
.B(n_163),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_386),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_333),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_325),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_352),
.B(n_326),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_327),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_314),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_328),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_339),
.B(n_278),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_329),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_353),
.B(n_233),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_449),
.B(n_420),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_370),
.B1(n_380),
.B2(n_332),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_358),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_359),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_436),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_404),
.A2(n_352),
.B1(n_268),
.B2(n_317),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_278),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

AND2x6_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_179),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_361),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_397),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_388),
.Y(n_479)
);

AND3x2_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_218),
.C(n_350),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_434),
.A2(n_376),
.B1(n_305),
.B2(n_232),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_436),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_449),
.B(n_362),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_392),
.A2(n_356),
.B1(n_334),
.B2(n_377),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_L g488 ( 
.A(n_389),
.B(n_308),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_446),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_391),
.B(n_363),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_433),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_446),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_305),
.B1(n_297),
.B2(n_298),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_434),
.A2(n_293),
.B1(n_298),
.B2(n_297),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_455),
.B(n_366),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_389),
.B(n_308),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_449),
.B(n_179),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_449),
.B(n_371),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_404),
.A2(n_266),
.B1(n_285),
.B2(n_257),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_391),
.B(n_190),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_391),
.B(n_374),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_449),
.B(n_190),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g512 ( 
.A1(n_404),
.A2(n_216),
.B1(n_184),
.B2(n_183),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_455),
.B(n_378),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_389),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_387),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_442),
.Y(n_516)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_449),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_434),
.B(n_197),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_451),
.B(n_335),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_434),
.A2(n_279),
.B1(n_293),
.B2(n_307),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_453),
.B(n_307),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_453),
.B(n_336),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_453),
.B(n_337),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_447),
.B(n_197),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_405),
.B(n_318),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_398),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_442),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_408),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_405),
.B(n_199),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_447),
.B(n_373),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_450),
.B(n_340),
.Y(n_536)
);

BUFx4f_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx4_ASAP7_75t_SL g539 ( 
.A(n_389),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_401),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_401),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_447),
.B(n_368),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

XNOR2x2_ASAP7_75t_L g544 ( 
.A(n_441),
.B(n_188),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_401),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_450),
.B(n_311),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_408),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_447),
.B(n_348),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_454),
.B(n_164),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_454),
.B(n_349),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_401),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_406),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_390),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_454),
.B(n_319),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_406),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_439),
.B(n_198),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_406),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_454),
.B(n_288),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_402),
.B(n_289),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_404),
.B(n_198),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_410),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_404),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_439),
.B(n_206),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_406),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_410),
.A2(n_452),
.B1(n_413),
.B2(n_419),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_410),
.B(n_290),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_398),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_398),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_452),
.B(n_206),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_452),
.B(n_210),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_406),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_406),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_411),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_441),
.B(n_448),
.Y(n_580)
);

BUFx4f_ASAP7_75t_L g581 ( 
.A(n_389),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_398),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_404),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_390),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_448),
.B(n_300),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_412),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_412),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_414),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_414),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_402),
.B(n_304),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_398),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_413),
.B(n_169),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_424),
.A2(n_192),
.B1(n_309),
.B2(n_306),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_400),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_417),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_402),
.B(n_210),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_404),
.B(n_171),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_413),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_417),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_418),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_389),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_406),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_418),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_413),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_409),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_413),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_566),
.B(n_233),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_490),
.B(n_402),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_566),
.B(n_537),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_490),
.B(n_415),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_494),
.B(n_415),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_498),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_537),
.B(n_233),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_494),
.B(n_415),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_534),
.B(n_571),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_543),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_543),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_422),
.C(n_395),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_537),
.B(n_308),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_533),
.B(n_415),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_583),
.A2(n_424),
.B1(n_422),
.B2(n_159),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_491),
.Y(n_623)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_550),
.B(n_421),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_546),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_415),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_499),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_562),
.B(n_308),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_464),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_546),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_562),
.B(n_308),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_503),
.B(n_428),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_513),
.B(n_428),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_549),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_562),
.B(n_308),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_554),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_549),
.B(n_419),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_569),
.B(n_419),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_569),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_579),
.B(n_419),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_554),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_579),
.B(n_419),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_500),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_515),
.B(n_476),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_500),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_536),
.B(n_436),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_464),
.A2(n_224),
.B1(n_221),
.B2(n_220),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_SL g649 ( 
.A(n_583),
.B(n_213),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_491),
.B(n_421),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_586),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_517),
.B(n_308),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_587),
.B(n_431),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_587),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_519),
.A2(n_431),
.B1(n_222),
.B2(n_225),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_588),
.B(n_431),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_554),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_588),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_548),
.B(n_176),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_540),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_540),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_589),
.B(n_431),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_589),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_595),
.B(n_431),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_510),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_541),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_510),
.B(n_427),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_554),
.Y(n_668)
);

BUFx8_ASAP7_75t_L g669 ( 
.A(n_461),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_595),
.B(n_396),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_606),
.B(n_427),
.Y(n_671)
);

INVxp33_ASAP7_75t_SL g672 ( 
.A(n_459),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_541),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_530),
.B(n_177),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_599),
.B(n_396),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_556),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_545),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_575),
.A2(n_236),
.B1(n_287),
.B2(n_273),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_599),
.B(n_432),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_600),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_517),
.B(n_308),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_600),
.B(n_432),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_517),
.A2(n_445),
.B(n_444),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_187),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_593),
.B(n_525),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_603),
.B(n_432),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_581),
.B(n_468),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_581),
.B(n_409),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_527),
.B(n_191),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_545),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_606),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_581),
.B(n_409),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_519),
.A2(n_230),
.B1(n_213),
.B2(n_222),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_559),
.A2(n_225),
.B1(n_230),
.B2(n_244),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_468),
.B(n_409),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_603),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_547),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_479),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_547),
.B(n_435),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_479),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_575),
.A2(n_576),
.B1(n_551),
.B2(n_524),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_468),
.B(n_409),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_556),
.B(n_235),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_435),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_576),
.A2(n_239),
.B(n_303),
.C(n_296),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_598),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_553),
.A2(n_389),
.B(n_244),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_483),
.B(n_435),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_483),
.B(n_440),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_SL g710 ( 
.A(n_551),
.B(n_248),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_559),
.A2(n_568),
.B1(n_544),
.B2(n_509),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_584),
.B(n_429),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_461),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_486),
.B(n_487),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_486),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_487),
.B(n_440),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_495),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_524),
.A2(n_248),
.B1(n_250),
.B2(n_296),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_544),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_495),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_598),
.B(n_409),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_482),
.B(n_429),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_496),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_496),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_598),
.B(n_409),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_504),
.B(n_409),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_502),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_502),
.B(n_440),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_504),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_552),
.B(n_430),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_516),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_520),
.B(n_425),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_524),
.B(n_430),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_520),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_568),
.B(n_444),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_524),
.A2(n_291),
.B1(n_287),
.B2(n_262),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_521),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_526),
.B(n_444),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_509),
.B(n_437),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_526),
.B(n_425),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_532),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_532),
.Y(n_742)
);

AND2x6_ASAP7_75t_L g743 ( 
.A(n_509),
.B(n_256),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_471),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_472),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_465),
.B(n_445),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_457),
.Y(n_747)
);

AND2x2_ASAP7_75t_SL g748 ( 
.A(n_488),
.B(n_256),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_485),
.B(n_395),
.C(n_195),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_460),
.A2(n_272),
.B1(n_295),
.B2(n_291),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_457),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_467),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_597),
.A2(n_295),
.B(n_272),
.C(n_273),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_467),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_462),
.B(n_425),
.Y(n_755)
);

NOR3xp33_ASAP7_75t_L g756 ( 
.A(n_469),
.B(n_276),
.C(n_211),
.Y(n_756)
);

AND2x6_ASAP7_75t_SL g757 ( 
.A(n_557),
.B(n_262),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_480),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_567),
.B(n_425),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_465),
.B(n_445),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_567),
.B(n_425),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_529),
.B(n_389),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_529),
.A2(n_303),
.B1(n_389),
.B2(n_425),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_465),
.B(n_425),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_466),
.B(n_425),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_473),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_466),
.B(n_437),
.Y(n_767)
);

NOR2x1p5_ASAP7_75t_L g768 ( 
.A(n_564),
.B(n_200),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_596),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_470),
.B(n_438),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_484),
.A2(n_443),
.B1(n_438),
.B2(n_426),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_473),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_567),
.B(n_400),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_470),
.B(n_443),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_604),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_463),
.B(n_400),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_687),
.A2(n_522),
.B(n_475),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_644),
.B(n_769),
.Y(n_778)
);

O2A1O1Ixp5_ASAP7_75t_L g779 ( 
.A1(n_652),
.A2(n_563),
.B(n_507),
.C(n_592),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_687),
.A2(n_522),
.B(n_475),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_719),
.A2(n_505),
.B(n_488),
.C(n_458),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_685),
.A2(n_590),
.B(n_585),
.C(n_542),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_659),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_629),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_689),
.B(n_529),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_705),
.A2(n_505),
.B(n_535),
.C(n_508),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_722),
.B(n_470),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_695),
.A2(n_522),
.B(n_475),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_650),
.B(n_470),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_615),
.A2(n_481),
.B(n_497),
.C(n_501),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_701),
.A2(n_604),
.B1(n_529),
.B2(n_565),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_735),
.A2(n_529),
.B(n_489),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_623),
.B(n_665),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_676),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_624),
.B(n_512),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_706),
.B(n_523),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_695),
.A2(n_702),
.B(n_608),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_667),
.B(n_565),
.Y(n_798)
);

BUFx12f_ASAP7_75t_L g799 ( 
.A(n_669),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_684),
.A2(n_489),
.B(n_466),
.C(n_493),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_712),
.B(n_565),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_711),
.A2(n_565),
.B1(n_604),
.B2(n_489),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_632),
.B(n_217),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_702),
.A2(n_755),
.B(n_725),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_670),
.B(n_529),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_669),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_672),
.B(n_471),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_691),
.Y(n_808)
);

BUFx4f_ASAP7_75t_L g809 ( 
.A(n_703),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_721),
.A2(n_518),
.B(n_478),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_609),
.A2(n_518),
.B(n_478),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_706),
.B(n_463),
.Y(n_812)
);

BUFx24_ASAP7_75t_L g813 ( 
.A(n_669),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_609),
.A2(n_518),
.B(n_478),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_647),
.B(n_249),
.C(n_234),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_675),
.B(n_472),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_634),
.B(n_472),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_706),
.B(n_463),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_251),
.C(n_238),
.Y(n_819)
);

OAI321xp33_ASAP7_75t_L g820 ( 
.A1(n_750),
.A2(n_407),
.A3(n_416),
.B1(n_423),
.B2(n_426),
.C(n_294),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_775),
.B(n_739),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_699),
.A2(n_518),
.B(n_478),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_639),
.B(n_645),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_660),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_706),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_737),
.B(n_471),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_704),
.A2(n_518),
.B(n_478),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_674),
.B(n_471),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_748),
.A2(n_474),
.B1(n_477),
.B2(n_492),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_739),
.B(n_539),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_710),
.A2(n_474),
.B(n_477),
.C(n_492),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_661),
.A2(n_471),
.B(n_463),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_715),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_713),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_770),
.B(n_237),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_710),
.A2(n_616),
.B1(n_625),
.B2(n_617),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_661),
.A2(n_514),
.B(n_601),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_472),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_654),
.B(n_472),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_666),
.A2(n_514),
.B(n_601),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_666),
.A2(n_514),
.B(n_601),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_673),
.A2(n_514),
.B(n_601),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_768),
.B(n_493),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_764),
.A2(n_765),
.B(n_760),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_677),
.A2(n_601),
.B(n_573),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_774),
.B(n_247),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_733),
.B(n_254),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_677),
.A2(n_573),
.B(n_602),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_717),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_622),
.B(n_255),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_630),
.A2(n_511),
.B1(n_472),
.B2(n_506),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_703),
.B(n_264),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_690),
.A2(n_573),
.B(n_602),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_691),
.B(n_539),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_658),
.B(n_506),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_663),
.B(n_506),
.Y(n_857)
);

OAI321xp33_ASAP7_75t_L g858 ( 
.A1(n_753),
.A2(n_426),
.A3(n_423),
.B1(n_416),
.B2(n_407),
.C(n_281),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_690),
.A2(n_573),
.B(n_555),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_680),
.B(n_265),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_652),
.A2(n_605),
.B(n_555),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_696),
.B(n_506),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_698),
.B(n_269),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_SL g864 ( 
.A(n_745),
.B(n_573),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_SL g865 ( 
.A(n_756),
.B(n_270),
.C(n_277),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_697),
.A2(n_605),
.B(n_558),
.Y(n_866)
);

NOR2x1_ASAP7_75t_L g867 ( 
.A(n_636),
.B(n_528),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_703),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_739),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_636),
.B(n_528),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_648),
.B(n_286),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_746),
.A2(n_594),
.B(n_591),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_705),
.A2(n_423),
.B(n_407),
.C(n_416),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_671),
.B(n_539),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_671),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_671),
.A2(n_511),
.B1(n_506),
.B2(n_561),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_714),
.A2(n_570),
.B(n_558),
.C(n_560),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_697),
.A2(n_570),
.B(n_560),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_744),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_691),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_748),
.A2(n_577),
.B1(n_561),
.B2(n_578),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_717),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_720),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_620),
.A2(n_577),
.B(n_578),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_700),
.B(n_292),
.Y(n_885)
);

BUFx4f_ASAP7_75t_L g886 ( 
.A(n_743),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_727),
.B(n_301),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_757),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_753),
.A2(n_594),
.B(n_591),
.C(n_582),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_621),
.A2(n_626),
.B(n_637),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_310),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_723),
.B(n_506),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_758),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_758),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_723),
.B(n_724),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_724),
.B(n_591),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_759),
.A2(n_538),
.B(n_582),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_638),
.A2(n_511),
.B(n_594),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_636),
.B(n_539),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_759),
.A2(n_582),
.B(n_574),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_761),
.A2(n_574),
.B(n_538),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_641),
.B(n_574),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_612),
.B(n_511),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_761),
.A2(n_538),
.B(n_531),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_729),
.B(n_531),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_607),
.A2(n_531),
.B(n_528),
.C(n_511),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_773),
.A2(n_400),
.B(n_511),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_731),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_612),
.B(n_400),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_641),
.B(n_151),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_744),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_734),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_773),
.A2(n_400),
.B(n_142),
.Y(n_913)
);

CKINVDCx14_ASAP7_75t_R g914 ( 
.A(n_758),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_649),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_618),
.B(n_627),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_607),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_683),
.A2(n_400),
.B(n_141),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_619),
.B(n_6),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_613),
.A2(n_642),
.B(n_640),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_613),
.A2(n_140),
.B(n_136),
.Y(n_921)
);

CKINVDCx11_ASAP7_75t_R g922 ( 
.A(n_749),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_649),
.A2(n_6),
.B(n_11),
.C(n_12),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_653),
.A2(n_132),
.B(n_128),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_657),
.B(n_118),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_643),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_741),
.Y(n_927)
);

BUFx8_ASAP7_75t_SL g928 ( 
.A(n_643),
.Y(n_928)
);

BUFx4f_ASAP7_75t_L g929 ( 
.A(n_743),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_620),
.A2(n_113),
.B(n_112),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_657),
.B(n_111),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_656),
.A2(n_107),
.B(n_105),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_662),
.A2(n_12),
.B(n_15),
.C(n_19),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_646),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_664),
.A2(n_744),
.B(n_692),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_742),
.B(n_20),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_657),
.B(n_21),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_646),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_771),
.B(n_25),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_767),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_668),
.B(n_92),
.Y(n_941)
);

NOR2x1_ASAP7_75t_R g942 ( 
.A(n_745),
.B(n_26),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_678),
.A2(n_27),
.B(n_28),
.C(n_31),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_668),
.B(n_90),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_655),
.B(n_28),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_679),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_744),
.A2(n_692),
.B(n_688),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_682),
.A2(n_31),
.B(n_32),
.C(n_35),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_668),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_718),
.A2(n_38),
.B(n_39),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_688),
.A2(n_91),
.B(n_89),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_693),
.B(n_87),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_743),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_686),
.B(n_708),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_709),
.B(n_716),
.Y(n_955)
);

CKINVDCx6p67_ASAP7_75t_R g956 ( 
.A(n_813),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_928),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_778),
.A2(n_628),
.B(n_631),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_784),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_834),
.Y(n_960)
);

NOR3xp33_ASAP7_75t_SL g961 ( 
.A(n_865),
.B(n_628),
.C(n_631),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_783),
.B(n_694),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_803),
.B(n_728),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_920),
.A2(n_635),
.B(n_681),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_851),
.B(n_736),
.C(n_635),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_946),
.B(n_743),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_954),
.A2(n_681),
.B(n_611),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_787),
.B(n_752),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_782),
.A2(n_610),
.B(n_614),
.C(n_766),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_807),
.A2(n_763),
.B1(n_772),
.B2(n_766),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_825),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_865),
.A2(n_743),
.B1(n_772),
.B2(n_747),
.Y(n_972)
);

XOR2x2_ASAP7_75t_SL g973 ( 
.A(n_939),
.B(n_38),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_883),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_801),
.A2(n_743),
.B1(n_762),
.B2(n_738),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_874),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_789),
.B(n_754),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_798),
.B(n_754),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_869),
.B(n_875),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_955),
.A2(n_762),
.B(n_707),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_833),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_835),
.B(n_751),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_786),
.A2(n_781),
.B(n_779),
.C(n_795),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_805),
.A2(n_752),
.B(n_751),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_940),
.B(n_823),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_948),
.A2(n_740),
.B(n_732),
.C(n_726),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_847),
.B(n_726),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_891),
.B(n_740),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_786),
.A2(n_781),
.B(n_779),
.C(n_915),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_908),
.B(n_732),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_794),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_893),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_794),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_869),
.B(n_776),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_912),
.B(n_41),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_825),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_837),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_785),
.A2(n_74),
.B(n_61),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_875),
.A2(n_83),
.B1(n_43),
.B2(n_48),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_799),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_828),
.A2(n_41),
.B1(n_48),
.B2(n_51),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_806),
.Y(n_1002)
);

INVx6_ASAP7_75t_L g1003 ( 
.A(n_825),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_793),
.B(n_52),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_850),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_828),
.A2(n_52),
.B(n_53),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_819),
.B(n_919),
.C(n_815),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_927),
.B(n_826),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_915),
.A2(n_848),
.B(n_804),
.C(n_790),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_SL g1010 ( 
.A1(n_796),
.A2(n_836),
.B(n_816),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_943),
.A2(n_917),
.B(n_923),
.C(n_950),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_825),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_922),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_848),
.A2(n_797),
.B(n_885),
.C(n_860),
.Y(n_1014)
);

INVx6_ASAP7_75t_L g1015 ( 
.A(n_830),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_890),
.A2(n_792),
.B(n_935),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_860),
.B(n_863),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_895),
.A2(n_898),
.B(n_947),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_868),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_868),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_791),
.A2(n_802),
.B1(n_882),
.B2(n_929),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_894),
.Y(n_1022)
);

OR2x6_ASAP7_75t_SL g1023 ( 
.A(n_945),
.B(n_914),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_917),
.A2(n_831),
.B(n_933),
.C(n_873),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_863),
.B(n_885),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_822),
.A2(n_827),
.B(n_780),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_830),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_887),
.B(n_853),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_821),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_887),
.B(n_793),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_SL g1031 ( 
.A1(n_888),
.A2(n_821),
.B1(n_936),
.B2(n_910),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_871),
.B(n_809),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_880),
.B(n_824),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_809),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_910),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_844),
.B(n_944),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_944),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_937),
.A2(n_952),
.B1(n_874),
.B2(n_934),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_808),
.B(n_886),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_L g1040 ( 
.A(n_953),
.B(n_879),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_933),
.A2(n_873),
.B(n_877),
.C(n_820),
.Y(n_1041)
);

INVx3_ASAP7_75t_SL g1042 ( 
.A(n_953),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_879),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_926),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_938),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_777),
.A2(n_800),
.B(n_788),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_889),
.A2(n_906),
.B(n_857),
.C(n_862),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_949),
.B(n_855),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_916),
.B(n_896),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_879),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_896),
.A2(n_881),
.B(n_906),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_953),
.B(n_930),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_892),
.A2(n_849),
.B(n_854),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_949),
.A2(n_905),
.B1(n_953),
.B2(n_829),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_905),
.B(n_864),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_859),
.A2(n_811),
.B(n_814),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_909),
.A2(n_903),
.B(n_810),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_889),
.A2(n_858),
.B(n_817),
.C(n_840),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_839),
.A2(n_856),
.B(n_878),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_879),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_866),
.A2(n_900),
.B(n_897),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_884),
.A2(n_861),
.B(n_904),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_925),
.A2(n_941),
.B(n_931),
.C(n_951),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_867),
.B(n_911),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_SL g1065 ( 
.A1(n_942),
.A2(n_870),
.B1(n_876),
.B2(n_852),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_911),
.B(n_870),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_911),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_911),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_902),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_913),
.B(n_932),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_899),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_872),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_845),
.B(n_901),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_924),
.B(n_907),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_812),
.Y(n_1075)
);

INVx3_ASAP7_75t_SL g1076 ( 
.A(n_818),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_832),
.A2(n_846),
.B(n_918),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_921),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_838),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_841),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_842),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_843),
.B(n_778),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_783),
.A2(n_685),
.B1(n_580),
.B2(n_672),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_783),
.A2(n_685),
.B1(n_580),
.B2(n_672),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_783),
.A2(n_685),
.B1(n_580),
.B2(n_672),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_800),
.A2(n_613),
.B(n_785),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_778),
.A2(n_783),
.B1(n_685),
.B2(n_615),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_778),
.B(n_783),
.Y(n_1088)
);

NAND3xp33_ASAP7_75t_L g1089 ( 
.A(n_851),
.B(n_689),
.C(n_685),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_799),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_825),
.Y(n_1091)
);

AND2x2_ASAP7_75t_SL g1092 ( 
.A(n_809),
.B(n_647),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_883),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_778),
.A2(n_517),
.B(n_687),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_778),
.B(n_783),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_R g1096 ( 
.A(n_784),
.B(n_464),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1028),
.B(n_1083),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1089),
.A2(n_1017),
.B(n_1025),
.C(n_1014),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1099)
);

NAND3x1_ASAP7_75t_L g1100 ( 
.A(n_1032),
.B(n_1085),
.C(n_1084),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_984),
.A2(n_1077),
.B(n_1053),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_984),
.A2(n_1077),
.B(n_1053),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1092),
.B(n_1030),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_996),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_996),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1035),
.B(n_1029),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1043),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1026),
.A2(n_1056),
.B(n_1046),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1016),
.A2(n_1094),
.B(n_1070),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1027),
.B(n_1034),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_992),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_965),
.A2(n_963),
.B(n_1009),
.C(n_1011),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_L g1113 ( 
.A1(n_1087),
.A2(n_1011),
.B1(n_1001),
.B2(n_1004),
.C(n_1007),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_974),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_991),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1026),
.A2(n_1056),
.B(n_1046),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_985),
.B(n_982),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_983),
.A2(n_1010),
.B(n_961),
.C(n_989),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_962),
.A2(n_1041),
.B(n_958),
.C(n_1063),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_993),
.B(n_973),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1093),
.B(n_1037),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1008),
.B(n_987),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1051),
.A2(n_958),
.B(n_1047),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_1020),
.B(n_968),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_988),
.B(n_1036),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_976),
.B(n_1022),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1007),
.A2(n_1006),
.B1(n_1031),
.B2(n_999),
.C(n_1041),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1049),
.A2(n_1065),
.B1(n_981),
.B2(n_1005),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1016),
.A2(n_1073),
.A3(n_1051),
.B(n_1021),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_966),
.A2(n_1055),
.B(n_1039),
.C(n_1082),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_995),
.A2(n_979),
.B1(n_978),
.B2(n_977),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_1015),
.B(n_996),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1061),
.A2(n_1057),
.B(n_1062),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1061),
.A2(n_1057),
.B(n_1059),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_997),
.A2(n_1038),
.B1(n_975),
.B2(n_990),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1094),
.A2(n_980),
.B(n_1018),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_959),
.B(n_960),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_980),
.A2(n_1018),
.B(n_964),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1058),
.A2(n_967),
.B(n_964),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_957),
.A2(n_1019),
.B1(n_1013),
.B2(n_1000),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1054),
.A2(n_969),
.A3(n_1059),
.B(n_970),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_976),
.B(n_1033),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_SL g1143 ( 
.A(n_1042),
.B(n_1076),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1058),
.A2(n_1024),
.B(n_986),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_1006),
.A2(n_998),
.A3(n_1078),
.B(n_1080),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1063),
.A2(n_1040),
.B(n_1086),
.Y(n_1146)
);

AO21x2_ASAP7_75t_L g1147 ( 
.A1(n_1086),
.A2(n_1024),
.B(n_998),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_986),
.A2(n_1066),
.B(n_972),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1023),
.B(n_1015),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1012),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1048),
.A2(n_994),
.B(n_1044),
.Y(n_1151)
);

BUFx8_ASAP7_75t_L g1152 ( 
.A(n_1090),
.Y(n_1152)
);

AO22x2_ASAP7_75t_L g1153 ( 
.A1(n_1072),
.A2(n_1067),
.B1(n_1075),
.B2(n_1069),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1045),
.Y(n_1154)
);

AO32x2_ASAP7_75t_L g1155 ( 
.A1(n_1075),
.A2(n_1050),
.A3(n_1052),
.B1(n_1079),
.B2(n_971),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1060),
.A2(n_1081),
.B(n_1043),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1015),
.B(n_1064),
.Y(n_1157)
);

BUFx2_ASAP7_75t_R g1158 ( 
.A(n_1002),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1068),
.B(n_1064),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1012),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1012),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1071),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1071),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_956),
.B(n_1071),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1081),
.A2(n_1043),
.B(n_1050),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1003),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1091),
.B(n_1003),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1003),
.A2(n_1081),
.B1(n_1091),
.B2(n_1043),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_SL g1169 ( 
.A(n_1091),
.B(n_1096),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_R g1172 ( 
.A(n_959),
.B(n_395),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_L g1173 ( 
.A(n_1089),
.B(n_1025),
.C(n_1017),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1089),
.A2(n_1025),
.B(n_1017),
.C(n_685),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1089),
.A2(n_672),
.B1(n_647),
.B2(n_632),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_983),
.A2(n_989),
.A3(n_1016),
.B(n_1046),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1016),
.A2(n_1046),
.B(n_983),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1028),
.B(n_1083),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1089),
.B(n_1017),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_983),
.A2(n_989),
.A3(n_1016),
.B(n_1046),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1089),
.A2(n_1025),
.B(n_1017),
.C(n_685),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1087),
.Y(n_1186)
);

AOI221xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1011),
.A2(n_1025),
.B1(n_1017),
.B2(n_1001),
.C(n_950),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_983),
.A2(n_989),
.A3(n_1016),
.B(n_1046),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_992),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_983),
.A2(n_989),
.A3(n_1016),
.B(n_1046),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_991),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_991),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1196)
);

NAND3x1_ASAP7_75t_L g1197 ( 
.A(n_1032),
.B(n_647),
.C(n_619),
.Y(n_1197)
);

BUFx2_ASAP7_75t_R g1198 ( 
.A(n_959),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1035),
.B(n_1029),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_991),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1201)
);

AO32x2_ASAP7_75t_L g1202 ( 
.A1(n_1087),
.A2(n_719),
.A3(n_1021),
.B1(n_1001),
.B2(n_1065),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_991),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_974),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1205)
);

BUFx4f_ASAP7_75t_L g1206 ( 
.A(n_956),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1089),
.A2(n_1025),
.B(n_1017),
.C(n_685),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1089),
.C(n_685),
.Y(n_1208)
);

AO32x2_ASAP7_75t_L g1209 ( 
.A1(n_1087),
.A2(n_719),
.A3(n_1021),
.B1(n_1001),
.B2(n_1065),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1212)
);

AOI31xp67_ASAP7_75t_L g1213 ( 
.A1(n_1074),
.A2(n_1070),
.A3(n_1073),
.B(n_613),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1083),
.B(n_1084),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1089),
.A2(n_1025),
.B1(n_1017),
.B2(n_672),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1089),
.A2(n_1025),
.B1(n_1017),
.B2(n_672),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_991),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1089),
.C(n_685),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1089),
.B(n_1017),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_983),
.A2(n_989),
.A3(n_1016),
.B(n_1046),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1006),
.A2(n_1011),
.B(n_998),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1089),
.A2(n_1025),
.B(n_1017),
.C(n_685),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_976),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_959),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1016),
.A2(n_517),
.B(n_537),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_976),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_984),
.A2(n_872),
.B(n_1077),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_974),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1132),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1215),
.A2(n_1222),
.B1(n_1180),
.B2(n_1173),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1175),
.A2(n_1113),
.B1(n_1127),
.B2(n_1218),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1218),
.A2(n_1219),
.B1(n_1097),
.B2(n_1178),
.Y(n_1238)
);

CKINVDCx6p67_ASAP7_75t_R g1239 ( 
.A(n_1192),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1144),
.A2(n_1128),
.B1(n_1103),
.B2(n_1123),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1099),
.B(n_1181),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1114),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1191),
.B(n_1205),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1144),
.A2(n_1128),
.B1(n_1123),
.B2(n_1226),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1225),
.A2(n_1201),
.B1(n_1139),
.B2(n_1177),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1219),
.A2(n_1207),
.B1(n_1227),
.B2(n_1185),
.Y(n_1246)
);

CKINVDCx6p67_ASAP7_75t_R g1247 ( 
.A(n_1161),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1154),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1132),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1204),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1174),
.A2(n_1100),
.B1(n_1117),
.B2(n_1112),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1229),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1152),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1197),
.A2(n_1187),
.B1(n_1120),
.B2(n_1137),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1107),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1122),
.A2(n_1124),
.B1(n_1125),
.B2(n_1131),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1115),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1115),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1234),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1152),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1186),
.A2(n_1139),
.B1(n_1177),
.B2(n_1135),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1194),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1135),
.A2(n_1147),
.B1(n_1131),
.B2(n_1121),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1149),
.B(n_1159),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1126),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1142),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1132),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1111),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1098),
.A2(n_1118),
.B1(n_1221),
.B2(n_1208),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1153),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1187),
.B(n_1195),
.Y(n_1271)
);

BUFx2_ASAP7_75t_SL g1272 ( 
.A(n_1126),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1146),
.A2(n_1209),
.B1(n_1202),
.B2(n_1147),
.Y(n_1273)
);

CKINVDCx6p67_ASAP7_75t_R g1274 ( 
.A(n_1110),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1206),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1110),
.Y(n_1276)
);

OAI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1119),
.A2(n_1140),
.B(n_1200),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1169),
.A2(n_1110),
.B1(n_1209),
.B2(n_1202),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1202),
.A2(n_1209),
.B1(n_1206),
.B2(n_1148),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1143),
.Y(n_1280)
);

CKINVDCx16_ASAP7_75t_R g1281 ( 
.A(n_1159),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1164),
.A2(n_1106),
.B1(n_1199),
.B2(n_1157),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1220),
.A2(n_1109),
.B1(n_1138),
.B2(n_1228),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1167),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1168),
.A2(n_1162),
.B1(n_1163),
.B2(n_1199),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1176),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1153),
.A2(n_1198),
.B1(n_1106),
.B2(n_1107),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1232),
.A2(n_1136),
.B1(n_1166),
.B2(n_1116),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1232),
.A2(n_1108),
.B1(n_1151),
.B2(n_1190),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1130),
.A2(n_1160),
.B1(n_1104),
.B2(n_1105),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_SL g1291 ( 
.A(n_1104),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1105),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1171),
.A2(n_1179),
.B1(n_1196),
.B2(n_1210),
.Y(n_1293)
);

INVx6_ASAP7_75t_L g1294 ( 
.A(n_1105),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_1150),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1212),
.A2(n_1214),
.B1(n_1231),
.B2(n_1224),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1158),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1155),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1155),
.Y(n_1299)
);

INVx6_ASAP7_75t_L g1300 ( 
.A(n_1150),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1150),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1155),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1182),
.Y(n_1303)
);

AOI22x1_ASAP7_75t_SL g1304 ( 
.A1(n_1172),
.A2(n_1156),
.B1(n_1165),
.B2(n_1145),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1133),
.A2(n_1134),
.B1(n_1102),
.B2(n_1101),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1182),
.A2(n_1223),
.B1(n_1193),
.B2(n_1188),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1188),
.A2(n_1223),
.B1(n_1193),
.B2(n_1172),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1141),
.A2(n_1129),
.B1(n_1145),
.B2(n_1213),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1145),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1129),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1141),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1141),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1170),
.Y(n_1313)
);

BUFx4f_ASAP7_75t_L g1314 ( 
.A(n_1183),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1184),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1189),
.A2(n_1211),
.B1(n_1216),
.B2(n_1217),
.Y(n_1316)
);

CKINVDCx6p67_ASAP7_75t_R g1317 ( 
.A(n_1230),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1233),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1180),
.A2(n_1017),
.B1(n_1025),
.B2(n_672),
.Y(n_1319)
);

AO22x1_ASAP7_75t_L g1320 ( 
.A1(n_1180),
.A2(n_633),
.B1(n_632),
.B2(n_647),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1161),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1132),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1103),
.B(n_1097),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1161),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1099),
.B(n_1181),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1229),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1146),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1132),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1215),
.A2(n_1089),
.B1(n_1017),
.B2(n_1025),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1192),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1104),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1099),
.B(n_1181),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1115),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1180),
.A2(n_1017),
.B1(n_1025),
.B2(n_672),
.Y(n_1334)
);

CKINVDCx14_ASAP7_75t_R g1335 ( 
.A(n_1229),
.Y(n_1335)
);

INVx3_ASAP7_75t_SL g1336 ( 
.A(n_1229),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1180),
.A2(n_1017),
.B1(n_1025),
.B2(n_672),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1192),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1174),
.A2(n_1089),
.B(n_1025),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1175),
.A2(n_1089),
.B1(n_1084),
.B2(n_1085),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1161),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1192),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1180),
.A2(n_1025),
.B(n_1017),
.Y(n_1343)
);

BUFx8_ASAP7_75t_L g1344 ( 
.A(n_1203),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1229),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1103),
.B(n_1097),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1327),
.A2(n_1308),
.B(n_1309),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1270),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1249),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1320),
.B(n_1343),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1262),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1316),
.A2(n_1296),
.B(n_1293),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1312),
.B(n_1286),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1249),
.Y(n_1355)
);

AOI22x1_ASAP7_75t_SL g1356 ( 
.A1(n_1260),
.A2(n_1280),
.B1(n_1297),
.B2(n_1310),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1357)
);

NOR2x1_ASAP7_75t_R g1358 ( 
.A(n_1253),
.B(n_1338),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1283),
.B(n_1303),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1327),
.A2(n_1305),
.B(n_1314),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1316),
.A2(n_1296),
.B(n_1293),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1261),
.A2(n_1302),
.B(n_1298),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1286),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1269),
.A2(n_1246),
.B(n_1307),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1313),
.B(n_1315),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1333),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1299),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1338),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1306),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1306),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1273),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1318),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1271),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1314),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1273),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1289),
.A2(n_1288),
.B(n_1261),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1323),
.B(n_1346),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1245),
.B(n_1279),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1311),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1317),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1311),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1235),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1245),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1236),
.B(n_1256),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1237),
.A2(n_1340),
.B1(n_1337),
.B2(n_1319),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1237),
.A2(n_1337),
.B1(n_1319),
.B2(n_1334),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1279),
.B(n_1263),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1242),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1250),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1236),
.B(n_1256),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1235),
.Y(n_1391)
);

AO31x2_ASAP7_75t_L g1392 ( 
.A1(n_1251),
.A2(n_1259),
.A3(n_1266),
.B(n_1248),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1283),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1263),
.B(n_1278),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1339),
.A2(n_1285),
.B(n_1332),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1289),
.A2(n_1288),
.B(n_1278),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1322),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1334),
.A2(n_1329),
.B1(n_1277),
.B2(n_1238),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1304),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1249),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1238),
.A2(n_1254),
.B1(n_1258),
.B2(n_1257),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1287),
.B(n_1284),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1290),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1328),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1267),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1287),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1284),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1274),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1282),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1276),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1264),
.B(n_1281),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1272),
.B(n_1255),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1331),
.B(n_1295),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1344),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1291),
.A2(n_1300),
.B(n_1294),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1330),
.B(n_1342),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1300),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1275),
.A2(n_1301),
.B(n_1335),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1352),
.A2(n_1291),
.B(n_1252),
.Y(n_1421)
);

AOI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1385),
.A2(n_1335),
.B1(n_1336),
.B2(n_1326),
.C(n_1345),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1373),
.B(n_1336),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1388),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1386),
.A2(n_1399),
.B1(n_1350),
.B2(n_1411),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1411),
.A2(n_1257),
.B1(n_1258),
.B2(n_1344),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1352),
.A2(n_1292),
.B(n_1341),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1364),
.B(n_1321),
.Y(n_1428)
);

AO32x2_ASAP7_75t_L g1429 ( 
.A1(n_1349),
.A2(n_1324),
.A3(n_1341),
.B1(n_1265),
.B2(n_1247),
.Y(n_1429)
);

AO21x1_ASAP7_75t_L g1430 ( 
.A1(n_1384),
.A2(n_1239),
.B(n_1268),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1384),
.A2(n_1390),
.B(n_1400),
.C(n_1403),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1388),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_SL g1433 ( 
.A1(n_1390),
.A2(n_1400),
.B(n_1401),
.C(n_1404),
.Y(n_1433)
);

BUFx4f_ASAP7_75t_L g1434 ( 
.A(n_1368),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1353),
.A2(n_1357),
.B1(n_1383),
.B2(n_1387),
.C(n_1394),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1378),
.B(n_1369),
.Y(n_1437)
);

NAND2xp33_ASAP7_75t_L g1438 ( 
.A(n_1357),
.B(n_1397),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1369),
.B(n_1370),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1370),
.B(n_1371),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1377),
.B(n_1379),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1388),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_SL g1443 ( 
.A(n_1365),
.B(n_1395),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1366),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1376),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1387),
.A2(n_1397),
.B(n_1394),
.C(n_1360),
.Y(n_1446)
);

AO32x2_ASAP7_75t_L g1447 ( 
.A1(n_1349),
.A2(n_1402),
.A3(n_1373),
.B1(n_1348),
.B2(n_1371),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1408),
.A2(n_1375),
.B1(n_1409),
.B2(n_1393),
.C(n_1405),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1408),
.A2(n_1401),
.B1(n_1404),
.B2(n_1381),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1381),
.B(n_1413),
.Y(n_1450)
);

AOI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1420),
.A2(n_1405),
.B(n_1381),
.C(n_1410),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1363),
.Y(n_1452)
);

AO32x2_ASAP7_75t_L g1453 ( 
.A1(n_1349),
.A2(n_1402),
.A3(n_1348),
.B1(n_1375),
.B2(n_1362),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1410),
.A2(n_1412),
.B1(n_1420),
.B2(n_1418),
.Y(n_1454)
);

BUFx8_ASAP7_75t_SL g1455 ( 
.A(n_1368),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1374),
.B(n_1365),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1376),
.A2(n_1393),
.B(n_1359),
.C(n_1361),
.Y(n_1457)
);

AO32x2_ASAP7_75t_L g1458 ( 
.A1(n_1349),
.A2(n_1402),
.A3(n_1362),
.B1(n_1367),
.B2(n_1354),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1395),
.A2(n_1361),
.B(n_1376),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1359),
.A2(n_1417),
.B(n_1407),
.C(n_1355),
.Y(n_1460)
);

NAND2xp33_ASAP7_75t_L g1461 ( 
.A(n_1414),
.B(n_1412),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1351),
.B(n_1392),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1462),
.B(n_1362),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1457),
.B(n_1362),
.Y(n_1464)
);

NOR3xp33_ASAP7_75t_L g1465 ( 
.A(n_1431),
.B(n_1358),
.C(n_1414),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1424),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1425),
.A2(n_1368),
.B1(n_1407),
.B2(n_1402),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1432),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1436),
.B(n_1362),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1436),
.B(n_1396),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1457),
.B(n_1347),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1432),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1437),
.B(n_1396),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1437),
.B(n_1396),
.Y(n_1474)
);

AND2x4_ASAP7_75t_SL g1475 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1442),
.B(n_1380),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1442),
.Y(n_1477)
);

AND2x4_ASAP7_75t_SL g1478 ( 
.A(n_1456),
.B(n_1365),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1452),
.Y(n_1479)
);

AND2x4_ASAP7_75t_SL g1480 ( 
.A(n_1456),
.B(n_1365),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1443),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1459),
.B(n_1354),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1438),
.A2(n_1407),
.B1(n_1359),
.B2(n_1416),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1440),
.B(n_1396),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1441),
.B(n_1396),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1422),
.A2(n_1418),
.B1(n_1416),
.B2(n_1406),
.C(n_1398),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1439),
.B(n_1389),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1430),
.B(n_1380),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1438),
.A2(n_1359),
.B1(n_1416),
.B2(n_1382),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1435),
.A2(n_1391),
.B1(n_1406),
.B2(n_1372),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1450),
.A2(n_1391),
.B1(n_1372),
.B2(n_1419),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1476),
.B(n_1460),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1464),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1466),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1466),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1475),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1481),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1465),
.A2(n_1448),
.B1(n_1449),
.B2(n_1434),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1468),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1486),
.B(n_1423),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1463),
.B(n_1445),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1475),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1465),
.A2(n_1434),
.B1(n_1455),
.B2(n_1444),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1485),
.B(n_1458),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1472),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1479),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_1454),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1475),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1490),
.A2(n_1446),
.B1(n_1433),
.B2(n_1451),
.C(n_1461),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1485),
.B(n_1458),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1478),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1477),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1463),
.B(n_1445),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1470),
.B(n_1458),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1464),
.B(n_1427),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1470),
.B(n_1453),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1492),
.B(n_1481),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1494),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1492),
.B(n_1421),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1506),
.B(n_1473),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1499),
.B(n_1474),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1495),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1515),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1506),
.B(n_1474),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1509),
.B(n_1484),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1495),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1500),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1515),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1492),
.B(n_1476),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1520),
.B(n_1471),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1501),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1517),
.B(n_1471),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1503),
.B(n_1482),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1500),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1502),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1508),
.Y(n_1542)
);

AND2x4_ASAP7_75t_SL g1543 ( 
.A(n_1496),
.B(n_1504),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1507),
.B(n_1447),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1508),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1492),
.B(n_1496),
.Y(n_1546)
);

NOR2x1_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1488),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1528),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1521),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1521),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1543),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1523),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1523),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1527),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1527),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1536),
.A2(n_1510),
.B(n_1512),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1546),
.B(n_1492),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1546),
.B(n_1497),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1531),
.Y(n_1565)
);

OAI221xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1538),
.A2(n_1512),
.B1(n_1498),
.B2(n_1505),
.C(n_1510),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1543),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1532),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1525),
.B(n_1493),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1543),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1532),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1529),
.B(n_1493),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1503),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1528),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1503),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1539),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

OAI211xp5_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1498),
.B(n_1505),
.C(n_1493),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1540),
.Y(n_1582)
);

OR2x2_ASAP7_75t_SL g1583 ( 
.A(n_1547),
.B(n_1493),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1548),
.B(n_1493),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1548),
.B(n_1493),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1541),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1541),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1542),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1533),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1533),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1559),
.B(n_1562),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1552),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1571),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1576),
.B(n_1530),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1554),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1568),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1587),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1568),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1581),
.B(n_1554),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_1535),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1568),
.Y(n_1604)
);

AOI211xp5_ASAP7_75t_L g1605 ( 
.A1(n_1566),
.A2(n_1433),
.B(n_1519),
.C(n_1522),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1576),
.B(n_1583),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1534),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1583),
.B(n_1530),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1550),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1584),
.B(n_1516),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1550),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1586),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1551),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1555),
.B(n_1535),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1563),
.B(n_1564),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1585),
.B(n_1516),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1564),
.B(n_1467),
.C(n_1573),
.D(n_1426),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1551),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1563),
.B(n_1522),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1570),
.B(n_1535),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1575),
.B(n_1537),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1553),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1578),
.B(n_1516),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1563),
.B(n_1522),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1553),
.B(n_1461),
.C(n_1483),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1592),
.B(n_1573),
.Y(n_1626)
);

OAI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1591),
.A2(n_1524),
.B1(n_1434),
.B2(n_1497),
.C(n_1519),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1563),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1605),
.B(n_1522),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1617),
.B(n_1455),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1613),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1602),
.A2(n_1358),
.B(n_1522),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1613),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1625),
.A2(n_1524),
.B(n_1556),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1607),
.A2(n_1514),
.B1(n_1518),
.B2(n_1524),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1596),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1618),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1537),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1601),
.B(n_1537),
.Y(n_1639)
);

NAND2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1606),
.B(n_1608),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_1356),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1612),
.Y(n_1642)
);

INVxp33_ASAP7_75t_L g1643 ( 
.A(n_1606),
.Y(n_1643)
);

O2A1O1Ixp5_ASAP7_75t_L g1644 ( 
.A1(n_1597),
.A2(n_1608),
.B(n_1596),
.C(n_1612),
.Y(n_1644)
);

NAND2xp33_ASAP7_75t_SL g1645 ( 
.A(n_1597),
.B(n_1544),
.Y(n_1645)
);

AOI33xp33_ASAP7_75t_L g1646 ( 
.A1(n_1600),
.A2(n_1558),
.A3(n_1557),
.B1(n_1588),
.B2(n_1556),
.B3(n_1567),
.Y(n_1646)
);

AOI31xp33_ASAP7_75t_L g1647 ( 
.A1(n_1600),
.A2(n_1524),
.A3(n_1519),
.B(n_1489),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1615),
.A2(n_1511),
.B1(n_1496),
.B2(n_1504),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1618),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1609),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1636),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1631),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1644),
.A2(n_1622),
.B(n_1611),
.C(n_1597),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1640),
.A2(n_1595),
.B1(n_1598),
.B2(n_1599),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1632),
.B(n_1630),
.C(n_1626),
.D(n_1628),
.Y(n_1655)
);

OAI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1643),
.A2(n_1607),
.B(n_1603),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1643),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1633),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1649),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1640),
.A2(n_1599),
.B1(n_1595),
.B2(n_1598),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1634),
.A2(n_1614),
.B1(n_1621),
.B2(n_1620),
.C(n_1594),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1619),
.Y(n_1663)
);

AO22x1_ASAP7_75t_L g1664 ( 
.A1(n_1641),
.A2(n_1624),
.B1(n_1619),
.B2(n_1572),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1638),
.Y(n_1665)
);

XOR2x2_ASAP7_75t_L g1666 ( 
.A(n_1629),
.B(n_1624),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1650),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1650),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1646),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1657),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1663),
.B(n_1639),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1642),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1651),
.B(n_1647),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1665),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1669),
.A2(n_1645),
.B1(n_1627),
.B2(n_1648),
.Y(n_1675)
);

OAI21xp33_ASAP7_75t_L g1676 ( 
.A1(n_1656),
.A2(n_1635),
.B(n_1594),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1666),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1667),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1645),
.B(n_1558),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1653),
.A2(n_1565),
.B(n_1557),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1672),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_1673),
.C(n_1679),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1672),
.B(n_1654),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1677),
.B(n_1655),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1671),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1675),
.B(n_1661),
.C(n_1664),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1674),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_SL g1688 ( 
.A(n_1675),
.B(n_1662),
.C(n_1660),
.D(n_1659),
.Y(n_1688)
);

OAI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1680),
.A2(n_1668),
.B(n_1658),
.C(n_1652),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_L g1690 ( 
.A(n_1676),
.B(n_1662),
.C(n_1616),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1565),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1681),
.B(n_1526),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1683),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1684),
.Y(n_1694)
);

AOI222xp33_ASAP7_75t_L g1695 ( 
.A1(n_1682),
.A2(n_1588),
.B1(n_1574),
.B2(n_1572),
.C1(n_1569),
.C2(n_1567),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_R g1696 ( 
.A(n_1688),
.B(n_1419),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1686),
.A2(n_1623),
.B(n_1616),
.Y(n_1697)
);

AOI222xp33_ASAP7_75t_L g1698 ( 
.A1(n_1693),
.A2(n_1689),
.B1(n_1687),
.B2(n_1685),
.C1(n_1691),
.C2(n_1690),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1696),
.Y(n_1699)
);

AOI211xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1694),
.A2(n_1623),
.B(n_1610),
.C(n_1580),
.Y(n_1700)
);

AOI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1697),
.A2(n_1610),
.B(n_1574),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1692),
.A2(n_1578),
.B1(n_1569),
.B2(n_1582),
.C(n_1580),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1695),
.A2(n_1582),
.B1(n_1579),
.B2(n_1356),
.Y(n_1703)
);

NOR2x1p5_ASAP7_75t_L g1704 ( 
.A(n_1698),
.B(n_1579),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1699),
.B(n_1561),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1700),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1703),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1701),
.Y(n_1708)
);

NAND4xp25_ASAP7_75t_L g1709 ( 
.A(n_1707),
.B(n_1702),
.C(n_1511),
.D(n_1504),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1706),
.B(n_1561),
.Y(n_1710)
);

AOI31xp33_ASAP7_75t_L g1711 ( 
.A1(n_1708),
.A2(n_1705),
.A3(n_1704),
.B(n_1706),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1710),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1712),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1713),
.A2(n_1708),
.B1(n_1712),
.B2(n_1711),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1713),
.B(n_1705),
.Y(n_1715)
);

NOR2xp67_ASAP7_75t_L g1716 ( 
.A(n_1715),
.B(n_1709),
.Y(n_1716)
);

OAI22x1_ASAP7_75t_L g1717 ( 
.A1(n_1714),
.A2(n_1577),
.B1(n_1589),
.B2(n_1590),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1716),
.B(n_1577),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1717),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1719),
.B(n_1549),
.Y(n_1720)
);

AOI22x1_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1718),
.B1(n_1590),
.B2(n_1589),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1589),
.B1(n_1549),
.B2(n_1590),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_R g1723 ( 
.A1(n_1722),
.A2(n_1549),
.B1(n_1429),
.B2(n_1491),
.C(n_1533),
.Y(n_1723)
);

AOI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1415),
.B(n_1542),
.C(n_1545),
.Y(n_1724)
);


endmodule