module real_jpeg_18612_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_419),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_1),
.B(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_34),
.B1(n_52),
.B2(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_55),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g230 ( 
.A1(n_2),
.A2(n_55),
.B1(n_231),
.B2(n_234),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_2),
.A2(n_55),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_3),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_5),
.A2(n_119),
.B1(n_244),
.B2(n_355),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_82),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_82),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_7),
.Y(n_420)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_8),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_8),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_10),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_23)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_11),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_11),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_11),
.A2(n_101),
.A3(n_215),
.B1(n_217),
.B2(n_220),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_153),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_11),
.B(n_127),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_11),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_11),
.B(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_205),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_203),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_186),
.Y(n_17)
);

NOR2xp67_ASAP7_75t_L g204 ( 
.A(n_18),
.B(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.C(n_147),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_19),
.A2(n_128),
.B1(n_129),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_19),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_56),
.B2(n_57),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_20),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_21),
.B(n_236),
.C(n_324),
.Y(n_401)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_22),
.Y(n_188)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_22),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_22),
.A2(n_326),
.B1(n_377),
.B2(n_378),
.Y(n_384)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_42),
.B2(n_51),
.Y(n_22)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_23),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_23),
.A2(n_32),
.B1(n_42),
.B2(n_51),
.Y(n_202)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_27),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_27),
.B(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_28),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_28),
.B(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_32),
.B(n_42),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_38),
.B(n_42),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_33),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_34),
.Y(n_343)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_42),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_42)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_44),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_44),
.Y(n_340)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_87),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_58),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_58),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_78),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_60),
.A2(n_133),
.B(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_60),
.A2(n_68),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2x1p5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_61),
.A2(n_78),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g229 ( 
.A1(n_61),
.A2(n_69),
.B1(n_152),
.B2(n_230),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_61),
.A2(n_69),
.B1(n_152),
.B2(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_61),
.B(n_293),
.Y(n_292)
);

AO22x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_65),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_65),
.Y(n_245)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_65),
.Y(n_247)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_73),
.Y(n_258)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_86),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_87),
.B(n_188),
.C(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_98),
.B1(n_117),
.B2(n_127),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_99),
.B1(n_111),
.B2(n_140),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_89),
.A2(n_99),
.B1(n_111),
.B2(n_140),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_89),
.A2(n_99),
.B(n_111),
.Y(n_378)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_98),
.A2(n_117),
.B1(n_127),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2x1p5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_111)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_114),
.Y(n_233)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_118),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_123),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_129),
.A2(n_130),
.B(n_139),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_139),
.A2(n_309),
.B1(n_310),
.B2(n_314),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_139),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_139),
.B(n_289),
.C(n_312),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_139),
.B(n_202),
.C(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_139),
.A2(n_201),
.B1(n_202),
.B2(n_314),
.Y(n_395)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_146),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_147),
.B(n_416),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_161),
.B(n_182),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_149),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_160),
.Y(n_149)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_150),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_152),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_157),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_157),
.A2(n_255),
.A3(n_259),
.B1(n_261),
.B2(n_266),
.Y(n_254)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_160),
.A2(n_161),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_161),
.A2(n_162),
.B1(n_182),
.B2(n_183),
.Y(n_363)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_163),
.A2(n_242),
.B1(n_354),
.B2(n_357),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_170),
.B(n_223),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_174),
.Y(n_260)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_176),
.Y(n_271)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_178),
.A2(n_243),
.B(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_188),
.Y(n_376)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_201),
.B2(n_202),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_201),
.A2(n_202),
.B1(n_228),
.B2(n_236),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_202),
.B(n_228),
.C(n_352),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_413),
.B(n_418),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AO221x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_347),
.B1(n_349),
.B2(n_406),
.C(n_412),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_318),
.B(n_346),
.Y(n_208)
);

AOI21x1_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_302),
.B(n_317),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_251),
.B(n_301),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_238),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_212),
.B(n_238),
.Y(n_301)
);

XOR2x2_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_213),
.B(n_229),
.C(n_236),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_214),
.B(n_221),
.Y(n_305)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_242),
.B1(n_243),
.B2(n_248),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_228),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_228),
.A2(n_236),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_229),
.A2(n_237),
.B1(n_254),
.B2(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_229),
.B(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_229),
.A2(n_237),
.B1(n_372),
.B2(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_250),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_239),
.A2(n_240),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_305),
.C(n_307),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_239),
.A2(n_240),
.B1(n_353),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_240),
.B(n_353),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_292),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_241),
.A2(n_273),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_276),
.B(n_300),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_272),
.Y(n_252)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_253),
.B(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_273),
.B(n_331),
.Y(n_389)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_295),
.B(n_299),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_291),
.B(n_294),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_289),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_296),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_290),
.A2(n_354),
.B(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_297),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_316),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_307),
.B1(n_308),
.B2(n_315),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_320),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_327),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_328),
.C(n_329),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_341),
.B1(n_344),
.B2(n_345),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_390),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_379),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_364),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_364),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_360),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_351),
.B(n_361),
.C(n_362),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_366),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.C(n_370),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_367),
.Y(n_381)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.C(n_377),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_382),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.C(n_388),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_386),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_389),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_402),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_393),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_398),
.C(n_400),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_400),
.B2(n_401),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_409),
.Y(n_408)
);

NAND2x1_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_405),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B(n_410),
.C(n_411),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_415),
.Y(n_418)
);


endmodule