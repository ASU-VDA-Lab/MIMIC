module fake_jpeg_11274_n_584 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_584);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_21),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_76),
.Y(n_136)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_72),
.Y(n_153)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_86),
.Y(n_127)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_16),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_82),
.Y(n_192)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_13),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_14),
.B1(n_13),
.B2(n_10),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_48),
.B1(n_120),
.B2(n_84),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_39),
.B(n_14),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_108),
.B(n_115),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_112),
.B(n_119),
.Y(n_185)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_52),
.Y(n_159)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_118),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_48),
.B(n_14),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_120),
.B(n_8),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_133),
.A2(n_140),
.B1(n_166),
.B2(n_45),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_27),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_41),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_68),
.B(n_55),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_157),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_70),
.B(n_55),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_159),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_89),
.A2(n_17),
.B1(n_50),
.B2(n_46),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_97),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_174),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_74),
.A2(n_26),
.B1(n_42),
.B2(n_53),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_172),
.A2(n_179),
.B1(n_37),
.B2(n_1),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_62),
.B(n_33),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_53),
.C(n_36),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_191),
.C(n_118),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_85),
.A2(n_29),
.B1(n_36),
.B2(n_46),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_63),
.A2(n_33),
.B1(n_35),
.B2(n_43),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_181),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_92),
.A2(n_29),
.B(n_50),
.C(n_43),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_184),
.A2(n_37),
.B1(n_45),
.B2(n_52),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_131),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_59),
.B(n_35),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_189),
.B(n_193),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_88),
.A2(n_45),
.B1(n_52),
.B2(n_14),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_87),
.B(n_10),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_87),
.B(n_9),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_9),
.Y(n_199)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_197),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_198),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_199),
.B(n_211),
.Y(n_273)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_201),
.Y(n_287)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_202),
.Y(n_298)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_203),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_64),
.B1(n_79),
.B2(n_80),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_204),
.A2(n_225),
.B1(n_137),
.B2(n_155),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_159),
.A2(n_82),
.B1(n_90),
.B2(n_81),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_205),
.A2(n_222),
.B1(n_263),
.B2(n_170),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_208),
.Y(n_310)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_209),
.Y(n_302)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_224),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_114),
.C(n_107),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_212),
.B(n_205),
.C(n_240),
.Y(n_301)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_213),
.Y(n_313)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_214),
.Y(n_318)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_179),
.A2(n_102),
.B1(n_96),
.B2(n_94),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_142),
.A2(n_103),
.B1(n_176),
.B2(n_151),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_229),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_227),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_228),
.A2(n_236),
.B1(n_240),
.B2(n_242),
.Y(n_279)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_129),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_231),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_162),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_234),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_156),
.A2(n_8),
.B1(n_45),
.B2(n_52),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

INVx13_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_169),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_243),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_156),
.A2(n_52),
.B1(n_45),
.B2(n_37),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_244),
.Y(n_291)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_143),
.Y(n_243)
);

INVx5_ASAP7_75t_SL g244 ( 
.A(n_153),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_246),
.Y(n_283)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_144),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_131),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_248),
.Y(n_288)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_139),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_250),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_183),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_136),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_251),
.A2(n_195),
.B1(n_137),
.B2(n_122),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_125),
.B(n_0),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_252),
.B(n_257),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_280)
);

INVx5_ASAP7_75t_SL g254 ( 
.A(n_184),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_146),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_178),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_123),
.B(n_2),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_260),
.B(n_3),
.Y(n_285)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_130),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_130),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_161),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_265),
.A2(n_244),
.B1(n_217),
.B2(n_243),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_215),
.B(n_172),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_270),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_122),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_272),
.A2(n_281),
.B1(n_284),
.B2(n_294),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_207),
.B(n_138),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_289),
.Y(n_343)
);

NOR4xp25_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_165),
.C(n_155),
.D(n_194),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_285),
.C(n_4),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_2),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_282),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_204),
.A2(n_194),
.B1(n_149),
.B2(n_147),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_206),
.B(n_211),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_290),
.A2(n_306),
.B1(n_309),
.B2(n_314),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_234),
.A2(n_149),
.B1(n_147),
.B2(n_192),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_227),
.C(n_236),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_206),
.B(n_152),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_319),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_222),
.A2(n_192),
.B1(n_152),
.B2(n_158),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_229),
.A2(n_170),
.B1(n_158),
.B2(n_190),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_311),
.A2(n_267),
.B1(n_203),
.B2(n_200),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_225),
.A2(n_190),
.B1(n_173),
.B2(n_5),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_5),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_4),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_223),
.B(n_4),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_7),
.Y(n_357)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_275),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_324),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_303),
.B(n_265),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_323),
.B(n_332),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_289),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_358),
.C(n_307),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_270),
.B(n_256),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_339),
.Y(n_384)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_268),
.Y(n_328)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_227),
.C(n_248),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_329),
.B(n_337),
.C(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_336),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_273),
.B(n_237),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_269),
.A2(n_238),
.B(n_245),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_345),
.B(n_283),
.Y(n_370)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_266),
.B(n_201),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_219),
.C(n_228),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_297),
.B(n_214),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_346),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_312),
.B1(n_284),
.B2(n_282),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_360),
.B1(n_362),
.B2(n_316),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_293),
.A2(n_242),
.B(n_246),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_297),
.B(n_253),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_355),
.Y(n_388)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_349),
.Y(n_386)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_282),
.A2(n_5),
.B(n_6),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_351),
.A2(n_359),
.B(n_287),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_352),
.B(n_357),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_353),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_6),
.C(n_7),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_276),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_291),
.B(n_7),
.C(n_305),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_280),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_282),
.B1(n_294),
.B2(n_281),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_285),
.B(n_320),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_298),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_272),
.A2(n_290),
.B1(n_291),
.B2(n_306),
.Y(n_362)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_291),
.A3(n_278),
.B1(n_273),
.B2(n_319),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_389),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_325),
.A2(n_286),
.B1(n_279),
.B2(n_296),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_366),
.A2(n_370),
.B(n_372),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_340),
.A2(n_309),
.B1(n_315),
.B2(n_314),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_367),
.A2(n_377),
.B1(n_380),
.B2(n_382),
.Y(n_414)
);

AOI32xp33_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_267),
.A3(n_304),
.B1(n_308),
.B2(n_295),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_296),
.B1(n_300),
.B2(n_271),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_383),
.B1(n_387),
.B2(n_396),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_359),
.A2(n_304),
.B(n_308),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_375),
.A2(n_330),
.B(n_354),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_360),
.A2(n_318),
.B1(n_300),
.B2(n_310),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_378),
.A2(n_393),
.B(n_351),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_356),
.A2(n_313),
.B1(n_292),
.B2(n_302),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_327),
.A2(n_310),
.B1(n_316),
.B2(n_313),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_358),
.A2(n_302),
.B1(n_298),
.B2(n_287),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_266),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_390),
.B(n_361),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_355),
.C(n_326),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_307),
.B(n_317),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_356),
.A2(n_307),
.B1(n_317),
.B2(n_334),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_397),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_317),
.B1(n_330),
.B2(n_329),
.Y(n_396)
);

OAI22x1_ASAP7_75t_SL g397 ( 
.A1(n_345),
.A2(n_321),
.B1(n_339),
.B2(n_347),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_386),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_400),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_379),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_405),
.C(n_420),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_363),
.B(n_390),
.Y(n_403)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_350),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_408),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_350),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_409),
.B(n_416),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_410),
.A2(n_370),
.B(n_373),
.Y(n_457)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_396),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_388),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_364),
.B(n_332),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_422),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_418),
.A2(n_426),
.B(n_375),
.Y(n_435)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_328),
.C(n_338),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_378),
.A2(n_348),
.B(n_341),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_383),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_342),
.Y(n_424)
);

NAND2x1_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_372),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_374),
.A2(n_357),
.B1(n_346),
.B2(n_335),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_380),
.B1(n_377),
.B2(n_382),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_352),
.B(n_349),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_398),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_430),
.Y(n_462)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_363),
.B(n_353),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_431),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_395),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_440),
.C(n_441),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_435),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_438),
.B(n_458),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_420),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_391),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_414),
.B1(n_429),
.B2(n_408),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_388),
.C(n_389),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_445),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_400),
.A2(n_404),
.B1(n_414),
.B2(n_416),
.Y(n_448)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_431),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_413),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_451),
.A2(n_457),
.B(n_407),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_397),
.B1(n_367),
.B2(n_384),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_453),
.A2(n_456),
.B1(n_429),
.B2(n_422),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_406),
.A2(n_384),
.B1(n_376),
.B2(n_366),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_403),
.B(n_365),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_456),
.Y(n_505)
);

NOR3xp33_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_373),
.C(n_447),
.Y(n_465)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_487),
.C(n_460),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_399),
.Y(n_467)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_467),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_462),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_468),
.B(n_473),
.Y(n_503)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_462),
.Y(n_469)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_474),
.B1(n_415),
.B2(n_371),
.Y(n_512)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_472),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_449),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_439),
.B(n_409),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_475),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_449),
.A2(n_424),
.B1(n_401),
.B2(n_421),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_476),
.A2(n_482),
.B1(n_485),
.B2(n_453),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_430),
.Y(n_478)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_424),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_479),
.Y(n_491)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_434),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_481),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_436),
.A2(n_401),
.B(n_407),
.C(n_424),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_436),
.A2(n_410),
.B1(n_425),
.B2(n_428),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_483),
.A2(n_484),
.B1(n_488),
.B2(n_460),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_432),
.A2(n_427),
.B1(n_411),
.B2(n_423),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_437),
.B(n_419),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_451),
.A2(n_418),
.B(n_426),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_489),
.A2(n_435),
.B(n_451),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_492),
.A2(n_511),
.B(n_477),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_493),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_486),
.B(n_438),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_496),
.B(n_505),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_466),
.B(n_443),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_498),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_472),
.B(n_443),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_433),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_387),
.Y(n_529)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_507),
.Y(n_520)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_463),
.A2(n_442),
.B1(n_444),
.B2(n_458),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_474),
.B1(n_470),
.B2(n_489),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_487),
.B(n_441),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_510),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_463),
.A2(n_459),
.B1(n_452),
.B2(n_446),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_477),
.A2(n_459),
.B(n_452),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_482),
.B1(n_476),
.B2(n_468),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_513),
.A2(n_505),
.B1(n_501),
.B2(n_494),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_502),
.A2(n_467),
.B1(n_473),
.B2(n_469),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_519),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_529),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_495),
.B(n_478),
.Y(n_518)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_518),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_471),
.C(n_440),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_521),
.A2(n_525),
.B1(n_526),
.B2(n_490),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_486),
.C(n_464),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_523),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_479),
.C(n_483),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_493),
.A2(n_479),
.B1(n_481),
.B2(n_480),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_490),
.A2(n_488),
.B1(n_485),
.B2(n_371),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_504),
.B(n_385),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_504),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_517),
.A2(n_522),
.B1(n_528),
.B2(n_513),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_532),
.A2(n_545),
.B1(n_526),
.B2(n_524),
.Y(n_557)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_518),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_535),
.B(n_538),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_542),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_512),
.C(n_491),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_521),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_514),
.B(n_495),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_540),
.B(n_541),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_491),
.C(n_511),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_503),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_520),
.B(n_507),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_543),
.B(n_494),
.Y(n_555)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_530),
.B(n_503),
.CI(n_492),
.CON(n_545),
.SN(n_545)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_531),
.A2(n_517),
.B1(n_528),
.B2(n_501),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_548),
.B(n_551),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_536),
.A2(n_516),
.B(n_527),
.Y(n_549)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_549),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_554),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_525),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_542),
.C(n_532),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_552),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_524),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_555),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_533),
.Y(n_563)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_563),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_556),
.A2(n_537),
.B1(n_545),
.B2(n_539),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_564),
.B(n_565),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g565 ( 
.A1(n_553),
.A2(n_545),
.B(n_533),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_546),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_552),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_567),
.A2(n_571),
.B(n_558),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_547),
.C(n_551),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_570),
.B(n_572),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_547),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_561),
.B(n_550),
.Y(n_572)
);

OAI21xp33_ASAP7_75t_L g573 ( 
.A1(n_568),
.A2(n_562),
.B(n_560),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_573),
.A2(n_574),
.B(n_576),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_559),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_575),
.B(n_569),
.C(n_563),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_578),
.A2(n_554),
.B(n_564),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_579),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_580),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_577),
.B(n_369),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_369),
.C(n_353),
.Y(n_583)
);

O2A1O1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_583),
.A2(n_369),
.B(n_392),
.C(n_577),
.Y(n_584)
);


endmodule