module real_aes_684_n_12 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10, n_11, n_12);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
input n_10;
input n_11;
output n_12;
wire n_28;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_19;
wire n_25;
wire n_30;
wire n_14;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_0), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_1), .B(n_5), .C(n_21), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_2), .Y(n_21) );
AOI22xp33_ASAP7_75t_SL g12 ( .A1(n_3), .A2(n_9), .B1(n_13), .B2(n_28), .Y(n_12) );
NAND3xp33_ASAP7_75t_SL g24 ( .A(n_4), .B(n_25), .C(n_26), .Y(n_24) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_6), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_7), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_8), .B(n_16), .Y(n_15) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_8), .B(n_30), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_10), .Y(n_23) );
NAND2xp33_ASAP7_75t_SL g31 ( .A(n_10), .B(n_18), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_11), .B(n_27), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
OR2x2_ASAP7_75t_L g16 ( .A(n_17), .B(n_24), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_18), .B(n_23), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g19 ( .A(n_20), .B(n_22), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_24), .B(n_31), .Y(n_30) );
CKINVDCx14_ASAP7_75t_R g28 ( .A(n_29), .Y(n_28) );
endmodule