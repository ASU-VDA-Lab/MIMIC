module real_jpeg_33463_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_12;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22x1_ASAP7_75t_SL g21 ( 
.A1(n_0),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

OAI22x1_ASAP7_75t_SL g93 ( 
.A1(n_0),
.A2(n_25),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

AOI22x1_ASAP7_75t_L g176 ( 
.A1(n_0),
.A2(n_25),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_0),
.A2(n_203),
.A3(n_209),
.B1(n_213),
.B2(n_221),
.Y(n_202)
);

NAND2xp67_ASAP7_75t_SL g276 ( 
.A(n_0),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_0),
.B(n_240),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_1),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_4),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_4),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_5),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_5),
.Y(n_317)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_6),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22x1_ASAP7_75t_L g79 ( 
.A1(n_8),
.A2(n_60),
.B1(n_80),
.B2(n_84),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_8),
.A2(n_60),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_8),
.A2(n_60),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_9),
.Y(n_163)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_9),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_297),
.Y(n_11)
);

INVxp67_ASAP7_75t_SL g12 ( 
.A(n_13),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_231),
.B(n_294),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_186),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_15),
.B(n_186),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_132),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_99),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_17),
.B(n_132),
.C(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_64),
.C(n_71),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_18),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_18),
.B(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_19),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B1(n_44),
.B2(n_55),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22x1_ASAP7_75t_L g183 ( 
.A1(n_21),
.A2(n_31),
.B1(n_45),
.B2(n_56),
.Y(n_183)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_25),
.B(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_25),
.A2(n_121),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_25),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_25),
.B(n_32),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_25),
.B(n_262),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_SL g267 ( 
.A1(n_25),
.A2(n_167),
.B(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_46),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_33),
.B(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_33),
.Y(n_264)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_35),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_35),
.Y(n_199)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_38),
.Y(n_217)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_49),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_64),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_190)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_71),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_71),
.B(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_72),
.B(n_275),
.Y(n_274)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B(n_88),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_77),
.Y(n_277)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_79),
.A2(n_89),
.B1(n_93),
.B2(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_83),
.Y(n_272)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_87),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_88),
.A2(n_314),
.B(n_321),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

NOR2x1_ASAP7_75t_R g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_90),
.Y(n_230)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_93),
.B(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_95),
.Y(n_316)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_99),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_126),
.B1(n_127),
.B2(n_131),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_101),
.B(n_126),
.Y(n_304)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.A3(n_109),
.B1(n_114),
.B2(n_121),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_106),
.A3(n_109),
.B1(n_114),
.B2(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_126),
.B(n_192),
.C(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_126),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_R g280 ( 
.A(n_127),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_127),
.B(n_281),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_156),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_135),
.B(n_157),
.C(n_185),
.Y(n_311)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_144),
.B(n_145),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_137),
.A2(n_144),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_146),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_149),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_175),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.Y(n_158)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_167),
.B(n_170),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_166),
.B1(n_176),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_160),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_R g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

AOI22x1_ASAP7_75t_L g238 ( 
.A1(n_175),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_182),
.A2(n_185),
.B1(n_237),
.B2(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.C(n_200),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_200),
.B1(n_201),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_192),
.A2(n_193),
.B1(n_253),
.B2(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_227),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_227),
.Y(n_242)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_243),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_243),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.C(n_242),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_251),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_260),
.Y(n_285)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_237),
.B(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_292),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_254),
.B(n_290),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_284),
.B(n_289),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_273),
.B(n_283),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_265),
.B(n_267),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_280),
.B(n_282),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_324),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_302),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx4f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);


endmodule