module real_aes_8575_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_730, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_730;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_725;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g464 ( .A1(n_0), .A2(n_202), .B(n_465), .C(n_468), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_1), .B(n_459), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_1), .A2(n_715), .B1(n_716), .B2(n_724), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_1), .Y(n_724) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g237 ( .A(n_3), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_4), .B(n_154), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_5), .A2(n_454), .B(n_542), .Y(n_541) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_6), .A2(n_177), .B(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_7), .A2(n_38), .B1(n_147), .B2(n_171), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_8), .B(n_177), .Y(n_249) );
AND2x6_ASAP7_75t_L g162 ( .A(n_9), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_10), .A2(n_162), .B(n_445), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_11), .B(n_39), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_11), .B(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_13), .B(n_152), .Y(n_185) );
INVx1_ASAP7_75t_L g229 ( .A(n_14), .Y(n_229) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_15), .A2(n_76), .B1(n_718), .B2(n_719), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_15), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_16), .B(n_154), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_17), .B(n_178), .Y(n_216) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_18), .A2(n_176), .A3(n_177), .B1(n_200), .B2(n_204), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_19), .B(n_147), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_20), .B(n_178), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_21), .A2(n_56), .B1(n_147), .B2(n_171), .Y(n_203) );
AOI22xp33_ASAP7_75t_SL g174 ( .A1(n_22), .A2(n_82), .B1(n_147), .B2(n_152), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_23), .B(n_147), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_24), .A2(n_176), .B(n_445), .C(n_492), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_25), .A2(n_176), .B(n_445), .C(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_26), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_27), .B(n_139), .Y(n_258) );
OAI22xp5_ASAP7_75t_SL g701 ( .A1(n_28), .A2(n_94), .B1(n_702), .B2(n_703), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_28), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_29), .A2(n_700), .B1(n_701), .B2(n_704), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_29), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_30), .A2(n_454), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_31), .B(n_139), .Y(n_164) );
INVx2_ASAP7_75t_L g149 ( .A(n_32), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_33), .A2(n_451), .B(n_477), .C(n_478), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_34), .B(n_147), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_35), .B(n_139), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_36), .A2(n_43), .B1(n_435), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_36), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_37), .B(n_187), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_40), .B(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_41), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_42), .B(n_154), .Y(n_530) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_43), .A2(n_130), .B1(n_435), .B2(n_436), .Y(n_129) );
INVx1_ASAP7_75t_L g435 ( .A(n_43), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_44), .B(n_454), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_45), .B(n_118), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_46), .A2(n_451), .B(n_477), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_47), .B(n_147), .Y(n_244) );
INVx1_ASAP7_75t_L g466 ( .A(n_48), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_49), .A2(n_92), .B1(n_171), .B2(n_172), .Y(n_170) );
INVx1_ASAP7_75t_L g529 ( .A(n_50), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_51), .B(n_147), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_52), .B(n_147), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_53), .A2(n_698), .B1(n_699), .B2(n_705), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_53), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_54), .B(n_454), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_55), .B(n_235), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g220 ( .A1(n_57), .A2(n_61), .B1(n_147), .B2(n_152), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_58), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_59), .B(n_147), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_60), .B(n_147), .Y(n_257) );
INVx1_ASAP7_75t_L g163 ( .A(n_62), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_63), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_64), .B(n_459), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_65), .A2(n_232), .B(n_235), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_66), .B(n_147), .Y(n_238) );
INVx1_ASAP7_75t_L g142 ( .A(n_67), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_68), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_69), .B(n_154), .Y(n_482) );
AO32x2_ASAP7_75t_L g168 ( .A1(n_70), .A2(n_169), .A3(n_175), .B1(n_176), .B2(n_177), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_71), .B(n_155), .Y(n_519) );
INVx1_ASAP7_75t_L g256 ( .A(n_72), .Y(n_256) );
INVx1_ASAP7_75t_L g150 ( .A(n_73), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_74), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_75), .B(n_481), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_76), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_77), .A2(n_445), .B(n_447), .C(n_451), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_78), .B(n_152), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_79), .Y(n_543) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_81), .B(n_480), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_83), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_84), .B(n_171), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_85), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_86), .B(n_152), .Y(n_159) );
INVx2_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_88), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_89), .B(n_173), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_90), .B(n_152), .Y(n_245) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_91), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g120 ( .A(n_91), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g128 ( .A(n_91), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_93), .A2(n_104), .B1(n_152), .B2(n_153), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_94), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_95), .B(n_454), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_96), .Y(n_479) );
INVxp67_ASAP7_75t_L g546 ( .A(n_97), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_98), .A2(n_106), .B1(n_116), .B2(n_728), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_99), .B(n_152), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_100), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g448 ( .A(n_101), .Y(n_448) );
INVx1_ASAP7_75t_L g515 ( .A(n_102), .Y(n_515) );
AND2x2_ASAP7_75t_L g531 ( .A(n_103), .B(n_139), .Y(n_531) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g728 ( .A(n_108), .Y(n_728) );
CKINVDCx12_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x2_ASAP7_75t_L g122 ( .A(n_112), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
NAND2x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_124), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g727 ( .A(n_120), .Y(n_727) );
NOR2x2_ASAP7_75t_L g710 ( .A(n_121), .B(n_128), .Y(n_710) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g125 ( .A1(n_122), .A2(n_126), .B1(n_127), .B2(n_697), .C(n_706), .Y(n_125) );
OAI321xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_707), .A3(n_711), .B1(n_714), .B2(n_725), .C(n_726), .Y(n_124) );
INVx1_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
AO22x2_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_129), .B1(n_437), .B2(n_696), .Y(n_127) );
INVx1_ASAP7_75t_L g696 ( .A(n_128), .Y(n_696) );
INVx1_ASAP7_75t_L g436 ( .A(n_130), .Y(n_436) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_130), .A2(n_436), .B1(n_721), .B2(n_722), .Y(n_720) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_356), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_305), .C(n_347), .Y(n_131) );
AOI211xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_210), .B(n_259), .C(n_281), .Y(n_132) );
OAI211xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_165), .B(n_193), .C(n_205), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_135), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g368 ( .A(n_135), .B(n_285), .Y(n_368) );
BUFx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g270 ( .A(n_136), .B(n_196), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_136), .B(n_181), .Y(n_387) );
INVx1_ASAP7_75t_L g405 ( .A(n_136), .Y(n_405) );
AND2x2_ASAP7_75t_L g414 ( .A(n_136), .B(n_302), .Y(n_414) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g297 ( .A(n_137), .B(n_181), .Y(n_297) );
AND2x2_ASAP7_75t_L g355 ( .A(n_137), .B(n_302), .Y(n_355) );
INVx1_ASAP7_75t_L g399 ( .A(n_137), .Y(n_399) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g276 ( .A(n_138), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g284 ( .A(n_138), .Y(n_284) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_138), .Y(n_324) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .B(n_164), .Y(n_138) );
INVx2_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_139), .A2(n_182), .B(n_192), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_139), .A2(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g498 ( .A(n_139), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_139), .A2(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_L g178 ( .A(n_140), .B(n_141), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_157), .B(n_162), .Y(n_144) );
O2A1O1Ixp5_ASAP7_75t_SL g145 ( .A1(n_146), .A2(n_150), .B(n_151), .C(n_154), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_147), .Y(n_450) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AND2x6_ASAP7_75t_L g445 ( .A(n_148), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g153 ( .A(n_149), .Y(n_153) );
INVx1_ASAP7_75t_L g236 ( .A(n_149), .Y(n_236) );
INVx2_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_154), .A2(n_244), .B(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_154), .A2(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_154), .B(n_546), .Y(n_545) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_155), .A2(n_170), .B1(n_173), .B2(n_174), .Y(n_169) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
INVx1_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
INVx1_ASAP7_75t_L g446 ( .A(n_156), .Y(n_446) );
AND2x2_ASAP7_75t_L g455 ( .A(n_156), .B(n_236), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_160), .Y(n_157) );
INVx1_ASAP7_75t_L g232 ( .A(n_160), .Y(n_232) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g481 ( .A(n_161), .Y(n_481) );
BUFx3_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_162), .A2(n_183), .B(n_188), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_162), .A2(n_228), .B(n_233), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_162), .A2(n_243), .B(n_246), .Y(n_242) );
INVx4_ASAP7_75t_SL g452 ( .A(n_162), .Y(n_452) );
AND2x4_ASAP7_75t_L g454 ( .A(n_162), .B(n_455), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_162), .B(n_455), .Y(n_516) );
INVxp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
AND2x2_ASAP7_75t_L g263 ( .A(n_167), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g296 ( .A(n_167), .Y(n_296) );
OR2x2_ASAP7_75t_L g422 ( .A(n_167), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_167), .B(n_181), .Y(n_426) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
INVx1_ASAP7_75t_L g208 ( .A(n_168), .Y(n_208) );
AND2x2_ASAP7_75t_L g285 ( .A(n_168), .B(n_198), .Y(n_285) );
AND2x2_ASAP7_75t_L g325 ( .A(n_168), .B(n_199), .Y(n_325) );
INVx2_ASAP7_75t_L g468 ( .A(n_172), .Y(n_468) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_172), .Y(n_483) );
INVx2_ASAP7_75t_L g191 ( .A(n_173), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_173), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_173), .A2(n_202), .B1(n_219), .B2(n_220), .Y(n_218) );
INVx4_ASAP7_75t_L g467 ( .A(n_173), .Y(n_467) );
INVx1_ASAP7_75t_L g495 ( .A(n_175), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g217 ( .A(n_176), .B(n_218), .C(n_221), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_176), .A2(n_252), .B(n_255), .Y(n_251) );
INVx4_ASAP7_75t_L g221 ( .A(n_177), .Y(n_221) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_177), .A2(n_242), .B(n_249), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_177), .A2(n_505), .B(n_506), .Y(n_504) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_177), .Y(n_540) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
INVxp67_ASAP7_75t_L g367 ( .A(n_179), .Y(n_367) );
AND2x4_ASAP7_75t_L g392 ( .A(n_179), .B(n_285), .Y(n_392) );
BUFx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_SL g283 ( .A(n_180), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g197 ( .A(n_181), .B(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g271 ( .A(n_181), .B(n_199), .Y(n_271) );
INVx1_ASAP7_75t_L g277 ( .A(n_181), .Y(n_277) );
INVx2_ASAP7_75t_L g303 ( .A(n_181), .Y(n_303) );
AND2x2_ASAP7_75t_L g319 ( .A(n_181), .B(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
O2A1O1Ixp5_ASAP7_75t_L g255 ( .A1(n_191), .A2(n_234), .B(n_256), .C(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_194), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_197), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g274 ( .A(n_196), .Y(n_274) );
AND2x2_ASAP7_75t_L g382 ( .A(n_196), .B(n_198), .Y(n_382) );
AND2x2_ASAP7_75t_L g299 ( .A(n_197), .B(n_284), .Y(n_299) );
AND2x2_ASAP7_75t_L g398 ( .A(n_197), .B(n_399), .Y(n_398) );
NOR2xp67_ASAP7_75t_L g320 ( .A(n_198), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g423 ( .A(n_198), .B(n_284), .Y(n_423) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx2_ASAP7_75t_L g209 ( .A(n_199), .Y(n_209) );
AND2x2_ASAP7_75t_L g302 ( .A(n_199), .B(n_303), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_202), .A2(n_234), .B(n_237), .C(n_238), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_202), .A2(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g226 ( .A(n_204), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_204), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_209), .Y(n_206) );
AND2x2_ASAP7_75t_L g348 ( .A(n_207), .B(n_283), .Y(n_348) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_208), .B(n_284), .Y(n_333) );
INVx2_ASAP7_75t_L g332 ( .A(n_209), .Y(n_332) );
OAI222xp33_ASAP7_75t_L g336 ( .A1(n_209), .A2(n_276), .B1(n_337), .B2(n_339), .C1(n_340), .C2(n_343), .Y(n_336) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g261 ( .A(n_214), .Y(n_261) );
OR2x2_ASAP7_75t_L g372 ( .A(n_214), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g294 ( .A(n_215), .Y(n_294) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_215), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g351 ( .A(n_215), .B(n_265), .Y(n_351) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
INVx1_ASAP7_75t_L g312 ( .A(n_216), .Y(n_312) );
AO21x1_ASAP7_75t_L g311 ( .A1(n_218), .A2(n_221), .B(n_312), .Y(n_311) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_221), .A2(n_443), .B(n_456), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_221), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g459 ( .A(n_221), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_221), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_221), .A2(n_514), .B(n_521), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_222), .A2(n_315), .B1(n_354), .B2(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_240), .Y(n_222) );
INVx3_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
OR2x2_ASAP7_75t_L g420 ( .A(n_223), .B(n_296), .Y(n_420) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g293 ( .A(n_224), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_224), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g317 ( .A(n_224), .B(n_265), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_224), .B(n_241), .Y(n_373) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g264 ( .A(n_225), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g268 ( .A(n_225), .B(n_241), .Y(n_268) );
AND2x2_ASAP7_75t_L g344 ( .A(n_225), .B(n_291), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_225), .B(n_250), .Y(n_384) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_239), .Y(n_225) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_226), .A2(n_251), .B(n_258), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .C(n_232), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_230), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_230), .A2(n_519), .B(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_232), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_234), .A2(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_240), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g300 ( .A(n_240), .B(n_261), .Y(n_300) );
AND2x2_ASAP7_75t_L g304 ( .A(n_240), .B(n_294), .Y(n_304) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
INVx3_ASAP7_75t_L g265 ( .A(n_241), .Y(n_265) );
AND2x2_ASAP7_75t_L g290 ( .A(n_241), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g425 ( .A(n_241), .B(n_408), .Y(n_425) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_250), .Y(n_279) );
INVx2_ASAP7_75t_L g291 ( .A(n_250), .Y(n_291) );
AND2x2_ASAP7_75t_L g335 ( .A(n_250), .B(n_311), .Y(n_335) );
INVx1_ASAP7_75t_L g378 ( .A(n_250), .Y(n_378) );
OR2x2_ASAP7_75t_L g409 ( .A(n_250), .B(n_311), .Y(n_409) );
AND2x2_ASAP7_75t_L g429 ( .A(n_250), .B(n_265), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B(n_266), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g267 ( .A(n_261), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_261), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g386 ( .A(n_263), .Y(n_386) );
INVx2_ASAP7_75t_SL g280 ( .A(n_264), .Y(n_280) );
AND2x2_ASAP7_75t_L g400 ( .A(n_264), .B(n_294), .Y(n_400) );
INVx2_ASAP7_75t_L g346 ( .A(n_265), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_265), .B(n_378), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_269), .B1(n_272), .B2(n_278), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_268), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g434 ( .A(n_268), .Y(n_434) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g359 ( .A(n_270), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_270), .B(n_302), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_271), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g375 ( .A(n_271), .B(n_324), .Y(n_375) );
INVx2_ASAP7_75t_L g431 ( .A(n_271), .Y(n_431) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g301 ( .A(n_274), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_274), .B(n_319), .Y(n_352) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_276), .B(n_296), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g413 ( .A(n_279), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_SL g363 ( .A1(n_280), .A2(n_364), .B(n_366), .C(n_369), .Y(n_363) );
OR2x2_ASAP7_75t_L g390 ( .A(n_280), .B(n_294), .Y(n_390) );
OAI221xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_286), .B1(n_288), .B2(n_295), .C(n_298), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_283), .B(n_332), .Y(n_339) );
AND2x2_ASAP7_75t_L g381 ( .A(n_283), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g417 ( .A(n_283), .Y(n_417) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
INVx1_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
NOR2xp67_ASAP7_75t_L g341 ( .A(n_287), .B(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g395 ( .A(n_287), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_287), .B(n_335), .Y(n_411) );
INVx2_ASAP7_75t_L g397 ( .A(n_288), .Y(n_397) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g338 ( .A(n_290), .B(n_309), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_290), .A2(n_306), .B(n_348), .C(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g316 ( .A(n_291), .B(n_311), .Y(n_316) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_295), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OR2x2_ASAP7_75t_L g364 ( .A(n_296), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_301), .B2(n_304), .Y(n_298) );
INVx1_ASAP7_75t_L g418 ( .A(n_300), .Y(n_418) );
INVx1_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
INVx1_ASAP7_75t_L g416 ( .A(n_304), .Y(n_416) );
AOI211xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_309), .B(n_313), .C(n_336), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g328 ( .A(n_308), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g379 ( .A(n_309), .Y(n_379) );
AND2x2_ASAP7_75t_L g428 ( .A(n_309), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B(n_326), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_316), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g334 ( .A(n_317), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g410 ( .A(n_317), .Y(n_410) );
OAI32xp33_ASAP7_75t_L g421 ( .A1(n_317), .A2(n_369), .A3(n_376), .B1(n_417), .B2(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_SL g389 ( .A(n_319), .Y(n_389) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g329 ( .A(n_325), .Y(n_329) );
OAI21xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B(n_334), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_328), .A2(n_376), .B1(n_402), .B2(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_332), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g362 ( .A(n_346), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_401), .Y(n_396) );
NAND5xp2_ASAP7_75t_L g356 ( .A(n_357), .B(n_380), .C(n_396), .D(n_406), .E(n_424), .Y(n_356) );
AOI211xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_360), .B(n_363), .C(n_370), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g427 ( .A(n_364), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_374), .B2(n_376), .Y(n_370) );
INVx1_ASAP7_75t_SL g403 ( .A(n_373), .Y(n_403) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_376), .A2(n_386), .A3(n_387), .B1(n_388), .B2(n_389), .C1(n_390), .C2(n_391), .Y(n_385) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g388 ( .A(n_378), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_378), .B(n_403), .Y(n_402) );
AOI211xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_383), .B(n_385), .C(n_393), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_389), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_415) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_414), .B1(n_415), .B2(n_419), .C(n_421), .Y(n_406) );
OAI211xp5_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_410), .B(n_411), .C(n_412), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g433 ( .A(n_409), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_427), .B2(n_428), .C(n_430), .Y(n_424) );
AOI21xp33_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_432), .B(n_433), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_438), .B(n_639), .Y(n_437) );
AND4x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_579), .C(n_594), .D(n_619), .Y(n_438) );
NOR2xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_552), .Y(n_439) );
OAI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_470), .B(n_532), .Y(n_440) );
AND2x2_ASAP7_75t_L g582 ( .A(n_441), .B(n_487), .Y(n_582) );
AND2x2_ASAP7_75t_L g595 ( .A(n_441), .B(n_486), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_441), .B(n_471), .Y(n_645) );
INVx1_ASAP7_75t_L g649 ( .A(n_441), .Y(n_649) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_458), .Y(n_441) );
INVx2_ASAP7_75t_L g566 ( .A(n_442), .Y(n_566) );
BUFx2_ASAP7_75t_L g593 ( .A(n_442), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_453), .Y(n_443) );
INVx5_ASAP7_75t_L g463 ( .A(n_445), .Y(n_463) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_SL g461 ( .A1(n_452), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_452), .A2(n_463), .B(n_543), .C(n_544), .Y(n_542) );
BUFx2_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
AND2x2_ASAP7_75t_L g533 ( .A(n_458), .B(n_487), .Y(n_533) );
INVx2_ASAP7_75t_L g549 ( .A(n_458), .Y(n_549) );
AND2x2_ASAP7_75t_L g558 ( .A(n_458), .B(n_486), .Y(n_558) );
AND2x2_ASAP7_75t_L g637 ( .A(n_458), .B(n_566), .Y(n_637) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_469), .Y(n_458) );
INVx2_ASAP7_75t_L g477 ( .A(n_463), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_499), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_471), .B(n_564), .Y(n_602) );
INVx1_ASAP7_75t_L g690 ( .A(n_471), .Y(n_690) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_486), .Y(n_471) );
AND2x2_ASAP7_75t_L g548 ( .A(n_472), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g562 ( .A(n_472), .B(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_472), .Y(n_591) );
OR2x2_ASAP7_75t_L g623 ( .A(n_472), .B(n_565), .Y(n_623) );
AND2x2_ASAP7_75t_L g631 ( .A(n_472), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g664 ( .A(n_472), .B(n_633), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_472), .B(n_533), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_472), .B(n_593), .Y(n_689) );
AND2x2_ASAP7_75t_L g695 ( .A(n_472), .B(n_582), .Y(n_695) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g555 ( .A(n_473), .Y(n_555) );
AND2x2_ASAP7_75t_L g585 ( .A(n_473), .B(n_565), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_473), .B(n_578), .Y(n_618) );
AND2x2_ASAP7_75t_L g638 ( .A(n_473), .B(n_487), .Y(n_638) );
AND2x2_ASAP7_75t_L g672 ( .A(n_473), .B(n_538), .Y(n_672) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_482), .C(n_483), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_480), .A2(n_483), .B(n_529), .C(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g578 ( .A(n_486), .B(n_549), .Y(n_578) );
AND2x2_ASAP7_75t_L g589 ( .A(n_486), .B(n_585), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_486), .B(n_565), .Y(n_628) );
INVx2_ASAP7_75t_L g643 ( .A(n_486), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_486), .B(n_577), .Y(n_666) );
AND2x2_ASAP7_75t_L g685 ( .A(n_486), .B(n_637), .Y(n_685) );
INVx5_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_487), .Y(n_584) );
AND2x2_ASAP7_75t_L g592 ( .A(n_487), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g633 ( .A(n_487), .B(n_549), .Y(n_633) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
AOI21xp5_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_491), .B(n_495), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
AND2x2_ASAP7_75t_L g556 ( .A(n_501), .B(n_539), .Y(n_556) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_502), .B(n_513), .Y(n_536) );
OR2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_539), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_502), .B(n_539), .Y(n_574) );
AND2x2_ASAP7_75t_L g601 ( .A(n_502), .B(n_538), .Y(n_601) );
AND2x2_ASAP7_75t_L g653 ( .A(n_502), .B(n_512), .Y(n_653) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_503), .B(n_523), .Y(n_561) );
AND2x2_ASAP7_75t_L g597 ( .A(n_503), .B(n_513), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_510), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g587 ( .A(n_511), .B(n_569), .Y(n_587) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
OAI322xp33_ASAP7_75t_L g552 ( .A1(n_512), .A2(n_553), .A3(n_557), .B1(n_559), .B2(n_562), .C1(n_567), .C2(n_575), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_512), .B(n_538), .Y(n_560) );
OR2x2_ASAP7_75t_L g570 ( .A(n_512), .B(n_524), .Y(n_570) );
AND2x2_ASAP7_75t_L g572 ( .A(n_512), .B(n_524), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_512), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_512), .B(n_539), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_512), .B(n_668), .Y(n_667) );
INVx5_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_513), .B(n_556), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_523), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g550 ( .A(n_523), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_523), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g612 ( .A(n_523), .B(n_539), .Y(n_612) );
AOI211xp5_ASAP7_75t_SL g640 ( .A1(n_523), .A2(n_641), .B(n_644), .C(n_656), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_523), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g678 ( .A(n_523), .B(n_653), .Y(n_678) );
INVx5_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g606 ( .A(n_524), .B(n_539), .Y(n_606) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_524), .Y(n_615) );
AND2x2_ASAP7_75t_L g655 ( .A(n_524), .B(n_653), .Y(n_655) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_524), .B(n_556), .Y(n_686) );
AND2x2_ASAP7_75t_L g693 ( .A(n_524), .B(n_652), .Y(n_693) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B1(n_548), .B2(n_550), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_533), .B(n_555), .Y(n_603) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g551 ( .A(n_536), .Y(n_551) );
OR2x2_ASAP7_75t_L g611 ( .A(n_536), .B(n_612), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_536), .A2(n_660), .B1(n_662), .B2(n_663), .C(n_665), .Y(n_659) );
INVx2_ASAP7_75t_L g598 ( .A(n_537), .Y(n_598) );
AND2x2_ASAP7_75t_L g571 ( .A(n_538), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g661 ( .A(n_538), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_538), .B(n_653), .Y(n_674) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_L g616 ( .A(n_539), .Y(n_616) );
AND2x2_ASAP7_75t_L g652 ( .A(n_539), .B(n_653), .Y(n_652) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_547), .Y(n_539) );
AND2x2_ASAP7_75t_L g654 ( .A(n_548), .B(n_593), .Y(n_654) );
AND2x2_ASAP7_75t_L g564 ( .A(n_549), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_549), .B(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g635 ( .A(n_551), .B(n_598), .Y(n_635) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g641 ( .A(n_554), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
OR2x2_ASAP7_75t_L g627 ( .A(n_555), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g692 ( .A(n_555), .B(n_637), .Y(n_692) );
INVx2_ASAP7_75t_L g625 ( .A(n_556), .Y(n_625) );
NAND4xp25_ASAP7_75t_SL g688 ( .A(n_557), .B(n_689), .C(n_690), .D(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_558), .B(n_622), .Y(n_657) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_SL g694 ( .A(n_561), .Y(n_694) );
O2A1O1Ixp33_ASAP7_75t_SL g656 ( .A1(n_562), .A2(n_625), .B(n_629), .C(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g651 ( .A(n_564), .B(n_643), .Y(n_651) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_565), .Y(n_577) );
INVx1_ASAP7_75t_L g632 ( .A(n_565), .Y(n_632) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_566), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_571), .C(n_573), .Y(n_567) );
AND2x2_ASAP7_75t_L g588 ( .A(n_568), .B(n_572), .Y(n_588) );
OAI322xp33_ASAP7_75t_SL g626 ( .A1(n_568), .A2(n_627), .A3(n_629), .B1(n_630), .B2(n_634), .C1(n_635), .C2(n_636), .Y(n_626) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g648 ( .A(n_570), .B(n_574), .Y(n_648) );
INVx1_ASAP7_75t_L g629 ( .A(n_572), .Y(n_629) );
INVx1_ASAP7_75t_SL g647 ( .A(n_574), .Y(n_647) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_586), .B1(n_588), .B2(n_589), .C1(n_590), .C2(n_730), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_581), .B(n_583), .Y(n_580) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_581), .A2(n_643), .A3(n_648), .B1(n_670), .B2(n_671), .C1(n_673), .C2(n_674), .Y(n_669) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_582), .A2(n_596), .B1(n_620), .B2(n_624), .C(n_626), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
OAI222xp33_ASAP7_75t_L g599 ( .A1(n_587), .A2(n_600), .B1(n_602), .B2(n_603), .C1(n_604), .C2(n_607), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_589), .A2(n_596), .B1(n_666), .B2(n_667), .Y(n_665) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AOI211xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_599), .C(n_610), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g675 ( .A1(n_596), .A2(n_633), .B(n_676), .C(n_679), .Y(n_675) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g605 ( .A(n_597), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g668 ( .A(n_601), .Y(n_668) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_608), .B(n_633), .Y(n_662) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B(n_617), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_611), .A2(n_680), .B1(n_681), .B2(n_682), .C(n_683), .Y(n_679) );
INVxp33_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_615), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_622), .B(n_633), .Y(n_673) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g684 ( .A(n_637), .B(n_643), .Y(n_684) );
AND4x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_658), .C(n_675), .D(n_687), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_646), .B1(n_648), .B2(n_649), .C(n_650), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_654), .B2(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g680 ( .A(n_651), .Y(n_680) );
INVx1_ASAP7_75t_SL g670 ( .A(n_655), .Y(n_670) );
NOR2xp33_ASAP7_75t_SL g658 ( .A(n_659), .B(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_671), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_678), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g706 ( .A(n_697), .Y(n_706) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx3_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g725 ( .A(n_713), .Y(n_725) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
XNOR2xp5_ASAP7_75t_SL g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
endmodule